magic
tech sky130A
magscale 1 2
timestamp 1698513452
<< nmos >>
rect -1132 -100 -932 100
rect -874 -100 -674 100
rect -616 -100 -416 100
rect -358 -100 -158 100
rect -100 -100 100 100
rect 158 -100 358 100
rect 416 -100 616 100
rect 674 -100 874 100
rect 932 -100 1132 100
<< ndiff >>
rect -1190 88 -1132 100
rect -1190 -88 -1178 88
rect -1144 -88 -1132 88
rect -1190 -100 -1132 -88
rect -932 88 -874 100
rect -932 -88 -920 88
rect -886 -88 -874 88
rect -932 -100 -874 -88
rect -674 88 -616 100
rect -674 -88 -662 88
rect -628 -88 -616 88
rect -674 -100 -616 -88
rect -416 88 -358 100
rect -416 -88 -404 88
rect -370 -88 -358 88
rect -416 -100 -358 -88
rect -158 88 -100 100
rect -158 -88 -146 88
rect -112 -88 -100 88
rect -158 -100 -100 -88
rect 100 88 158 100
rect 100 -88 112 88
rect 146 -88 158 88
rect 100 -100 158 -88
rect 358 88 416 100
rect 358 -88 370 88
rect 404 -88 416 88
rect 358 -100 416 -88
rect 616 88 674 100
rect 616 -88 628 88
rect 662 -88 674 88
rect 616 -100 674 -88
rect 874 88 932 100
rect 874 -88 886 88
rect 920 -88 932 88
rect 874 -100 932 -88
rect 1132 88 1190 100
rect 1132 -88 1144 88
rect 1178 -88 1190 88
rect 1132 -100 1190 -88
<< ndiffc >>
rect -1178 -88 -1144 88
rect -920 -88 -886 88
rect -662 -88 -628 88
rect -404 -88 -370 88
rect -146 -88 -112 88
rect 112 -88 146 88
rect 370 -88 404 88
rect 628 -88 662 88
rect 886 -88 920 88
rect 1144 -88 1178 88
<< poly >>
rect -1132 172 -932 188
rect -1132 138 -1116 172
rect -948 138 -932 172
rect -1132 100 -932 138
rect -874 172 -674 188
rect -874 138 -858 172
rect -690 138 -674 172
rect -874 100 -674 138
rect -616 172 -416 188
rect -616 138 -600 172
rect -432 138 -416 172
rect -616 100 -416 138
rect -358 172 -158 188
rect -358 138 -342 172
rect -174 138 -158 172
rect -358 100 -158 138
rect -100 172 100 188
rect -100 138 -84 172
rect 84 138 100 172
rect -100 100 100 138
rect 158 172 358 188
rect 158 138 174 172
rect 342 138 358 172
rect 158 100 358 138
rect 416 172 616 188
rect 416 138 432 172
rect 600 138 616 172
rect 416 100 616 138
rect 674 172 874 188
rect 674 138 690 172
rect 858 138 874 172
rect 674 100 874 138
rect 932 172 1132 188
rect 932 138 948 172
rect 1116 138 1132 172
rect 932 100 1132 138
rect -1132 -138 -932 -100
rect -1132 -172 -1116 -138
rect -948 -172 -932 -138
rect -1132 -188 -932 -172
rect -874 -138 -674 -100
rect -874 -172 -858 -138
rect -690 -172 -674 -138
rect -874 -188 -674 -172
rect -616 -138 -416 -100
rect -616 -172 -600 -138
rect -432 -172 -416 -138
rect -616 -188 -416 -172
rect -358 -138 -158 -100
rect -358 -172 -342 -138
rect -174 -172 -158 -138
rect -358 -188 -158 -172
rect -100 -138 100 -100
rect -100 -172 -84 -138
rect 84 -172 100 -138
rect -100 -188 100 -172
rect 158 -138 358 -100
rect 158 -172 174 -138
rect 342 -172 358 -138
rect 158 -188 358 -172
rect 416 -138 616 -100
rect 416 -172 432 -138
rect 600 -172 616 -138
rect 416 -188 616 -172
rect 674 -138 874 -100
rect 674 -172 690 -138
rect 858 -172 874 -138
rect 674 -188 874 -172
rect 932 -138 1132 -100
rect 932 -172 948 -138
rect 1116 -172 1132 -138
rect 932 -188 1132 -172
<< polycont >>
rect -1116 138 -948 172
rect -858 138 -690 172
rect -600 138 -432 172
rect -342 138 -174 172
rect -84 138 84 172
rect 174 138 342 172
rect 432 138 600 172
rect 690 138 858 172
rect 948 138 1116 172
rect -1116 -172 -948 -138
rect -858 -172 -690 -138
rect -600 -172 -432 -138
rect -342 -172 -174 -138
rect -84 -172 84 -138
rect 174 -172 342 -138
rect 432 -172 600 -138
rect 690 -172 858 -138
rect 948 -172 1116 -138
<< locali >>
rect -1132 138 -1116 172
rect -948 138 -932 172
rect -874 138 -858 172
rect -690 138 -674 172
rect -616 138 -600 172
rect -432 138 -416 172
rect -358 138 -342 172
rect -174 138 -158 172
rect -100 138 -84 172
rect 84 138 100 172
rect 158 138 174 172
rect 342 138 358 172
rect 416 138 432 172
rect 600 138 616 172
rect 674 138 690 172
rect 858 138 874 172
rect 932 138 948 172
rect 1116 138 1132 172
rect -1178 88 -1144 104
rect -1178 -104 -1144 -88
rect -920 88 -886 104
rect -920 -104 -886 -88
rect -662 88 -628 104
rect -662 -104 -628 -88
rect -404 88 -370 104
rect -404 -104 -370 -88
rect -146 88 -112 104
rect -146 -104 -112 -88
rect 112 88 146 104
rect 112 -104 146 -88
rect 370 88 404 104
rect 370 -104 404 -88
rect 628 88 662 104
rect 628 -104 662 -88
rect 886 88 920 104
rect 886 -104 920 -88
rect 1144 88 1178 104
rect 1144 -104 1178 -88
rect -1132 -172 -1116 -138
rect -948 -172 -932 -138
rect -874 -172 -858 -138
rect -690 -172 -674 -138
rect -616 -172 -600 -138
rect -432 -172 -416 -138
rect -358 -172 -342 -138
rect -174 -172 -158 -138
rect -100 -172 -84 -138
rect 84 -172 100 -138
rect 158 -172 174 -138
rect 342 -172 358 -138
rect 416 -172 432 -138
rect 600 -172 616 -138
rect 674 -172 690 -138
rect 858 -172 874 -138
rect 932 -172 948 -138
rect 1116 -172 1132 -138
<< viali >>
rect -1116 138 -948 172
rect -858 138 -690 172
rect -600 138 -432 172
rect -342 138 -174 172
rect -84 138 84 172
rect 174 138 342 172
rect 432 138 600 172
rect 690 138 858 172
rect 948 138 1116 172
rect -1178 -17 -1144 71
rect -920 -71 -886 17
rect -662 -17 -628 71
rect -404 -71 -370 17
rect -146 -17 -112 71
rect 112 -71 146 17
rect 370 -17 404 71
rect 628 -71 662 17
rect 886 -17 920 71
rect 1144 -71 1178 17
rect -1116 -172 -948 -138
rect -858 -172 -690 -138
rect -600 -172 -432 -138
rect -342 -172 -174 -138
rect -84 -172 84 -138
rect 174 -172 342 -138
rect 432 -172 600 -138
rect 690 -172 858 -138
rect 948 -172 1116 -138
<< metal1 >>
rect -1128 172 -936 178
rect -1128 138 -1116 172
rect -948 138 -936 172
rect -1128 132 -936 138
rect -870 172 -678 178
rect -870 138 -858 172
rect -690 138 -678 172
rect -870 132 -678 138
rect -612 172 -420 178
rect -612 138 -600 172
rect -432 138 -420 172
rect -612 132 -420 138
rect -354 172 -162 178
rect -354 138 -342 172
rect -174 138 -162 172
rect -354 132 -162 138
rect -96 172 96 178
rect -96 138 -84 172
rect 84 138 96 172
rect -96 132 96 138
rect 162 172 354 178
rect 162 138 174 172
rect 342 138 354 172
rect 162 132 354 138
rect 420 172 612 178
rect 420 138 432 172
rect 600 138 612 172
rect 420 132 612 138
rect 678 172 870 178
rect 678 138 690 172
rect 858 138 870 172
rect 678 132 870 138
rect 936 172 1128 178
rect 936 138 948 172
rect 1116 138 1128 172
rect 936 132 1128 138
rect -1184 71 -1138 83
rect -1184 -17 -1178 71
rect -1144 -17 -1138 71
rect -668 71 -622 83
rect -1184 -29 -1138 -17
rect -926 17 -880 29
rect -926 -71 -920 17
rect -886 -71 -880 17
rect -668 -17 -662 71
rect -628 -17 -622 71
rect -152 71 -106 83
rect -668 -29 -622 -17
rect -410 17 -364 29
rect -926 -83 -880 -71
rect -410 -71 -404 17
rect -370 -71 -364 17
rect -152 -17 -146 71
rect -112 -17 -106 71
rect 364 71 410 83
rect -152 -29 -106 -17
rect 106 17 152 29
rect -410 -83 -364 -71
rect 106 -71 112 17
rect 146 -71 152 17
rect 364 -17 370 71
rect 404 -17 410 71
rect 880 71 926 83
rect 364 -29 410 -17
rect 622 17 668 29
rect 106 -83 152 -71
rect 622 -71 628 17
rect 662 -71 668 17
rect 880 -17 886 71
rect 920 -17 926 71
rect 880 -29 926 -17
rect 1138 17 1184 29
rect 622 -83 668 -71
rect 1138 -71 1144 17
rect 1178 -71 1184 17
rect 1138 -83 1184 -71
rect -1128 -138 -936 -132
rect -1128 -172 -1116 -138
rect -948 -172 -936 -138
rect -1128 -178 -936 -172
rect -870 -138 -678 -132
rect -870 -172 -858 -138
rect -690 -172 -678 -138
rect -870 -178 -678 -172
rect -612 -138 -420 -132
rect -612 -172 -600 -138
rect -432 -172 -420 -138
rect -612 -178 -420 -172
rect -354 -138 -162 -132
rect -354 -172 -342 -138
rect -174 -172 -162 -138
rect -354 -178 -162 -172
rect -96 -138 96 -132
rect -96 -172 -84 -138
rect 84 -172 96 -138
rect -96 -178 96 -172
rect 162 -138 354 -132
rect 162 -172 174 -138
rect 342 -172 354 -138
rect 162 -178 354 -172
rect 420 -138 612 -132
rect 420 -172 432 -138
rect 600 -172 612 -138
rect 420 -178 612 -172
rect 678 -138 870 -132
rect 678 -172 690 -138
rect 858 -172 870 -138
rect 678 -178 870 -172
rect 936 -138 1128 -132
rect 936 -172 948 -138
rect 1116 -172 1128 -138
rect 936 -178 1128 -172
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 1.0 m 1 nf 9 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc +50 viadrn -50 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
