magic
tech sky130A
magscale 1 2
timestamp 1698511094
<< metal3 >>
rect -2550 1472 2549 1500
rect -2550 -1472 2465 1472
rect 2529 -1472 2549 1472
rect -2550 -1500 2549 -1472
<< via3 >>
rect 2465 -1472 2529 1472
<< mimcap >>
rect -2450 1360 2350 1400
rect -2450 -1360 -2410 1360
rect 2310 -1360 2350 1360
rect -2450 -1400 2350 -1360
<< mimcapcontact >>
rect -2410 -1360 2310 1360
<< metal4 >>
rect 2449 1472 2545 1488
rect -2411 1360 2311 1361
rect -2411 -1360 -2410 1360
rect 2310 -1360 2311 1360
rect -2411 -1361 2311 -1360
rect 2449 -1472 2465 1472
rect 2529 -1472 2545 1472
rect 2449 -1488 2545 -1472
<< properties >>
string FIXED_BBOX -2550 -1500 2450 1500
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 24 l 14 val 686.44 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
