magic
tech sky130A
magscale 1 2
timestamp 1698520721
<< pwell >>
rect -201 -650 201 650
<< psubdiff >>
rect -165 580 -69 614
rect 69 580 165 614
rect -165 518 -131 580
rect 131 518 165 580
rect -165 -580 -131 -518
rect 131 -580 165 -518
rect -165 -614 -69 -580
rect 69 -614 165 -580
<< psubdiffcont >>
rect -69 580 69 614
rect -165 -518 -131 518
rect 131 -518 165 518
rect -69 -614 69 -580
<< xpolycontact >>
rect -35 52 35 484
rect -35 -484 35 -52
<< xpolyres >>
rect -35 -52 35 52
<< locali >>
rect -165 580 -69 614
rect 69 580 165 614
rect -165 518 -131 580
rect 131 518 165 580
rect -165 -580 -131 -518
rect 131 -580 165 -518
rect -165 -614 -69 -580
rect 69 -614 165 -580
<< viali >>
rect -19 69 19 466
rect -19 -466 19 -69
<< metal1 >>
rect -25 466 25 478
rect -25 69 -19 466
rect 19 69 25 466
rect -25 57 25 69
rect -25 -69 25 -57
rect -25 -466 -19 -69
rect 19 -466 25 -69
rect -25 -478 25 -466
<< res0p35 >>
rect -37 -54 37 54
<< properties >>
string FIXED_BBOX -148 -597 148 597
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 0.52 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 4.046k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
