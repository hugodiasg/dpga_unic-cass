magic
tech sky130A
magscale 1 2
timestamp 1698520721
<< error_p >>
rect -461 581 -403 587
rect -269 581 -211 587
rect -77 581 -19 587
rect 115 581 173 587
rect 307 581 365 587
rect 499 581 557 587
rect -461 547 -449 581
rect -269 547 -257 581
rect -77 547 -65 581
rect 115 547 127 581
rect 307 547 319 581
rect 499 547 511 581
rect -461 541 -403 547
rect -269 541 -211 547
rect -77 541 -19 547
rect 115 541 173 547
rect 307 541 365 547
rect 499 541 557 547
rect -557 -547 -499 -541
rect -365 -547 -307 -541
rect -173 -547 -115 -541
rect 19 -547 77 -541
rect 211 -547 269 -541
rect 403 -547 461 -541
rect -557 -581 -545 -547
rect -365 -581 -353 -547
rect -173 -581 -161 -547
rect 19 -581 31 -547
rect 211 -581 223 -547
rect 403 -581 415 -547
rect -557 -587 -499 -581
rect -365 -587 -307 -581
rect -173 -587 -115 -581
rect 19 -587 77 -581
rect 211 -587 269 -581
rect 403 -587 461 -581
<< nwell >>
rect -743 -719 743 719
<< pmos >>
rect -543 -500 -513 500
rect -447 -500 -417 500
rect -351 -500 -321 500
rect -255 -500 -225 500
rect -159 -500 -129 500
rect -63 -500 -33 500
rect 33 -500 63 500
rect 129 -500 159 500
rect 225 -500 255 500
rect 321 -500 351 500
rect 417 -500 447 500
rect 513 -500 543 500
<< pdiff >>
rect -605 488 -543 500
rect -605 -488 -593 488
rect -559 -488 -543 488
rect -605 -500 -543 -488
rect -513 488 -447 500
rect -513 -488 -497 488
rect -463 -488 -447 488
rect -513 -500 -447 -488
rect -417 488 -351 500
rect -417 -488 -401 488
rect -367 -488 -351 488
rect -417 -500 -351 -488
rect -321 488 -255 500
rect -321 -488 -305 488
rect -271 -488 -255 488
rect -321 -500 -255 -488
rect -225 488 -159 500
rect -225 -488 -209 488
rect -175 -488 -159 488
rect -225 -500 -159 -488
rect -129 488 -63 500
rect -129 -488 -113 488
rect -79 -488 -63 488
rect -129 -500 -63 -488
rect -33 488 33 500
rect -33 -488 -17 488
rect 17 -488 33 488
rect -33 -500 33 -488
rect 63 488 129 500
rect 63 -488 79 488
rect 113 -488 129 488
rect 63 -500 129 -488
rect 159 488 225 500
rect 159 -488 175 488
rect 209 -488 225 488
rect 159 -500 225 -488
rect 255 488 321 500
rect 255 -488 271 488
rect 305 -488 321 488
rect 255 -500 321 -488
rect 351 488 417 500
rect 351 -488 367 488
rect 401 -488 417 488
rect 351 -500 417 -488
rect 447 488 513 500
rect 447 -488 463 488
rect 497 -488 513 488
rect 447 -500 513 -488
rect 543 488 605 500
rect 543 -488 559 488
rect 593 -488 605 488
rect 543 -500 605 -488
<< pdiffc >>
rect -593 -488 -559 488
rect -497 -488 -463 488
rect -401 -488 -367 488
rect -305 -488 -271 488
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
rect 271 -488 305 488
rect 367 -488 401 488
rect 463 -488 497 488
rect 559 -488 593 488
<< nsubdiff >>
rect -707 649 -611 683
rect 611 649 707 683
rect -707 587 -673 649
rect 673 587 707 649
rect -707 -649 -673 -587
rect 673 -649 707 -587
rect -707 -683 -611 -649
rect 611 -683 707 -649
<< nsubdiffcont >>
rect -611 649 611 683
rect -707 -587 -673 587
rect 673 -587 707 587
rect -611 -683 611 -649
<< poly >>
rect -465 581 -399 597
rect -465 547 -449 581
rect -415 547 -399 581
rect -465 531 -399 547
rect -273 581 -207 597
rect -273 547 -257 581
rect -223 547 -207 581
rect -273 531 -207 547
rect -81 581 -15 597
rect -81 547 -65 581
rect -31 547 -15 581
rect -81 531 -15 547
rect 111 581 177 597
rect 111 547 127 581
rect 161 547 177 581
rect 111 531 177 547
rect 303 581 369 597
rect 303 547 319 581
rect 353 547 369 581
rect 303 531 369 547
rect 495 581 561 597
rect 495 547 511 581
rect 545 547 561 581
rect 495 531 561 547
rect -543 500 -513 526
rect -447 500 -417 531
rect -351 500 -321 526
rect -255 500 -225 531
rect -159 500 -129 526
rect -63 500 -33 531
rect 33 500 63 526
rect 129 500 159 531
rect 225 500 255 526
rect 321 500 351 531
rect 417 500 447 526
rect 513 500 543 531
rect -543 -531 -513 -500
rect -447 -526 -417 -500
rect -351 -531 -321 -500
rect -255 -526 -225 -500
rect -159 -531 -129 -500
rect -63 -526 -33 -500
rect 33 -531 63 -500
rect 129 -526 159 -500
rect 225 -531 255 -500
rect 321 -526 351 -500
rect 417 -531 447 -500
rect 513 -526 543 -500
rect -561 -547 -495 -531
rect -561 -581 -545 -547
rect -511 -581 -495 -547
rect -561 -597 -495 -581
rect -369 -547 -303 -531
rect -369 -581 -353 -547
rect -319 -581 -303 -547
rect -369 -597 -303 -581
rect -177 -547 -111 -531
rect -177 -581 -161 -547
rect -127 -581 -111 -547
rect -177 -597 -111 -581
rect 15 -547 81 -531
rect 15 -581 31 -547
rect 65 -581 81 -547
rect 15 -597 81 -581
rect 207 -547 273 -531
rect 207 -581 223 -547
rect 257 -581 273 -547
rect 207 -597 273 -581
rect 399 -547 465 -531
rect 399 -581 415 -547
rect 449 -581 465 -547
rect 399 -597 465 -581
<< polycont >>
rect -449 547 -415 581
rect -257 547 -223 581
rect -65 547 -31 581
rect 127 547 161 581
rect 319 547 353 581
rect 511 547 545 581
rect -545 -581 -511 -547
rect -353 -581 -319 -547
rect -161 -581 -127 -547
rect 31 -581 65 -547
rect 223 -581 257 -547
rect 415 -581 449 -547
<< locali >>
rect -707 649 -611 683
rect 611 649 707 683
rect -707 587 -673 649
rect 673 587 707 649
rect -465 547 -449 581
rect -415 547 -399 581
rect -273 547 -257 581
rect -223 547 -207 581
rect -81 547 -65 581
rect -31 547 -15 581
rect 111 547 127 581
rect 161 547 177 581
rect 303 547 319 581
rect 353 547 369 581
rect 495 547 511 581
rect 545 547 561 581
rect -593 488 -559 504
rect -593 -504 -559 -488
rect -497 488 -463 504
rect -497 -504 -463 -488
rect -401 488 -367 504
rect -401 -504 -367 -488
rect -305 488 -271 504
rect -305 -504 -271 -488
rect -209 488 -175 504
rect -209 -504 -175 -488
rect -113 488 -79 504
rect -113 -504 -79 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 79 488 113 504
rect 79 -504 113 -488
rect 175 488 209 504
rect 175 -504 209 -488
rect 271 488 305 504
rect 271 -504 305 -488
rect 367 488 401 504
rect 367 -504 401 -488
rect 463 488 497 504
rect 463 -504 497 -488
rect 559 488 593 504
rect 559 -504 593 -488
rect -561 -581 -545 -547
rect -511 -581 -495 -547
rect -369 -581 -353 -547
rect -319 -581 -303 -547
rect -177 -581 -161 -547
rect -127 -581 -111 -547
rect 15 -581 31 -547
rect 65 -581 81 -547
rect 207 -581 223 -547
rect 257 -581 273 -547
rect 399 -581 415 -547
rect 449 -581 465 -547
rect -707 -649 -673 -587
rect 673 -649 707 -587
rect -707 -683 -611 -649
rect 611 -683 707 -649
<< viali >>
rect -449 547 -415 581
rect -257 547 -223 581
rect -65 547 -31 581
rect 127 547 161 581
rect 319 547 353 581
rect 511 547 545 581
rect -593 -488 -559 488
rect -497 -488 -463 488
rect -401 -488 -367 488
rect -305 -488 -271 488
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
rect 271 -488 305 488
rect 367 -488 401 488
rect 463 -488 497 488
rect 559 -488 593 488
rect -545 -581 -511 -547
rect -353 -581 -319 -547
rect -161 -581 -127 -547
rect 31 -581 65 -547
rect 223 -581 257 -547
rect 415 -581 449 -547
<< metal1 >>
rect -461 581 -403 587
rect -461 547 -449 581
rect -415 547 -403 581
rect -461 541 -403 547
rect -269 581 -211 587
rect -269 547 -257 581
rect -223 547 -211 581
rect -269 541 -211 547
rect -77 581 -19 587
rect -77 547 -65 581
rect -31 547 -19 581
rect -77 541 -19 547
rect 115 581 173 587
rect 115 547 127 581
rect 161 547 173 581
rect 115 541 173 547
rect 307 581 365 587
rect 307 547 319 581
rect 353 547 365 581
rect 307 541 365 547
rect 499 581 557 587
rect 499 547 511 581
rect 545 547 557 581
rect 499 541 557 547
rect -599 488 -553 500
rect -599 -488 -593 488
rect -559 -488 -553 488
rect -599 -500 -553 -488
rect -503 488 -457 500
rect -503 -488 -497 488
rect -463 -488 -457 488
rect -503 -500 -457 -488
rect -407 488 -361 500
rect -407 -488 -401 488
rect -367 -488 -361 488
rect -407 -500 -361 -488
rect -311 488 -265 500
rect -311 -488 -305 488
rect -271 -488 -265 488
rect -311 -500 -265 -488
rect -215 488 -169 500
rect -215 -488 -209 488
rect -175 -488 -169 488
rect -215 -500 -169 -488
rect -119 488 -73 500
rect -119 -488 -113 488
rect -79 -488 -73 488
rect -119 -500 -73 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 73 488 119 500
rect 73 -488 79 488
rect 113 -488 119 488
rect 73 -500 119 -488
rect 169 488 215 500
rect 169 -488 175 488
rect 209 -488 215 488
rect 169 -500 215 -488
rect 265 488 311 500
rect 265 -488 271 488
rect 305 -488 311 488
rect 265 -500 311 -488
rect 361 488 407 500
rect 361 -488 367 488
rect 401 -488 407 488
rect 361 -500 407 -488
rect 457 488 503 500
rect 457 -488 463 488
rect 497 -488 503 488
rect 457 -500 503 -488
rect 553 488 599 500
rect 553 -488 559 488
rect 593 -488 599 488
rect 553 -500 599 -488
rect -557 -547 -499 -541
rect -557 -581 -545 -547
rect -511 -581 -499 -547
rect -557 -587 -499 -581
rect -365 -547 -307 -541
rect -365 -581 -353 -547
rect -319 -581 -307 -547
rect -365 -587 -307 -581
rect -173 -547 -115 -541
rect -173 -581 -161 -547
rect -127 -581 -115 -547
rect -173 -587 -115 -581
rect 19 -547 77 -541
rect 19 -581 31 -547
rect 65 -581 77 -547
rect 19 -587 77 -581
rect 211 -547 269 -541
rect 211 -581 223 -547
rect 257 -581 269 -547
rect 211 -587 269 -581
rect 403 -547 461 -541
rect 403 -581 415 -547
rect 449 -581 461 -547
rect 403 -587 461 -581
<< properties >>
string FIXED_BBOX -690 -666 690 666
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.0 l 0.15 m 1 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
