magic
tech sky130A
magscale 1 2
timestamp 1698430755
<< viali >>
rect 2421 17221 2455 17255
rect 15393 17221 15427 17255
rect 11161 17153 11195 17187
rect 2513 16949 2547 16983
rect 10977 16949 11011 16983
rect 15485 16949 15519 16983
rect 5917 5117 5951 5151
rect 8401 5117 8435 5151
rect 5273 4981 5307 5015
rect 7849 4981 7883 5015
rect 6837 4709 6871 4743
rect 8401 4641 8435 4675
rect 10425 4641 10459 4675
rect 4997 4573 5031 4607
rect 7021 4573 7055 4607
rect 8217 4573 8251 4607
rect 10241 4573 10275 4607
rect 5273 4505 5307 4539
rect 6745 4437 6779 4471
rect 7849 4437 7883 4471
rect 8309 4437 8343 4471
rect 9873 4437 9907 4471
rect 10333 4437 10367 4471
rect 5273 4233 5307 4267
rect 5641 4233 5675 4267
rect 6101 4233 6135 4267
rect 7297 4165 7331 4199
rect 4813 4097 4847 4131
rect 5089 4097 5123 4131
rect 5733 4097 5767 4131
rect 6377 4097 6411 4131
rect 9137 4097 9171 4131
rect 5457 4029 5491 4063
rect 7021 4029 7055 4063
rect 9413 4029 9447 4063
rect 9689 4029 9723 4063
rect 9321 3961 9355 3995
rect 4997 3893 5031 3927
rect 8585 3893 8619 3927
rect 11161 3893 11195 3927
rect 4721 3689 4755 3723
rect 5089 3689 5123 3723
rect 8401 3689 8435 3723
rect 10885 3689 10919 3723
rect 4169 3553 4203 3587
rect 6653 3553 6687 3587
rect 4353 3485 4387 3519
rect 6561 3485 6595 3519
rect 8585 3485 8619 3519
rect 9597 3485 9631 3519
rect 11621 3485 11655 3519
rect 6929 3417 6963 3451
rect 4261 3349 4295 3383
rect 8769 3349 8803 3383
rect 11437 3349 11471 3383
rect 4353 3145 4387 3179
rect 6745 3077 6779 3111
rect 4445 3009 4479 3043
rect 6837 3009 6871 3043
rect 9045 3009 9079 3043
rect 9137 3009 9171 3043
rect 3709 2941 3743 2975
rect 4721 2941 4755 2975
rect 6561 2941 6595 2975
rect 8769 2941 8803 2975
rect 9413 2941 9447 2975
rect 10885 2941 10919 2975
rect 12081 2941 12115 2975
rect 7205 2873 7239 2907
rect 6193 2805 6227 2839
rect 7297 2805 7331 2839
rect 11529 2805 11563 2839
rect 6561 2601 6595 2635
rect 7297 2601 7331 2635
rect 9137 2601 9171 2635
rect 11069 2601 11103 2635
rect 10793 2533 10827 2567
rect 4445 2465 4479 2499
rect 5917 2465 5951 2499
rect 6193 2465 6227 2499
rect 7113 2465 7147 2499
rect 9689 2465 9723 2499
rect 10149 2465 10183 2499
rect 10333 2465 10367 2499
rect 1777 2397 1811 2431
rect 4169 2397 4203 2431
rect 7481 2397 7515 2431
rect 7941 2397 7975 2431
rect 8217 2397 8251 2431
rect 9505 2397 9539 2431
rect 10425 2397 10459 2431
rect 12081 2397 12115 2431
rect 16037 2397 16071 2431
rect 1409 2329 1443 2363
rect 3801 2329 3835 2363
rect 10977 2329 11011 2363
rect 14197 2329 14231 2363
rect 7665 2261 7699 2295
rect 8309 2261 8343 2295
rect 9597 2261 9631 2295
rect 12173 2261 12207 2295
rect 14289 2261 14323 2295
<< metal1 >>
rect 1104 17434 16376 17456
rect 1104 17382 3519 17434
rect 3571 17382 3583 17434
rect 3635 17382 3647 17434
rect 3699 17382 3711 17434
rect 3763 17382 3775 17434
rect 3827 17382 7337 17434
rect 7389 17382 7401 17434
rect 7453 17382 7465 17434
rect 7517 17382 7529 17434
rect 7581 17382 7593 17434
rect 7645 17382 11155 17434
rect 11207 17382 11219 17434
rect 11271 17382 11283 17434
rect 11335 17382 11347 17434
rect 11399 17382 11411 17434
rect 11463 17382 14973 17434
rect 15025 17382 15037 17434
rect 15089 17382 15101 17434
rect 15153 17382 15165 17434
rect 15217 17382 15229 17434
rect 15281 17382 16376 17434
rect 1104 17360 16376 17382
rect 11054 17280 11060 17332
rect 11112 17280 11118 17332
rect 2222 17212 2228 17264
rect 2280 17252 2286 17264
rect 2409 17255 2467 17261
rect 2409 17252 2421 17255
rect 2280 17224 2421 17252
rect 2280 17212 2286 17224
rect 2409 17221 2421 17224
rect 2455 17221 2467 17255
rect 2409 17215 2467 17221
rect 11072 17184 11100 17280
rect 15378 17212 15384 17264
rect 15436 17212 15442 17264
rect 11149 17187 11207 17193
rect 11149 17184 11161 17187
rect 11072 17156 11161 17184
rect 11149 17153 11161 17156
rect 11195 17153 11207 17187
rect 11149 17147 11207 17153
rect 2498 16940 2504 16992
rect 2556 16940 2562 16992
rect 10226 16940 10232 16992
rect 10284 16980 10290 16992
rect 10965 16983 11023 16989
rect 10965 16980 10977 16983
rect 10284 16952 10977 16980
rect 10284 16940 10290 16952
rect 10965 16949 10977 16952
rect 11011 16949 11023 16983
rect 10965 16943 11023 16949
rect 15470 16940 15476 16992
rect 15528 16940 15534 16992
rect 1104 16890 16376 16912
rect 1104 16838 2859 16890
rect 2911 16838 2923 16890
rect 2975 16838 2987 16890
rect 3039 16838 3051 16890
rect 3103 16838 3115 16890
rect 3167 16838 6677 16890
rect 6729 16838 6741 16890
rect 6793 16838 6805 16890
rect 6857 16838 6869 16890
rect 6921 16838 6933 16890
rect 6985 16838 10495 16890
rect 10547 16838 10559 16890
rect 10611 16838 10623 16890
rect 10675 16838 10687 16890
rect 10739 16838 10751 16890
rect 10803 16838 14313 16890
rect 14365 16838 14377 16890
rect 14429 16838 14441 16890
rect 14493 16838 14505 16890
rect 14557 16838 14569 16890
rect 14621 16838 16376 16890
rect 1104 16816 16376 16838
rect 1104 16346 16376 16368
rect 1104 16294 3519 16346
rect 3571 16294 3583 16346
rect 3635 16294 3647 16346
rect 3699 16294 3711 16346
rect 3763 16294 3775 16346
rect 3827 16294 7337 16346
rect 7389 16294 7401 16346
rect 7453 16294 7465 16346
rect 7517 16294 7529 16346
rect 7581 16294 7593 16346
rect 7645 16294 11155 16346
rect 11207 16294 11219 16346
rect 11271 16294 11283 16346
rect 11335 16294 11347 16346
rect 11399 16294 11411 16346
rect 11463 16294 14973 16346
rect 15025 16294 15037 16346
rect 15089 16294 15101 16346
rect 15153 16294 15165 16346
rect 15217 16294 15229 16346
rect 15281 16294 16376 16346
rect 1104 16272 16376 16294
rect 1104 15802 16376 15824
rect 1104 15750 2859 15802
rect 2911 15750 2923 15802
rect 2975 15750 2987 15802
rect 3039 15750 3051 15802
rect 3103 15750 3115 15802
rect 3167 15750 6677 15802
rect 6729 15750 6741 15802
rect 6793 15750 6805 15802
rect 6857 15750 6869 15802
rect 6921 15750 6933 15802
rect 6985 15750 10495 15802
rect 10547 15750 10559 15802
rect 10611 15750 10623 15802
rect 10675 15750 10687 15802
rect 10739 15750 10751 15802
rect 10803 15750 14313 15802
rect 14365 15750 14377 15802
rect 14429 15750 14441 15802
rect 14493 15750 14505 15802
rect 14557 15750 14569 15802
rect 14621 15750 16376 15802
rect 1104 15728 16376 15750
rect 6546 15308 6552 15360
rect 6604 15348 6610 15360
rect 7190 15348 7196 15360
rect 6604 15320 7196 15348
rect 6604 15308 6610 15320
rect 7190 15308 7196 15320
rect 7248 15308 7254 15360
rect 1104 15258 16376 15280
rect 1104 15206 3519 15258
rect 3571 15206 3583 15258
rect 3635 15206 3647 15258
rect 3699 15206 3711 15258
rect 3763 15206 3775 15258
rect 3827 15206 7337 15258
rect 7389 15206 7401 15258
rect 7453 15206 7465 15258
rect 7517 15206 7529 15258
rect 7581 15206 7593 15258
rect 7645 15206 11155 15258
rect 11207 15206 11219 15258
rect 11271 15206 11283 15258
rect 11335 15206 11347 15258
rect 11399 15206 11411 15258
rect 11463 15206 14973 15258
rect 15025 15206 15037 15258
rect 15089 15206 15101 15258
rect 15153 15206 15165 15258
rect 15217 15206 15229 15258
rect 15281 15206 16376 15258
rect 1104 15184 16376 15206
rect 1104 14714 16376 14736
rect 1104 14662 2859 14714
rect 2911 14662 2923 14714
rect 2975 14662 2987 14714
rect 3039 14662 3051 14714
rect 3103 14662 3115 14714
rect 3167 14662 6677 14714
rect 6729 14662 6741 14714
rect 6793 14662 6805 14714
rect 6857 14662 6869 14714
rect 6921 14662 6933 14714
rect 6985 14662 10495 14714
rect 10547 14662 10559 14714
rect 10611 14662 10623 14714
rect 10675 14662 10687 14714
rect 10739 14662 10751 14714
rect 10803 14662 14313 14714
rect 14365 14662 14377 14714
rect 14429 14662 14441 14714
rect 14493 14662 14505 14714
rect 14557 14662 14569 14714
rect 14621 14662 16376 14714
rect 1104 14640 16376 14662
rect 1104 14170 16376 14192
rect 1104 14118 3519 14170
rect 3571 14118 3583 14170
rect 3635 14118 3647 14170
rect 3699 14118 3711 14170
rect 3763 14118 3775 14170
rect 3827 14118 7337 14170
rect 7389 14118 7401 14170
rect 7453 14118 7465 14170
rect 7517 14118 7529 14170
rect 7581 14118 7593 14170
rect 7645 14118 11155 14170
rect 11207 14118 11219 14170
rect 11271 14118 11283 14170
rect 11335 14118 11347 14170
rect 11399 14118 11411 14170
rect 11463 14118 14973 14170
rect 15025 14118 15037 14170
rect 15089 14118 15101 14170
rect 15153 14118 15165 14170
rect 15217 14118 15229 14170
rect 15281 14118 16376 14170
rect 1104 14096 16376 14118
rect 1104 13626 16376 13648
rect 1104 13574 2859 13626
rect 2911 13574 2923 13626
rect 2975 13574 2987 13626
rect 3039 13574 3051 13626
rect 3103 13574 3115 13626
rect 3167 13574 6677 13626
rect 6729 13574 6741 13626
rect 6793 13574 6805 13626
rect 6857 13574 6869 13626
rect 6921 13574 6933 13626
rect 6985 13574 10495 13626
rect 10547 13574 10559 13626
rect 10611 13574 10623 13626
rect 10675 13574 10687 13626
rect 10739 13574 10751 13626
rect 10803 13574 14313 13626
rect 14365 13574 14377 13626
rect 14429 13574 14441 13626
rect 14493 13574 14505 13626
rect 14557 13574 14569 13626
rect 14621 13574 16376 13626
rect 1104 13552 16376 13574
rect 1104 13082 16376 13104
rect 1104 13030 3519 13082
rect 3571 13030 3583 13082
rect 3635 13030 3647 13082
rect 3699 13030 3711 13082
rect 3763 13030 3775 13082
rect 3827 13030 7337 13082
rect 7389 13030 7401 13082
rect 7453 13030 7465 13082
rect 7517 13030 7529 13082
rect 7581 13030 7593 13082
rect 7645 13030 11155 13082
rect 11207 13030 11219 13082
rect 11271 13030 11283 13082
rect 11335 13030 11347 13082
rect 11399 13030 11411 13082
rect 11463 13030 14973 13082
rect 15025 13030 15037 13082
rect 15089 13030 15101 13082
rect 15153 13030 15165 13082
rect 15217 13030 15229 13082
rect 15281 13030 16376 13082
rect 1104 13008 16376 13030
rect 1104 12538 16376 12560
rect 1104 12486 2859 12538
rect 2911 12486 2923 12538
rect 2975 12486 2987 12538
rect 3039 12486 3051 12538
rect 3103 12486 3115 12538
rect 3167 12486 6677 12538
rect 6729 12486 6741 12538
rect 6793 12486 6805 12538
rect 6857 12486 6869 12538
rect 6921 12486 6933 12538
rect 6985 12486 10495 12538
rect 10547 12486 10559 12538
rect 10611 12486 10623 12538
rect 10675 12486 10687 12538
rect 10739 12486 10751 12538
rect 10803 12486 14313 12538
rect 14365 12486 14377 12538
rect 14429 12486 14441 12538
rect 14493 12486 14505 12538
rect 14557 12486 14569 12538
rect 14621 12486 16376 12538
rect 1104 12464 16376 12486
rect 1104 11994 16376 12016
rect 1104 11942 3519 11994
rect 3571 11942 3583 11994
rect 3635 11942 3647 11994
rect 3699 11942 3711 11994
rect 3763 11942 3775 11994
rect 3827 11942 7337 11994
rect 7389 11942 7401 11994
rect 7453 11942 7465 11994
rect 7517 11942 7529 11994
rect 7581 11942 7593 11994
rect 7645 11942 11155 11994
rect 11207 11942 11219 11994
rect 11271 11942 11283 11994
rect 11335 11942 11347 11994
rect 11399 11942 11411 11994
rect 11463 11942 14973 11994
rect 15025 11942 15037 11994
rect 15089 11942 15101 11994
rect 15153 11942 15165 11994
rect 15217 11942 15229 11994
rect 15281 11942 16376 11994
rect 1104 11920 16376 11942
rect 1104 11450 16376 11472
rect 1104 11398 2859 11450
rect 2911 11398 2923 11450
rect 2975 11398 2987 11450
rect 3039 11398 3051 11450
rect 3103 11398 3115 11450
rect 3167 11398 6677 11450
rect 6729 11398 6741 11450
rect 6793 11398 6805 11450
rect 6857 11398 6869 11450
rect 6921 11398 6933 11450
rect 6985 11398 10495 11450
rect 10547 11398 10559 11450
rect 10611 11398 10623 11450
rect 10675 11398 10687 11450
rect 10739 11398 10751 11450
rect 10803 11398 14313 11450
rect 14365 11398 14377 11450
rect 14429 11398 14441 11450
rect 14493 11398 14505 11450
rect 14557 11398 14569 11450
rect 14621 11398 16376 11450
rect 1104 11376 16376 11398
rect 1104 10906 16376 10928
rect 1104 10854 3519 10906
rect 3571 10854 3583 10906
rect 3635 10854 3647 10906
rect 3699 10854 3711 10906
rect 3763 10854 3775 10906
rect 3827 10854 7337 10906
rect 7389 10854 7401 10906
rect 7453 10854 7465 10906
rect 7517 10854 7529 10906
rect 7581 10854 7593 10906
rect 7645 10854 11155 10906
rect 11207 10854 11219 10906
rect 11271 10854 11283 10906
rect 11335 10854 11347 10906
rect 11399 10854 11411 10906
rect 11463 10854 14973 10906
rect 15025 10854 15037 10906
rect 15089 10854 15101 10906
rect 15153 10854 15165 10906
rect 15217 10854 15229 10906
rect 15281 10854 16376 10906
rect 1104 10832 16376 10854
rect 1104 10362 16376 10384
rect 1104 10310 2859 10362
rect 2911 10310 2923 10362
rect 2975 10310 2987 10362
rect 3039 10310 3051 10362
rect 3103 10310 3115 10362
rect 3167 10310 6677 10362
rect 6729 10310 6741 10362
rect 6793 10310 6805 10362
rect 6857 10310 6869 10362
rect 6921 10310 6933 10362
rect 6985 10310 10495 10362
rect 10547 10310 10559 10362
rect 10611 10310 10623 10362
rect 10675 10310 10687 10362
rect 10739 10310 10751 10362
rect 10803 10310 14313 10362
rect 14365 10310 14377 10362
rect 14429 10310 14441 10362
rect 14493 10310 14505 10362
rect 14557 10310 14569 10362
rect 14621 10310 16376 10362
rect 1104 10288 16376 10310
rect 1104 9818 16376 9840
rect 1104 9766 3519 9818
rect 3571 9766 3583 9818
rect 3635 9766 3647 9818
rect 3699 9766 3711 9818
rect 3763 9766 3775 9818
rect 3827 9766 7337 9818
rect 7389 9766 7401 9818
rect 7453 9766 7465 9818
rect 7517 9766 7529 9818
rect 7581 9766 7593 9818
rect 7645 9766 11155 9818
rect 11207 9766 11219 9818
rect 11271 9766 11283 9818
rect 11335 9766 11347 9818
rect 11399 9766 11411 9818
rect 11463 9766 14973 9818
rect 15025 9766 15037 9818
rect 15089 9766 15101 9818
rect 15153 9766 15165 9818
rect 15217 9766 15229 9818
rect 15281 9766 16376 9818
rect 1104 9744 16376 9766
rect 1104 9274 16376 9296
rect 1104 9222 2859 9274
rect 2911 9222 2923 9274
rect 2975 9222 2987 9274
rect 3039 9222 3051 9274
rect 3103 9222 3115 9274
rect 3167 9222 6677 9274
rect 6729 9222 6741 9274
rect 6793 9222 6805 9274
rect 6857 9222 6869 9274
rect 6921 9222 6933 9274
rect 6985 9222 10495 9274
rect 10547 9222 10559 9274
rect 10611 9222 10623 9274
rect 10675 9222 10687 9274
rect 10739 9222 10751 9274
rect 10803 9222 14313 9274
rect 14365 9222 14377 9274
rect 14429 9222 14441 9274
rect 14493 9222 14505 9274
rect 14557 9222 14569 9274
rect 14621 9222 16376 9274
rect 1104 9200 16376 9222
rect 1104 8730 16376 8752
rect 1104 8678 3519 8730
rect 3571 8678 3583 8730
rect 3635 8678 3647 8730
rect 3699 8678 3711 8730
rect 3763 8678 3775 8730
rect 3827 8678 7337 8730
rect 7389 8678 7401 8730
rect 7453 8678 7465 8730
rect 7517 8678 7529 8730
rect 7581 8678 7593 8730
rect 7645 8678 11155 8730
rect 11207 8678 11219 8730
rect 11271 8678 11283 8730
rect 11335 8678 11347 8730
rect 11399 8678 11411 8730
rect 11463 8678 14973 8730
rect 15025 8678 15037 8730
rect 15089 8678 15101 8730
rect 15153 8678 15165 8730
rect 15217 8678 15229 8730
rect 15281 8678 16376 8730
rect 1104 8656 16376 8678
rect 1104 8186 16376 8208
rect 1104 8134 2859 8186
rect 2911 8134 2923 8186
rect 2975 8134 2987 8186
rect 3039 8134 3051 8186
rect 3103 8134 3115 8186
rect 3167 8134 6677 8186
rect 6729 8134 6741 8186
rect 6793 8134 6805 8186
rect 6857 8134 6869 8186
rect 6921 8134 6933 8186
rect 6985 8134 10495 8186
rect 10547 8134 10559 8186
rect 10611 8134 10623 8186
rect 10675 8134 10687 8186
rect 10739 8134 10751 8186
rect 10803 8134 14313 8186
rect 14365 8134 14377 8186
rect 14429 8134 14441 8186
rect 14493 8134 14505 8186
rect 14557 8134 14569 8186
rect 14621 8134 16376 8186
rect 1104 8112 16376 8134
rect 1104 7642 16376 7664
rect 1104 7590 3519 7642
rect 3571 7590 3583 7642
rect 3635 7590 3647 7642
rect 3699 7590 3711 7642
rect 3763 7590 3775 7642
rect 3827 7590 7337 7642
rect 7389 7590 7401 7642
rect 7453 7590 7465 7642
rect 7517 7590 7529 7642
rect 7581 7590 7593 7642
rect 7645 7590 11155 7642
rect 11207 7590 11219 7642
rect 11271 7590 11283 7642
rect 11335 7590 11347 7642
rect 11399 7590 11411 7642
rect 11463 7590 14973 7642
rect 15025 7590 15037 7642
rect 15089 7590 15101 7642
rect 15153 7590 15165 7642
rect 15217 7590 15229 7642
rect 15281 7590 16376 7642
rect 1104 7568 16376 7590
rect 1104 7098 16376 7120
rect 1104 7046 2859 7098
rect 2911 7046 2923 7098
rect 2975 7046 2987 7098
rect 3039 7046 3051 7098
rect 3103 7046 3115 7098
rect 3167 7046 6677 7098
rect 6729 7046 6741 7098
rect 6793 7046 6805 7098
rect 6857 7046 6869 7098
rect 6921 7046 6933 7098
rect 6985 7046 10495 7098
rect 10547 7046 10559 7098
rect 10611 7046 10623 7098
rect 10675 7046 10687 7098
rect 10739 7046 10751 7098
rect 10803 7046 14313 7098
rect 14365 7046 14377 7098
rect 14429 7046 14441 7098
rect 14493 7046 14505 7098
rect 14557 7046 14569 7098
rect 14621 7046 16376 7098
rect 1104 7024 16376 7046
rect 1104 6554 16376 6576
rect 1104 6502 3519 6554
rect 3571 6502 3583 6554
rect 3635 6502 3647 6554
rect 3699 6502 3711 6554
rect 3763 6502 3775 6554
rect 3827 6502 7337 6554
rect 7389 6502 7401 6554
rect 7453 6502 7465 6554
rect 7517 6502 7529 6554
rect 7581 6502 7593 6554
rect 7645 6502 11155 6554
rect 11207 6502 11219 6554
rect 11271 6502 11283 6554
rect 11335 6502 11347 6554
rect 11399 6502 11411 6554
rect 11463 6502 14973 6554
rect 15025 6502 15037 6554
rect 15089 6502 15101 6554
rect 15153 6502 15165 6554
rect 15217 6502 15229 6554
rect 15281 6502 16376 6554
rect 1104 6480 16376 6502
rect 1104 6010 16376 6032
rect 1104 5958 2859 6010
rect 2911 5958 2923 6010
rect 2975 5958 2987 6010
rect 3039 5958 3051 6010
rect 3103 5958 3115 6010
rect 3167 5958 6677 6010
rect 6729 5958 6741 6010
rect 6793 5958 6805 6010
rect 6857 5958 6869 6010
rect 6921 5958 6933 6010
rect 6985 5958 10495 6010
rect 10547 5958 10559 6010
rect 10611 5958 10623 6010
rect 10675 5958 10687 6010
rect 10739 5958 10751 6010
rect 10803 5958 14313 6010
rect 14365 5958 14377 6010
rect 14429 5958 14441 6010
rect 14493 5958 14505 6010
rect 14557 5958 14569 6010
rect 14621 5958 16376 6010
rect 1104 5936 16376 5958
rect 1104 5466 16376 5488
rect 1104 5414 3519 5466
rect 3571 5414 3583 5466
rect 3635 5414 3647 5466
rect 3699 5414 3711 5466
rect 3763 5414 3775 5466
rect 3827 5414 7337 5466
rect 7389 5414 7401 5466
rect 7453 5414 7465 5466
rect 7517 5414 7529 5466
rect 7581 5414 7593 5466
rect 7645 5414 11155 5466
rect 11207 5414 11219 5466
rect 11271 5414 11283 5466
rect 11335 5414 11347 5466
rect 11399 5414 11411 5466
rect 11463 5414 14973 5466
rect 15025 5414 15037 5466
rect 15089 5414 15101 5466
rect 15153 5414 15165 5466
rect 15217 5414 15229 5466
rect 15281 5414 16376 5466
rect 1104 5392 16376 5414
rect 5902 5108 5908 5160
rect 5960 5108 5966 5160
rect 8386 5108 8392 5160
rect 8444 5108 8450 5160
rect 5166 4972 5172 5024
rect 5224 5012 5230 5024
rect 5261 5015 5319 5021
rect 5261 5012 5273 5015
rect 5224 4984 5273 5012
rect 5224 4972 5230 4984
rect 5261 4981 5273 4984
rect 5307 4981 5319 5015
rect 5261 4975 5319 4981
rect 7834 4972 7840 5024
rect 7892 4972 7898 5024
rect 1104 4922 16376 4944
rect 1104 4870 2859 4922
rect 2911 4870 2923 4922
rect 2975 4870 2987 4922
rect 3039 4870 3051 4922
rect 3103 4870 3115 4922
rect 3167 4870 6677 4922
rect 6729 4870 6741 4922
rect 6793 4870 6805 4922
rect 6857 4870 6869 4922
rect 6921 4870 6933 4922
rect 6985 4870 10495 4922
rect 10547 4870 10559 4922
rect 10611 4870 10623 4922
rect 10675 4870 10687 4922
rect 10739 4870 10751 4922
rect 10803 4870 14313 4922
rect 14365 4870 14377 4922
rect 14429 4870 14441 4922
rect 14493 4870 14505 4922
rect 14557 4870 14569 4922
rect 14621 4870 16376 4922
rect 1104 4848 16376 4870
rect 7834 4768 7840 4820
rect 7892 4808 7898 4820
rect 7892 4780 8248 4808
rect 7892 4768 7898 4780
rect 6270 4700 6276 4752
rect 6328 4740 6334 4752
rect 6825 4743 6883 4749
rect 6825 4740 6837 4743
rect 6328 4712 6837 4740
rect 6328 4700 6334 4712
rect 6825 4709 6837 4712
rect 6871 4709 6883 4743
rect 6825 4703 6883 4709
rect 4982 4564 4988 4616
rect 5040 4564 5046 4616
rect 7006 4564 7012 4616
rect 7064 4564 7070 4616
rect 8220 4613 8248 4780
rect 8389 4675 8447 4681
rect 8389 4641 8401 4675
rect 8435 4672 8447 4675
rect 9582 4672 9588 4684
rect 8435 4644 9588 4672
rect 8435 4641 8447 4644
rect 8389 4635 8447 4641
rect 8205 4607 8263 4613
rect 8205 4573 8217 4607
rect 8251 4573 8263 4607
rect 8205 4567 8263 4573
rect 5258 4496 5264 4548
rect 5316 4496 5322 4548
rect 5718 4496 5724 4548
rect 5776 4496 5782 4548
rect 8404 4536 8432 4635
rect 9582 4632 9588 4644
rect 9640 4672 9646 4684
rect 10413 4675 10471 4681
rect 10413 4672 10425 4675
rect 9640 4644 10425 4672
rect 9640 4632 9646 4644
rect 10413 4641 10425 4644
rect 10459 4641 10471 4675
rect 10413 4635 10471 4641
rect 10226 4564 10232 4616
rect 10284 4564 10290 4616
rect 6932 4508 8432 4536
rect 6932 4480 6960 4508
rect 5626 4428 5632 4480
rect 5684 4468 5690 4480
rect 6733 4471 6791 4477
rect 6733 4468 6745 4471
rect 5684 4440 6745 4468
rect 5684 4428 5690 4440
rect 6733 4437 6745 4440
rect 6779 4437 6791 4471
rect 6733 4431 6791 4437
rect 6914 4428 6920 4480
rect 6972 4428 6978 4480
rect 7834 4428 7840 4480
rect 7892 4428 7898 4480
rect 8202 4428 8208 4480
rect 8260 4468 8266 4480
rect 8297 4471 8355 4477
rect 8297 4468 8309 4471
rect 8260 4440 8309 4468
rect 8260 4428 8266 4440
rect 8297 4437 8309 4440
rect 8343 4437 8355 4471
rect 8297 4431 8355 4437
rect 9858 4428 9864 4480
rect 9916 4428 9922 4480
rect 10321 4471 10379 4477
rect 10321 4437 10333 4471
rect 10367 4468 10379 4471
rect 11054 4468 11060 4480
rect 10367 4440 11060 4468
rect 10367 4437 10379 4440
rect 10321 4431 10379 4437
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 1104 4378 16376 4400
rect 1104 4326 3519 4378
rect 3571 4326 3583 4378
rect 3635 4326 3647 4378
rect 3699 4326 3711 4378
rect 3763 4326 3775 4378
rect 3827 4326 7337 4378
rect 7389 4326 7401 4378
rect 7453 4326 7465 4378
rect 7517 4326 7529 4378
rect 7581 4326 7593 4378
rect 7645 4326 11155 4378
rect 11207 4326 11219 4378
rect 11271 4326 11283 4378
rect 11335 4326 11347 4378
rect 11399 4326 11411 4378
rect 11463 4326 14973 4378
rect 15025 4326 15037 4378
rect 15089 4326 15101 4378
rect 15153 4326 15165 4378
rect 15217 4326 15229 4378
rect 15281 4326 16376 4378
rect 1104 4304 16376 4326
rect 5166 4224 5172 4276
rect 5224 4224 5230 4276
rect 5258 4224 5264 4276
rect 5316 4224 5322 4276
rect 5626 4224 5632 4276
rect 5684 4224 5690 4276
rect 5902 4224 5908 4276
rect 5960 4264 5966 4276
rect 6089 4267 6147 4273
rect 6089 4264 6101 4267
rect 5960 4236 6101 4264
rect 5960 4224 5966 4236
rect 6089 4233 6101 4236
rect 6135 4233 6147 4267
rect 6089 4227 6147 4233
rect 9858 4224 9864 4276
rect 9916 4224 9922 4276
rect 4798 4088 4804 4140
rect 4856 4088 4862 4140
rect 5077 4131 5135 4137
rect 5077 4097 5089 4131
rect 5123 4128 5135 4131
rect 5184 4128 5212 4224
rect 7282 4156 7288 4208
rect 7340 4156 7346 4208
rect 9876 4196 9904 4224
rect 15470 4196 15476 4208
rect 9416 4168 9904 4196
rect 10902 4182 15476 4196
rect 10888 4168 15476 4182
rect 5123 4100 5212 4128
rect 5721 4131 5779 4137
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 5721 4097 5733 4131
rect 5767 4128 5779 4131
rect 6365 4131 6423 4137
rect 6365 4128 6377 4131
rect 5767 4100 6377 4128
rect 5767 4097 5779 4100
rect 5721 4091 5779 4097
rect 6365 4097 6377 4100
rect 6411 4097 6423 4131
rect 6365 4091 6423 4097
rect 9125 4131 9183 4137
rect 9125 4097 9137 4131
rect 9171 4128 9183 4131
rect 9416 4128 9444 4168
rect 9171 4100 9444 4128
rect 9171 4097 9183 4100
rect 9125 4091 9183 4097
rect 5445 4063 5503 4069
rect 5445 4060 5457 4063
rect 4172 4032 5457 4060
rect 4172 3936 4200 4032
rect 5445 4029 5457 4032
rect 5491 4060 5503 4063
rect 6454 4060 6460 4072
rect 5491 4032 6460 4060
rect 5491 4029 5503 4032
rect 5445 4023 5503 4029
rect 6454 4020 6460 4032
rect 6512 4060 6518 4072
rect 6914 4060 6920 4072
rect 6512 4032 6920 4060
rect 6512 4020 6518 4032
rect 6914 4020 6920 4032
rect 6972 4020 6978 4072
rect 7009 4063 7067 4069
rect 7009 4029 7021 4063
rect 7055 4060 7067 4063
rect 7098 4060 7104 4072
rect 7055 4032 7104 4060
rect 7055 4029 7067 4032
rect 7009 4023 7067 4029
rect 7098 4020 7104 4032
rect 7156 4020 7162 4072
rect 9398 4020 9404 4072
rect 9456 4020 9462 4072
rect 9677 4063 9735 4069
rect 9677 4060 9689 4063
rect 9508 4032 9689 4060
rect 9309 3995 9367 4001
rect 9309 3961 9321 3995
rect 9355 3961 9367 3995
rect 9309 3955 9367 3961
rect 4154 3884 4160 3936
rect 4212 3884 4218 3936
rect 4985 3927 5043 3933
rect 4985 3893 4997 3927
rect 5031 3924 5043 3927
rect 5534 3924 5540 3936
rect 5031 3896 5540 3924
rect 5031 3893 5043 3896
rect 4985 3887 5043 3893
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 6546 3884 6552 3936
rect 6604 3924 6610 3936
rect 8570 3924 8576 3936
rect 6604 3896 8576 3924
rect 6604 3884 6610 3896
rect 8570 3884 8576 3896
rect 8628 3884 8634 3936
rect 9324 3924 9352 3955
rect 9508 3924 9536 4032
rect 9677 4029 9689 4032
rect 9723 4029 9735 4063
rect 9677 4023 9735 4029
rect 10410 4020 10416 4072
rect 10468 4060 10474 4072
rect 10888 4060 10916 4168
rect 15470 4156 15476 4168
rect 15528 4156 15534 4208
rect 10468 4032 10916 4060
rect 10468 4020 10474 4032
rect 9324 3896 9536 3924
rect 11054 3884 11060 3936
rect 11112 3924 11118 3936
rect 11149 3927 11207 3933
rect 11149 3924 11161 3927
rect 11112 3896 11161 3924
rect 11112 3884 11118 3896
rect 11149 3893 11161 3896
rect 11195 3893 11207 3927
rect 11149 3887 11207 3893
rect 1104 3834 16376 3856
rect 1104 3782 2859 3834
rect 2911 3782 2923 3834
rect 2975 3782 2987 3834
rect 3039 3782 3051 3834
rect 3103 3782 3115 3834
rect 3167 3782 6677 3834
rect 6729 3782 6741 3834
rect 6793 3782 6805 3834
rect 6857 3782 6869 3834
rect 6921 3782 6933 3834
rect 6985 3782 10495 3834
rect 10547 3782 10559 3834
rect 10611 3782 10623 3834
rect 10675 3782 10687 3834
rect 10739 3782 10751 3834
rect 10803 3782 14313 3834
rect 14365 3782 14377 3834
rect 14429 3782 14441 3834
rect 14493 3782 14505 3834
rect 14557 3782 14569 3834
rect 14621 3782 16376 3834
rect 1104 3760 16376 3782
rect 4709 3723 4767 3729
rect 4709 3689 4721 3723
rect 4755 3720 4767 3723
rect 4798 3720 4804 3732
rect 4755 3692 4804 3720
rect 4755 3689 4767 3692
rect 4709 3683 4767 3689
rect 4798 3680 4804 3692
rect 4856 3680 4862 3732
rect 4982 3680 4988 3732
rect 5040 3720 5046 3732
rect 5077 3723 5135 3729
rect 5077 3720 5089 3723
rect 5040 3692 5089 3720
rect 5040 3680 5046 3692
rect 5077 3689 5089 3692
rect 5123 3689 5135 3723
rect 5077 3683 5135 3689
rect 2498 3544 2504 3596
rect 2556 3584 2562 3596
rect 4154 3584 4160 3596
rect 2556 3556 4160 3584
rect 2556 3544 2562 3556
rect 4154 3544 4160 3556
rect 4212 3544 4218 3596
rect 5092 3584 5120 3683
rect 8202 3680 8208 3732
rect 8260 3720 8266 3732
rect 8389 3723 8447 3729
rect 8389 3720 8401 3723
rect 8260 3692 8401 3720
rect 8260 3680 8266 3692
rect 8389 3689 8401 3692
rect 8435 3689 8447 3723
rect 8389 3683 8447 3689
rect 8570 3680 8576 3732
rect 8628 3680 8634 3732
rect 9398 3680 9404 3732
rect 9456 3720 9462 3732
rect 10873 3723 10931 3729
rect 10873 3720 10885 3723
rect 9456 3692 10885 3720
rect 9456 3680 9462 3692
rect 10873 3689 10885 3692
rect 10919 3689 10931 3723
rect 10873 3683 10931 3689
rect 6178 3584 6184 3596
rect 5092 3556 6184 3584
rect 6178 3544 6184 3556
rect 6236 3584 6242 3596
rect 6641 3587 6699 3593
rect 6641 3584 6653 3587
rect 6236 3556 6653 3584
rect 6236 3544 6242 3556
rect 6641 3553 6653 3556
rect 6687 3553 6699 3587
rect 8588 3584 8616 3680
rect 8588 3556 9628 3584
rect 6641 3547 6699 3553
rect 4338 3476 4344 3528
rect 4396 3516 4402 3528
rect 5626 3516 5632 3528
rect 4396 3488 5632 3516
rect 4396 3476 4402 3488
rect 5626 3476 5632 3488
rect 5684 3476 5690 3528
rect 6546 3476 6552 3528
rect 6604 3476 6610 3528
rect 8570 3476 8576 3528
rect 8628 3476 8634 3528
rect 9600 3525 9628 3556
rect 9585 3519 9643 3525
rect 9585 3485 9597 3519
rect 9631 3485 9643 3519
rect 9585 3479 9643 3485
rect 10410 3476 10416 3528
rect 10468 3476 10474 3528
rect 11606 3476 11612 3528
rect 11664 3476 11670 3528
rect 6917 3451 6975 3457
rect 6917 3417 6929 3451
rect 6963 3448 6975 3451
rect 7190 3448 7196 3460
rect 6963 3420 7196 3448
rect 6963 3417 6975 3420
rect 6917 3411 6975 3417
rect 7190 3408 7196 3420
rect 7248 3408 7254 3460
rect 10428 3448 10456 3476
rect 8142 3420 10456 3448
rect 4246 3340 4252 3392
rect 4304 3340 4310 3392
rect 6822 3340 6828 3392
rect 6880 3380 6886 3392
rect 8220 3380 8248 3420
rect 6880 3352 8248 3380
rect 6880 3340 6886 3352
rect 8754 3340 8760 3392
rect 8812 3340 8818 3392
rect 10686 3340 10692 3392
rect 10744 3380 10750 3392
rect 11425 3383 11483 3389
rect 11425 3380 11437 3383
rect 10744 3352 11437 3380
rect 10744 3340 10750 3352
rect 11425 3349 11437 3352
rect 11471 3349 11483 3383
rect 11425 3343 11483 3349
rect 1104 3290 16376 3312
rect 1104 3238 3519 3290
rect 3571 3238 3583 3290
rect 3635 3238 3647 3290
rect 3699 3238 3711 3290
rect 3763 3238 3775 3290
rect 3827 3238 7337 3290
rect 7389 3238 7401 3290
rect 7453 3238 7465 3290
rect 7517 3238 7529 3290
rect 7581 3238 7593 3290
rect 7645 3238 11155 3290
rect 11207 3238 11219 3290
rect 11271 3238 11283 3290
rect 11335 3238 11347 3290
rect 11399 3238 11411 3290
rect 11463 3238 14973 3290
rect 15025 3238 15037 3290
rect 15089 3238 15101 3290
rect 15153 3238 15165 3290
rect 15217 3238 15229 3290
rect 15281 3238 16376 3290
rect 1104 3216 16376 3238
rect 4246 3136 4252 3188
rect 4304 3176 4310 3188
rect 4341 3179 4399 3185
rect 4341 3176 4353 3179
rect 4304 3148 4353 3176
rect 4304 3136 4310 3148
rect 4341 3145 4353 3148
rect 4387 3145 4399 3179
rect 4341 3139 4399 3145
rect 4982 3136 4988 3188
rect 5040 3136 5046 3188
rect 6822 3176 6828 3188
rect 5828 3148 6828 3176
rect 5000 3108 5028 3136
rect 4448 3080 5028 3108
rect 4448 3049 4476 3080
rect 4433 3043 4491 3049
rect 4433 3009 4445 3043
rect 4479 3009 4491 3043
rect 4433 3003 4491 3009
rect 5718 3000 5724 3052
rect 5776 3040 5782 3052
rect 5828 3040 5856 3148
rect 6822 3136 6828 3148
rect 6880 3176 6886 3188
rect 6880 3148 7328 3176
rect 6880 3136 6886 3148
rect 6270 3068 6276 3120
rect 6328 3068 6334 3120
rect 6454 3068 6460 3120
rect 6512 3068 6518 3120
rect 6546 3068 6552 3120
rect 6604 3108 6610 3120
rect 6733 3111 6791 3117
rect 6733 3108 6745 3111
rect 6604 3080 6745 3108
rect 6604 3068 6610 3080
rect 6733 3077 6745 3080
rect 6779 3077 6791 3111
rect 7300 3108 7328 3148
rect 9398 3136 9404 3188
rect 9456 3136 9462 3188
rect 10686 3136 10692 3188
rect 10744 3136 10750 3188
rect 9416 3108 9444 3136
rect 7300 3080 7590 3108
rect 9140 3080 9444 3108
rect 6733 3071 6791 3077
rect 5776 3026 5856 3040
rect 5776 3012 5842 3026
rect 5776 3000 5782 3012
rect 3694 2932 3700 2984
rect 3752 2932 3758 2984
rect 4709 2975 4767 2981
rect 4709 2941 4721 2975
rect 4755 2972 4767 2975
rect 6288 2972 6316 3068
rect 4755 2944 6316 2972
rect 6472 2972 6500 3068
rect 9140 3049 9168 3080
rect 10410 3068 10416 3120
rect 10468 3068 10474 3120
rect 6825 3043 6883 3049
rect 6825 3009 6837 3043
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 9033 3043 9091 3049
rect 9033 3009 9045 3043
rect 9079 3040 9091 3043
rect 9125 3043 9183 3049
rect 9125 3040 9137 3043
rect 9079 3012 9137 3040
rect 9079 3009 9091 3012
rect 9033 3003 9091 3009
rect 9125 3009 9137 3012
rect 9171 3009 9183 3043
rect 9125 3003 9183 3009
rect 6549 2975 6607 2981
rect 6549 2972 6561 2975
rect 6472 2944 6561 2972
rect 4755 2941 4767 2944
rect 4709 2935 4767 2941
rect 6549 2941 6561 2944
rect 6595 2941 6607 2975
rect 6840 2972 6868 3003
rect 8202 2972 8208 2984
rect 6840 2944 8208 2972
rect 6549 2935 6607 2941
rect 8202 2932 8208 2944
rect 8260 2932 8266 2984
rect 8754 2932 8760 2984
rect 8812 2932 8818 2984
rect 9401 2975 9459 2981
rect 9401 2941 9413 2975
rect 9447 2972 9459 2975
rect 10704 2972 10732 3136
rect 9447 2944 10732 2972
rect 10873 2975 10931 2981
rect 9447 2941 9459 2944
rect 9401 2935 9459 2941
rect 10873 2941 10885 2975
rect 10919 2972 10931 2975
rect 12066 2972 12072 2984
rect 10919 2944 12072 2972
rect 10919 2941 10931 2944
rect 10873 2935 10931 2941
rect 12066 2932 12072 2944
rect 12124 2932 12130 2984
rect 7006 2864 7012 2916
rect 7064 2904 7070 2916
rect 7193 2907 7251 2913
rect 7193 2904 7205 2907
rect 7064 2876 7205 2904
rect 7064 2864 7070 2876
rect 7193 2873 7205 2876
rect 7239 2873 7251 2907
rect 7193 2867 7251 2873
rect 6181 2839 6239 2845
rect 6181 2805 6193 2839
rect 6227 2836 6239 2839
rect 7098 2836 7104 2848
rect 6227 2808 7104 2836
rect 6227 2805 6239 2808
rect 6181 2799 6239 2805
rect 7098 2796 7104 2808
rect 7156 2796 7162 2848
rect 7285 2839 7343 2845
rect 7285 2805 7297 2839
rect 7331 2836 7343 2839
rect 8386 2836 8392 2848
rect 7331 2808 8392 2836
rect 7331 2805 7343 2808
rect 7285 2799 7343 2805
rect 8386 2796 8392 2808
rect 8444 2796 8450 2848
rect 9766 2796 9772 2848
rect 9824 2836 9830 2848
rect 11054 2836 11060 2848
rect 9824 2808 11060 2836
rect 9824 2796 9830 2808
rect 11054 2796 11060 2808
rect 11112 2796 11118 2848
rect 11514 2796 11520 2848
rect 11572 2796 11578 2848
rect 1104 2746 16376 2768
rect 1104 2694 2859 2746
rect 2911 2694 2923 2746
rect 2975 2694 2987 2746
rect 3039 2694 3051 2746
rect 3103 2694 3115 2746
rect 3167 2694 6677 2746
rect 6729 2694 6741 2746
rect 6793 2694 6805 2746
rect 6857 2694 6869 2746
rect 6921 2694 6933 2746
rect 6985 2694 10495 2746
rect 10547 2694 10559 2746
rect 10611 2694 10623 2746
rect 10675 2694 10687 2746
rect 10739 2694 10751 2746
rect 10803 2694 14313 2746
rect 14365 2694 14377 2746
rect 14429 2694 14441 2746
rect 14493 2694 14505 2746
rect 14557 2694 14569 2746
rect 14621 2694 16376 2746
rect 1104 2672 16376 2694
rect 6546 2592 6552 2644
rect 6604 2592 6610 2644
rect 7190 2592 7196 2644
rect 7248 2632 7254 2644
rect 7285 2635 7343 2641
rect 7285 2632 7297 2635
rect 7248 2604 7297 2632
rect 7248 2592 7254 2604
rect 7285 2601 7297 2604
rect 7331 2601 7343 2635
rect 7285 2595 7343 2601
rect 8570 2592 8576 2644
rect 8628 2632 8634 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 8628 2604 9137 2632
rect 8628 2592 8634 2604
rect 9125 2601 9137 2604
rect 9171 2601 9183 2635
rect 9125 2595 9183 2601
rect 11054 2592 11060 2644
rect 11112 2592 11118 2644
rect 11606 2592 11612 2644
rect 11664 2592 11670 2644
rect 10781 2567 10839 2573
rect 10781 2533 10793 2567
rect 10827 2564 10839 2567
rect 11624 2564 11652 2592
rect 10827 2536 11652 2564
rect 10827 2533 10839 2536
rect 10781 2527 10839 2533
rect 4433 2499 4491 2505
rect 4433 2496 4445 2499
rect 3712 2468 4445 2496
rect 3712 2440 3740 2468
rect 4433 2465 4445 2468
rect 4479 2465 4491 2499
rect 4433 2459 4491 2465
rect 5534 2456 5540 2508
rect 5592 2496 5598 2508
rect 5905 2499 5963 2505
rect 5905 2496 5917 2499
rect 5592 2468 5917 2496
rect 5592 2456 5598 2468
rect 5905 2465 5917 2468
rect 5951 2465 5963 2499
rect 5905 2459 5963 2465
rect 6178 2456 6184 2508
rect 6236 2456 6242 2508
rect 7098 2456 7104 2508
rect 7156 2496 7162 2508
rect 7156 2468 8248 2496
rect 7156 2456 7162 2468
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2428 1823 2431
rect 3694 2428 3700 2440
rect 1811 2400 3700 2428
rect 1811 2397 1823 2400
rect 1765 2391 1823 2397
rect 3694 2388 3700 2400
rect 3752 2388 3758 2440
rect 4157 2431 4215 2437
rect 4157 2397 4169 2431
rect 4203 2428 4215 2431
rect 4338 2428 4344 2440
rect 4203 2400 4344 2428
rect 4203 2397 4215 2400
rect 4157 2391 4215 2397
rect 4338 2388 4344 2400
rect 4396 2388 4402 2440
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2428 7527 2431
rect 7834 2428 7840 2440
rect 7515 2400 7840 2428
rect 7515 2397 7527 2400
rect 7469 2391 7527 2397
rect 7834 2388 7840 2400
rect 7892 2388 7898 2440
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2428 7987 2431
rect 8110 2428 8116 2440
rect 7975 2400 8116 2428
rect 7975 2397 7987 2400
rect 7929 2391 7987 2397
rect 8110 2388 8116 2400
rect 8168 2388 8174 2440
rect 8220 2437 8248 2468
rect 9582 2456 9588 2508
rect 9640 2496 9646 2508
rect 9677 2499 9735 2505
rect 9677 2496 9689 2499
rect 9640 2468 9689 2496
rect 9640 2456 9646 2468
rect 9677 2465 9689 2468
rect 9723 2496 9735 2499
rect 10137 2499 10195 2505
rect 10137 2496 10149 2499
rect 9723 2468 10149 2496
rect 9723 2465 9735 2468
rect 9677 2459 9735 2465
rect 10137 2465 10149 2468
rect 10183 2465 10195 2499
rect 10137 2459 10195 2465
rect 10321 2499 10379 2505
rect 10321 2465 10333 2499
rect 10367 2496 10379 2499
rect 11514 2496 11520 2508
rect 10367 2468 11520 2496
rect 10367 2465 10379 2468
rect 10321 2459 10379 2465
rect 8205 2431 8263 2437
rect 8205 2397 8217 2431
rect 8251 2397 8263 2431
rect 8205 2391 8263 2397
rect 9493 2431 9551 2437
rect 9493 2397 9505 2431
rect 9539 2428 9551 2431
rect 10336 2428 10364 2459
rect 11514 2456 11520 2468
rect 11572 2456 11578 2508
rect 9539 2400 10364 2428
rect 10413 2431 10471 2437
rect 9539 2397 9551 2400
rect 9493 2391 9551 2397
rect 10413 2397 10425 2431
rect 10459 2428 10471 2431
rect 11146 2428 11152 2440
rect 10459 2400 11152 2428
rect 10459 2397 10471 2400
rect 10413 2391 10471 2397
rect 11146 2388 11152 2400
rect 11204 2428 11210 2440
rect 11204 2400 11560 2428
rect 11204 2388 11210 2400
rect 1302 2320 1308 2372
rect 1360 2360 1366 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 1360 2332 1409 2360
rect 1360 2320 1366 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 1397 2323 1455 2329
rect 3418 2320 3424 2372
rect 3476 2360 3482 2372
rect 3789 2363 3847 2369
rect 3789 2360 3801 2363
rect 3476 2332 3801 2360
rect 3476 2320 3482 2332
rect 3789 2329 3801 2332
rect 3835 2329 3847 2363
rect 5474 2332 5580 2360
rect 3789 2323 3847 2329
rect 5552 2292 5580 2332
rect 5626 2320 5632 2372
rect 5684 2360 5690 2372
rect 10965 2363 11023 2369
rect 10965 2360 10977 2363
rect 5684 2332 7788 2360
rect 5684 2320 5690 2332
rect 5718 2292 5724 2304
rect 5552 2264 5724 2292
rect 5718 2252 5724 2264
rect 5776 2252 5782 2304
rect 7650 2252 7656 2304
rect 7708 2252 7714 2304
rect 7760 2292 7788 2332
rect 9600 2332 10977 2360
rect 8297 2295 8355 2301
rect 8297 2292 8309 2295
rect 7760 2264 8309 2292
rect 8297 2261 8309 2264
rect 8343 2261 8355 2295
rect 8297 2255 8355 2261
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 9600 2301 9628 2332
rect 10965 2329 10977 2332
rect 11011 2329 11023 2363
rect 11532 2360 11560 2400
rect 12066 2388 12072 2440
rect 12124 2388 12130 2440
rect 16022 2388 16028 2440
rect 16080 2388 16086 2440
rect 14185 2363 14243 2369
rect 14185 2360 14197 2363
rect 11532 2332 14197 2360
rect 10965 2323 11023 2329
rect 14185 2329 14197 2332
rect 14231 2329 14243 2363
rect 14185 2323 14243 2329
rect 9585 2295 9643 2301
rect 9585 2292 9597 2295
rect 8444 2264 9597 2292
rect 8444 2252 8450 2264
rect 9585 2261 9597 2264
rect 9631 2261 9643 2295
rect 9585 2255 9643 2261
rect 11882 2252 11888 2304
rect 11940 2292 11946 2304
rect 12161 2295 12219 2301
rect 12161 2292 12173 2295
rect 11940 2264 12173 2292
rect 11940 2252 11946 2264
rect 12161 2261 12173 2264
rect 12207 2261 12219 2295
rect 12161 2255 12219 2261
rect 13998 2252 14004 2304
rect 14056 2292 14062 2304
rect 14277 2295 14335 2301
rect 14277 2292 14289 2295
rect 14056 2264 14289 2292
rect 14056 2252 14062 2264
rect 14277 2261 14289 2264
rect 14323 2261 14335 2295
rect 14277 2255 14335 2261
rect 1104 2202 16376 2224
rect 1104 2150 3519 2202
rect 3571 2150 3583 2202
rect 3635 2150 3647 2202
rect 3699 2150 3711 2202
rect 3763 2150 3775 2202
rect 3827 2150 7337 2202
rect 7389 2150 7401 2202
rect 7453 2150 7465 2202
rect 7517 2150 7529 2202
rect 7581 2150 7593 2202
rect 7645 2150 11155 2202
rect 11207 2150 11219 2202
rect 11271 2150 11283 2202
rect 11335 2150 11347 2202
rect 11399 2150 11411 2202
rect 11463 2150 14973 2202
rect 15025 2150 15037 2202
rect 15089 2150 15101 2202
rect 15153 2150 15165 2202
rect 15217 2150 15229 2202
rect 15281 2150 16376 2202
rect 1104 2128 16376 2150
<< via1 >>
rect 3519 17382 3571 17434
rect 3583 17382 3635 17434
rect 3647 17382 3699 17434
rect 3711 17382 3763 17434
rect 3775 17382 3827 17434
rect 7337 17382 7389 17434
rect 7401 17382 7453 17434
rect 7465 17382 7517 17434
rect 7529 17382 7581 17434
rect 7593 17382 7645 17434
rect 11155 17382 11207 17434
rect 11219 17382 11271 17434
rect 11283 17382 11335 17434
rect 11347 17382 11399 17434
rect 11411 17382 11463 17434
rect 14973 17382 15025 17434
rect 15037 17382 15089 17434
rect 15101 17382 15153 17434
rect 15165 17382 15217 17434
rect 15229 17382 15281 17434
rect 11060 17280 11112 17332
rect 2228 17212 2280 17264
rect 15384 17255 15436 17264
rect 15384 17221 15393 17255
rect 15393 17221 15427 17255
rect 15427 17221 15436 17255
rect 15384 17212 15436 17221
rect 2504 16983 2556 16992
rect 2504 16949 2513 16983
rect 2513 16949 2547 16983
rect 2547 16949 2556 16983
rect 2504 16940 2556 16949
rect 10232 16940 10284 16992
rect 15476 16983 15528 16992
rect 15476 16949 15485 16983
rect 15485 16949 15519 16983
rect 15519 16949 15528 16983
rect 15476 16940 15528 16949
rect 2859 16838 2911 16890
rect 2923 16838 2975 16890
rect 2987 16838 3039 16890
rect 3051 16838 3103 16890
rect 3115 16838 3167 16890
rect 6677 16838 6729 16890
rect 6741 16838 6793 16890
rect 6805 16838 6857 16890
rect 6869 16838 6921 16890
rect 6933 16838 6985 16890
rect 10495 16838 10547 16890
rect 10559 16838 10611 16890
rect 10623 16838 10675 16890
rect 10687 16838 10739 16890
rect 10751 16838 10803 16890
rect 14313 16838 14365 16890
rect 14377 16838 14429 16890
rect 14441 16838 14493 16890
rect 14505 16838 14557 16890
rect 14569 16838 14621 16890
rect 3519 16294 3571 16346
rect 3583 16294 3635 16346
rect 3647 16294 3699 16346
rect 3711 16294 3763 16346
rect 3775 16294 3827 16346
rect 7337 16294 7389 16346
rect 7401 16294 7453 16346
rect 7465 16294 7517 16346
rect 7529 16294 7581 16346
rect 7593 16294 7645 16346
rect 11155 16294 11207 16346
rect 11219 16294 11271 16346
rect 11283 16294 11335 16346
rect 11347 16294 11399 16346
rect 11411 16294 11463 16346
rect 14973 16294 15025 16346
rect 15037 16294 15089 16346
rect 15101 16294 15153 16346
rect 15165 16294 15217 16346
rect 15229 16294 15281 16346
rect 2859 15750 2911 15802
rect 2923 15750 2975 15802
rect 2987 15750 3039 15802
rect 3051 15750 3103 15802
rect 3115 15750 3167 15802
rect 6677 15750 6729 15802
rect 6741 15750 6793 15802
rect 6805 15750 6857 15802
rect 6869 15750 6921 15802
rect 6933 15750 6985 15802
rect 10495 15750 10547 15802
rect 10559 15750 10611 15802
rect 10623 15750 10675 15802
rect 10687 15750 10739 15802
rect 10751 15750 10803 15802
rect 14313 15750 14365 15802
rect 14377 15750 14429 15802
rect 14441 15750 14493 15802
rect 14505 15750 14557 15802
rect 14569 15750 14621 15802
rect 6552 15308 6604 15360
rect 7196 15308 7248 15360
rect 3519 15206 3571 15258
rect 3583 15206 3635 15258
rect 3647 15206 3699 15258
rect 3711 15206 3763 15258
rect 3775 15206 3827 15258
rect 7337 15206 7389 15258
rect 7401 15206 7453 15258
rect 7465 15206 7517 15258
rect 7529 15206 7581 15258
rect 7593 15206 7645 15258
rect 11155 15206 11207 15258
rect 11219 15206 11271 15258
rect 11283 15206 11335 15258
rect 11347 15206 11399 15258
rect 11411 15206 11463 15258
rect 14973 15206 15025 15258
rect 15037 15206 15089 15258
rect 15101 15206 15153 15258
rect 15165 15206 15217 15258
rect 15229 15206 15281 15258
rect 2859 14662 2911 14714
rect 2923 14662 2975 14714
rect 2987 14662 3039 14714
rect 3051 14662 3103 14714
rect 3115 14662 3167 14714
rect 6677 14662 6729 14714
rect 6741 14662 6793 14714
rect 6805 14662 6857 14714
rect 6869 14662 6921 14714
rect 6933 14662 6985 14714
rect 10495 14662 10547 14714
rect 10559 14662 10611 14714
rect 10623 14662 10675 14714
rect 10687 14662 10739 14714
rect 10751 14662 10803 14714
rect 14313 14662 14365 14714
rect 14377 14662 14429 14714
rect 14441 14662 14493 14714
rect 14505 14662 14557 14714
rect 14569 14662 14621 14714
rect 3519 14118 3571 14170
rect 3583 14118 3635 14170
rect 3647 14118 3699 14170
rect 3711 14118 3763 14170
rect 3775 14118 3827 14170
rect 7337 14118 7389 14170
rect 7401 14118 7453 14170
rect 7465 14118 7517 14170
rect 7529 14118 7581 14170
rect 7593 14118 7645 14170
rect 11155 14118 11207 14170
rect 11219 14118 11271 14170
rect 11283 14118 11335 14170
rect 11347 14118 11399 14170
rect 11411 14118 11463 14170
rect 14973 14118 15025 14170
rect 15037 14118 15089 14170
rect 15101 14118 15153 14170
rect 15165 14118 15217 14170
rect 15229 14118 15281 14170
rect 2859 13574 2911 13626
rect 2923 13574 2975 13626
rect 2987 13574 3039 13626
rect 3051 13574 3103 13626
rect 3115 13574 3167 13626
rect 6677 13574 6729 13626
rect 6741 13574 6793 13626
rect 6805 13574 6857 13626
rect 6869 13574 6921 13626
rect 6933 13574 6985 13626
rect 10495 13574 10547 13626
rect 10559 13574 10611 13626
rect 10623 13574 10675 13626
rect 10687 13574 10739 13626
rect 10751 13574 10803 13626
rect 14313 13574 14365 13626
rect 14377 13574 14429 13626
rect 14441 13574 14493 13626
rect 14505 13574 14557 13626
rect 14569 13574 14621 13626
rect 3519 13030 3571 13082
rect 3583 13030 3635 13082
rect 3647 13030 3699 13082
rect 3711 13030 3763 13082
rect 3775 13030 3827 13082
rect 7337 13030 7389 13082
rect 7401 13030 7453 13082
rect 7465 13030 7517 13082
rect 7529 13030 7581 13082
rect 7593 13030 7645 13082
rect 11155 13030 11207 13082
rect 11219 13030 11271 13082
rect 11283 13030 11335 13082
rect 11347 13030 11399 13082
rect 11411 13030 11463 13082
rect 14973 13030 15025 13082
rect 15037 13030 15089 13082
rect 15101 13030 15153 13082
rect 15165 13030 15217 13082
rect 15229 13030 15281 13082
rect 2859 12486 2911 12538
rect 2923 12486 2975 12538
rect 2987 12486 3039 12538
rect 3051 12486 3103 12538
rect 3115 12486 3167 12538
rect 6677 12486 6729 12538
rect 6741 12486 6793 12538
rect 6805 12486 6857 12538
rect 6869 12486 6921 12538
rect 6933 12486 6985 12538
rect 10495 12486 10547 12538
rect 10559 12486 10611 12538
rect 10623 12486 10675 12538
rect 10687 12486 10739 12538
rect 10751 12486 10803 12538
rect 14313 12486 14365 12538
rect 14377 12486 14429 12538
rect 14441 12486 14493 12538
rect 14505 12486 14557 12538
rect 14569 12486 14621 12538
rect 3519 11942 3571 11994
rect 3583 11942 3635 11994
rect 3647 11942 3699 11994
rect 3711 11942 3763 11994
rect 3775 11942 3827 11994
rect 7337 11942 7389 11994
rect 7401 11942 7453 11994
rect 7465 11942 7517 11994
rect 7529 11942 7581 11994
rect 7593 11942 7645 11994
rect 11155 11942 11207 11994
rect 11219 11942 11271 11994
rect 11283 11942 11335 11994
rect 11347 11942 11399 11994
rect 11411 11942 11463 11994
rect 14973 11942 15025 11994
rect 15037 11942 15089 11994
rect 15101 11942 15153 11994
rect 15165 11942 15217 11994
rect 15229 11942 15281 11994
rect 2859 11398 2911 11450
rect 2923 11398 2975 11450
rect 2987 11398 3039 11450
rect 3051 11398 3103 11450
rect 3115 11398 3167 11450
rect 6677 11398 6729 11450
rect 6741 11398 6793 11450
rect 6805 11398 6857 11450
rect 6869 11398 6921 11450
rect 6933 11398 6985 11450
rect 10495 11398 10547 11450
rect 10559 11398 10611 11450
rect 10623 11398 10675 11450
rect 10687 11398 10739 11450
rect 10751 11398 10803 11450
rect 14313 11398 14365 11450
rect 14377 11398 14429 11450
rect 14441 11398 14493 11450
rect 14505 11398 14557 11450
rect 14569 11398 14621 11450
rect 3519 10854 3571 10906
rect 3583 10854 3635 10906
rect 3647 10854 3699 10906
rect 3711 10854 3763 10906
rect 3775 10854 3827 10906
rect 7337 10854 7389 10906
rect 7401 10854 7453 10906
rect 7465 10854 7517 10906
rect 7529 10854 7581 10906
rect 7593 10854 7645 10906
rect 11155 10854 11207 10906
rect 11219 10854 11271 10906
rect 11283 10854 11335 10906
rect 11347 10854 11399 10906
rect 11411 10854 11463 10906
rect 14973 10854 15025 10906
rect 15037 10854 15089 10906
rect 15101 10854 15153 10906
rect 15165 10854 15217 10906
rect 15229 10854 15281 10906
rect 2859 10310 2911 10362
rect 2923 10310 2975 10362
rect 2987 10310 3039 10362
rect 3051 10310 3103 10362
rect 3115 10310 3167 10362
rect 6677 10310 6729 10362
rect 6741 10310 6793 10362
rect 6805 10310 6857 10362
rect 6869 10310 6921 10362
rect 6933 10310 6985 10362
rect 10495 10310 10547 10362
rect 10559 10310 10611 10362
rect 10623 10310 10675 10362
rect 10687 10310 10739 10362
rect 10751 10310 10803 10362
rect 14313 10310 14365 10362
rect 14377 10310 14429 10362
rect 14441 10310 14493 10362
rect 14505 10310 14557 10362
rect 14569 10310 14621 10362
rect 3519 9766 3571 9818
rect 3583 9766 3635 9818
rect 3647 9766 3699 9818
rect 3711 9766 3763 9818
rect 3775 9766 3827 9818
rect 7337 9766 7389 9818
rect 7401 9766 7453 9818
rect 7465 9766 7517 9818
rect 7529 9766 7581 9818
rect 7593 9766 7645 9818
rect 11155 9766 11207 9818
rect 11219 9766 11271 9818
rect 11283 9766 11335 9818
rect 11347 9766 11399 9818
rect 11411 9766 11463 9818
rect 14973 9766 15025 9818
rect 15037 9766 15089 9818
rect 15101 9766 15153 9818
rect 15165 9766 15217 9818
rect 15229 9766 15281 9818
rect 2859 9222 2911 9274
rect 2923 9222 2975 9274
rect 2987 9222 3039 9274
rect 3051 9222 3103 9274
rect 3115 9222 3167 9274
rect 6677 9222 6729 9274
rect 6741 9222 6793 9274
rect 6805 9222 6857 9274
rect 6869 9222 6921 9274
rect 6933 9222 6985 9274
rect 10495 9222 10547 9274
rect 10559 9222 10611 9274
rect 10623 9222 10675 9274
rect 10687 9222 10739 9274
rect 10751 9222 10803 9274
rect 14313 9222 14365 9274
rect 14377 9222 14429 9274
rect 14441 9222 14493 9274
rect 14505 9222 14557 9274
rect 14569 9222 14621 9274
rect 3519 8678 3571 8730
rect 3583 8678 3635 8730
rect 3647 8678 3699 8730
rect 3711 8678 3763 8730
rect 3775 8678 3827 8730
rect 7337 8678 7389 8730
rect 7401 8678 7453 8730
rect 7465 8678 7517 8730
rect 7529 8678 7581 8730
rect 7593 8678 7645 8730
rect 11155 8678 11207 8730
rect 11219 8678 11271 8730
rect 11283 8678 11335 8730
rect 11347 8678 11399 8730
rect 11411 8678 11463 8730
rect 14973 8678 15025 8730
rect 15037 8678 15089 8730
rect 15101 8678 15153 8730
rect 15165 8678 15217 8730
rect 15229 8678 15281 8730
rect 2859 8134 2911 8186
rect 2923 8134 2975 8186
rect 2987 8134 3039 8186
rect 3051 8134 3103 8186
rect 3115 8134 3167 8186
rect 6677 8134 6729 8186
rect 6741 8134 6793 8186
rect 6805 8134 6857 8186
rect 6869 8134 6921 8186
rect 6933 8134 6985 8186
rect 10495 8134 10547 8186
rect 10559 8134 10611 8186
rect 10623 8134 10675 8186
rect 10687 8134 10739 8186
rect 10751 8134 10803 8186
rect 14313 8134 14365 8186
rect 14377 8134 14429 8186
rect 14441 8134 14493 8186
rect 14505 8134 14557 8186
rect 14569 8134 14621 8186
rect 3519 7590 3571 7642
rect 3583 7590 3635 7642
rect 3647 7590 3699 7642
rect 3711 7590 3763 7642
rect 3775 7590 3827 7642
rect 7337 7590 7389 7642
rect 7401 7590 7453 7642
rect 7465 7590 7517 7642
rect 7529 7590 7581 7642
rect 7593 7590 7645 7642
rect 11155 7590 11207 7642
rect 11219 7590 11271 7642
rect 11283 7590 11335 7642
rect 11347 7590 11399 7642
rect 11411 7590 11463 7642
rect 14973 7590 15025 7642
rect 15037 7590 15089 7642
rect 15101 7590 15153 7642
rect 15165 7590 15217 7642
rect 15229 7590 15281 7642
rect 2859 7046 2911 7098
rect 2923 7046 2975 7098
rect 2987 7046 3039 7098
rect 3051 7046 3103 7098
rect 3115 7046 3167 7098
rect 6677 7046 6729 7098
rect 6741 7046 6793 7098
rect 6805 7046 6857 7098
rect 6869 7046 6921 7098
rect 6933 7046 6985 7098
rect 10495 7046 10547 7098
rect 10559 7046 10611 7098
rect 10623 7046 10675 7098
rect 10687 7046 10739 7098
rect 10751 7046 10803 7098
rect 14313 7046 14365 7098
rect 14377 7046 14429 7098
rect 14441 7046 14493 7098
rect 14505 7046 14557 7098
rect 14569 7046 14621 7098
rect 3519 6502 3571 6554
rect 3583 6502 3635 6554
rect 3647 6502 3699 6554
rect 3711 6502 3763 6554
rect 3775 6502 3827 6554
rect 7337 6502 7389 6554
rect 7401 6502 7453 6554
rect 7465 6502 7517 6554
rect 7529 6502 7581 6554
rect 7593 6502 7645 6554
rect 11155 6502 11207 6554
rect 11219 6502 11271 6554
rect 11283 6502 11335 6554
rect 11347 6502 11399 6554
rect 11411 6502 11463 6554
rect 14973 6502 15025 6554
rect 15037 6502 15089 6554
rect 15101 6502 15153 6554
rect 15165 6502 15217 6554
rect 15229 6502 15281 6554
rect 2859 5958 2911 6010
rect 2923 5958 2975 6010
rect 2987 5958 3039 6010
rect 3051 5958 3103 6010
rect 3115 5958 3167 6010
rect 6677 5958 6729 6010
rect 6741 5958 6793 6010
rect 6805 5958 6857 6010
rect 6869 5958 6921 6010
rect 6933 5958 6985 6010
rect 10495 5958 10547 6010
rect 10559 5958 10611 6010
rect 10623 5958 10675 6010
rect 10687 5958 10739 6010
rect 10751 5958 10803 6010
rect 14313 5958 14365 6010
rect 14377 5958 14429 6010
rect 14441 5958 14493 6010
rect 14505 5958 14557 6010
rect 14569 5958 14621 6010
rect 3519 5414 3571 5466
rect 3583 5414 3635 5466
rect 3647 5414 3699 5466
rect 3711 5414 3763 5466
rect 3775 5414 3827 5466
rect 7337 5414 7389 5466
rect 7401 5414 7453 5466
rect 7465 5414 7517 5466
rect 7529 5414 7581 5466
rect 7593 5414 7645 5466
rect 11155 5414 11207 5466
rect 11219 5414 11271 5466
rect 11283 5414 11335 5466
rect 11347 5414 11399 5466
rect 11411 5414 11463 5466
rect 14973 5414 15025 5466
rect 15037 5414 15089 5466
rect 15101 5414 15153 5466
rect 15165 5414 15217 5466
rect 15229 5414 15281 5466
rect 5908 5151 5960 5160
rect 5908 5117 5917 5151
rect 5917 5117 5951 5151
rect 5951 5117 5960 5151
rect 5908 5108 5960 5117
rect 8392 5151 8444 5160
rect 8392 5117 8401 5151
rect 8401 5117 8435 5151
rect 8435 5117 8444 5151
rect 8392 5108 8444 5117
rect 5172 4972 5224 5024
rect 7840 5015 7892 5024
rect 7840 4981 7849 5015
rect 7849 4981 7883 5015
rect 7883 4981 7892 5015
rect 7840 4972 7892 4981
rect 2859 4870 2911 4922
rect 2923 4870 2975 4922
rect 2987 4870 3039 4922
rect 3051 4870 3103 4922
rect 3115 4870 3167 4922
rect 6677 4870 6729 4922
rect 6741 4870 6793 4922
rect 6805 4870 6857 4922
rect 6869 4870 6921 4922
rect 6933 4870 6985 4922
rect 10495 4870 10547 4922
rect 10559 4870 10611 4922
rect 10623 4870 10675 4922
rect 10687 4870 10739 4922
rect 10751 4870 10803 4922
rect 14313 4870 14365 4922
rect 14377 4870 14429 4922
rect 14441 4870 14493 4922
rect 14505 4870 14557 4922
rect 14569 4870 14621 4922
rect 7840 4768 7892 4820
rect 6276 4700 6328 4752
rect 4988 4607 5040 4616
rect 4988 4573 4997 4607
rect 4997 4573 5031 4607
rect 5031 4573 5040 4607
rect 4988 4564 5040 4573
rect 7012 4607 7064 4616
rect 7012 4573 7021 4607
rect 7021 4573 7055 4607
rect 7055 4573 7064 4607
rect 7012 4564 7064 4573
rect 5264 4539 5316 4548
rect 5264 4505 5273 4539
rect 5273 4505 5307 4539
rect 5307 4505 5316 4539
rect 5264 4496 5316 4505
rect 5724 4496 5776 4548
rect 9588 4632 9640 4684
rect 10232 4607 10284 4616
rect 10232 4573 10241 4607
rect 10241 4573 10275 4607
rect 10275 4573 10284 4607
rect 10232 4564 10284 4573
rect 5632 4428 5684 4480
rect 6920 4428 6972 4480
rect 7840 4471 7892 4480
rect 7840 4437 7849 4471
rect 7849 4437 7883 4471
rect 7883 4437 7892 4471
rect 7840 4428 7892 4437
rect 8208 4428 8260 4480
rect 9864 4471 9916 4480
rect 9864 4437 9873 4471
rect 9873 4437 9907 4471
rect 9907 4437 9916 4471
rect 9864 4428 9916 4437
rect 11060 4428 11112 4480
rect 3519 4326 3571 4378
rect 3583 4326 3635 4378
rect 3647 4326 3699 4378
rect 3711 4326 3763 4378
rect 3775 4326 3827 4378
rect 7337 4326 7389 4378
rect 7401 4326 7453 4378
rect 7465 4326 7517 4378
rect 7529 4326 7581 4378
rect 7593 4326 7645 4378
rect 11155 4326 11207 4378
rect 11219 4326 11271 4378
rect 11283 4326 11335 4378
rect 11347 4326 11399 4378
rect 11411 4326 11463 4378
rect 14973 4326 15025 4378
rect 15037 4326 15089 4378
rect 15101 4326 15153 4378
rect 15165 4326 15217 4378
rect 15229 4326 15281 4378
rect 5172 4224 5224 4276
rect 5264 4267 5316 4276
rect 5264 4233 5273 4267
rect 5273 4233 5307 4267
rect 5307 4233 5316 4267
rect 5264 4224 5316 4233
rect 5632 4267 5684 4276
rect 5632 4233 5641 4267
rect 5641 4233 5675 4267
rect 5675 4233 5684 4267
rect 5632 4224 5684 4233
rect 5908 4224 5960 4276
rect 9864 4224 9916 4276
rect 4804 4131 4856 4140
rect 4804 4097 4813 4131
rect 4813 4097 4847 4131
rect 4847 4097 4856 4131
rect 4804 4088 4856 4097
rect 7288 4199 7340 4208
rect 7288 4165 7297 4199
rect 7297 4165 7331 4199
rect 7331 4165 7340 4199
rect 7288 4156 7340 4165
rect 6460 4020 6512 4072
rect 6920 4020 6972 4072
rect 7104 4020 7156 4072
rect 9404 4063 9456 4072
rect 9404 4029 9413 4063
rect 9413 4029 9447 4063
rect 9447 4029 9456 4063
rect 9404 4020 9456 4029
rect 4160 3884 4212 3936
rect 5540 3884 5592 3936
rect 6552 3884 6604 3936
rect 8576 3927 8628 3936
rect 8576 3893 8585 3927
rect 8585 3893 8619 3927
rect 8619 3893 8628 3927
rect 8576 3884 8628 3893
rect 10416 4020 10468 4072
rect 15476 4156 15528 4208
rect 11060 3884 11112 3936
rect 2859 3782 2911 3834
rect 2923 3782 2975 3834
rect 2987 3782 3039 3834
rect 3051 3782 3103 3834
rect 3115 3782 3167 3834
rect 6677 3782 6729 3834
rect 6741 3782 6793 3834
rect 6805 3782 6857 3834
rect 6869 3782 6921 3834
rect 6933 3782 6985 3834
rect 10495 3782 10547 3834
rect 10559 3782 10611 3834
rect 10623 3782 10675 3834
rect 10687 3782 10739 3834
rect 10751 3782 10803 3834
rect 14313 3782 14365 3834
rect 14377 3782 14429 3834
rect 14441 3782 14493 3834
rect 14505 3782 14557 3834
rect 14569 3782 14621 3834
rect 4804 3680 4856 3732
rect 4988 3680 5040 3732
rect 2504 3544 2556 3596
rect 4160 3587 4212 3596
rect 4160 3553 4169 3587
rect 4169 3553 4203 3587
rect 4203 3553 4212 3587
rect 4160 3544 4212 3553
rect 8208 3680 8260 3732
rect 8576 3680 8628 3732
rect 9404 3680 9456 3732
rect 6184 3544 6236 3596
rect 4344 3519 4396 3528
rect 4344 3485 4353 3519
rect 4353 3485 4387 3519
rect 4387 3485 4396 3519
rect 4344 3476 4396 3485
rect 5632 3476 5684 3528
rect 6552 3519 6604 3528
rect 6552 3485 6561 3519
rect 6561 3485 6595 3519
rect 6595 3485 6604 3519
rect 6552 3476 6604 3485
rect 8576 3519 8628 3528
rect 8576 3485 8585 3519
rect 8585 3485 8619 3519
rect 8619 3485 8628 3519
rect 8576 3476 8628 3485
rect 10416 3476 10468 3528
rect 11612 3519 11664 3528
rect 11612 3485 11621 3519
rect 11621 3485 11655 3519
rect 11655 3485 11664 3519
rect 11612 3476 11664 3485
rect 7196 3408 7248 3460
rect 4252 3383 4304 3392
rect 4252 3349 4261 3383
rect 4261 3349 4295 3383
rect 4295 3349 4304 3383
rect 4252 3340 4304 3349
rect 6828 3340 6880 3392
rect 8760 3383 8812 3392
rect 8760 3349 8769 3383
rect 8769 3349 8803 3383
rect 8803 3349 8812 3383
rect 8760 3340 8812 3349
rect 10692 3340 10744 3392
rect 3519 3238 3571 3290
rect 3583 3238 3635 3290
rect 3647 3238 3699 3290
rect 3711 3238 3763 3290
rect 3775 3238 3827 3290
rect 7337 3238 7389 3290
rect 7401 3238 7453 3290
rect 7465 3238 7517 3290
rect 7529 3238 7581 3290
rect 7593 3238 7645 3290
rect 11155 3238 11207 3290
rect 11219 3238 11271 3290
rect 11283 3238 11335 3290
rect 11347 3238 11399 3290
rect 11411 3238 11463 3290
rect 14973 3238 15025 3290
rect 15037 3238 15089 3290
rect 15101 3238 15153 3290
rect 15165 3238 15217 3290
rect 15229 3238 15281 3290
rect 4252 3136 4304 3188
rect 4988 3136 5040 3188
rect 5724 3000 5776 3052
rect 6828 3136 6880 3188
rect 6276 3068 6328 3120
rect 6460 3068 6512 3120
rect 6552 3068 6604 3120
rect 9404 3136 9456 3188
rect 10692 3136 10744 3188
rect 3700 2975 3752 2984
rect 3700 2941 3709 2975
rect 3709 2941 3743 2975
rect 3743 2941 3752 2975
rect 3700 2932 3752 2941
rect 10416 3068 10468 3120
rect 8208 2932 8260 2984
rect 8760 2975 8812 2984
rect 8760 2941 8769 2975
rect 8769 2941 8803 2975
rect 8803 2941 8812 2975
rect 8760 2932 8812 2941
rect 12072 2975 12124 2984
rect 12072 2941 12081 2975
rect 12081 2941 12115 2975
rect 12115 2941 12124 2975
rect 12072 2932 12124 2941
rect 7012 2864 7064 2916
rect 7104 2796 7156 2848
rect 8392 2796 8444 2848
rect 9772 2796 9824 2848
rect 11060 2796 11112 2848
rect 11520 2839 11572 2848
rect 11520 2805 11529 2839
rect 11529 2805 11563 2839
rect 11563 2805 11572 2839
rect 11520 2796 11572 2805
rect 2859 2694 2911 2746
rect 2923 2694 2975 2746
rect 2987 2694 3039 2746
rect 3051 2694 3103 2746
rect 3115 2694 3167 2746
rect 6677 2694 6729 2746
rect 6741 2694 6793 2746
rect 6805 2694 6857 2746
rect 6869 2694 6921 2746
rect 6933 2694 6985 2746
rect 10495 2694 10547 2746
rect 10559 2694 10611 2746
rect 10623 2694 10675 2746
rect 10687 2694 10739 2746
rect 10751 2694 10803 2746
rect 14313 2694 14365 2746
rect 14377 2694 14429 2746
rect 14441 2694 14493 2746
rect 14505 2694 14557 2746
rect 14569 2694 14621 2746
rect 6552 2635 6604 2644
rect 6552 2601 6561 2635
rect 6561 2601 6595 2635
rect 6595 2601 6604 2635
rect 6552 2592 6604 2601
rect 7196 2592 7248 2644
rect 8576 2592 8628 2644
rect 11060 2635 11112 2644
rect 11060 2601 11069 2635
rect 11069 2601 11103 2635
rect 11103 2601 11112 2635
rect 11060 2592 11112 2601
rect 11612 2592 11664 2644
rect 5540 2456 5592 2508
rect 6184 2499 6236 2508
rect 6184 2465 6193 2499
rect 6193 2465 6227 2499
rect 6227 2465 6236 2499
rect 6184 2456 6236 2465
rect 7104 2499 7156 2508
rect 7104 2465 7113 2499
rect 7113 2465 7147 2499
rect 7147 2465 7156 2499
rect 7104 2456 7156 2465
rect 3700 2388 3752 2440
rect 4344 2388 4396 2440
rect 7840 2388 7892 2440
rect 8116 2388 8168 2440
rect 9588 2456 9640 2508
rect 11520 2456 11572 2508
rect 11152 2388 11204 2440
rect 1308 2320 1360 2372
rect 3424 2320 3476 2372
rect 5632 2320 5684 2372
rect 5724 2252 5776 2304
rect 7656 2295 7708 2304
rect 7656 2261 7665 2295
rect 7665 2261 7699 2295
rect 7699 2261 7708 2295
rect 7656 2252 7708 2261
rect 8392 2252 8444 2304
rect 12072 2431 12124 2440
rect 12072 2397 12081 2431
rect 12081 2397 12115 2431
rect 12115 2397 12124 2431
rect 12072 2388 12124 2397
rect 16028 2431 16080 2440
rect 16028 2397 16037 2431
rect 16037 2397 16071 2431
rect 16071 2397 16080 2431
rect 16028 2388 16080 2397
rect 11888 2252 11940 2304
rect 14004 2252 14056 2304
rect 3519 2150 3571 2202
rect 3583 2150 3635 2202
rect 3647 2150 3699 2202
rect 3711 2150 3763 2202
rect 3775 2150 3827 2202
rect 7337 2150 7389 2202
rect 7401 2150 7453 2202
rect 7465 2150 7517 2202
rect 7529 2150 7581 2202
rect 7593 2150 7645 2202
rect 11155 2150 11207 2202
rect 11219 2150 11271 2202
rect 11283 2150 11335 2202
rect 11347 2150 11399 2202
rect 11411 2150 11463 2202
rect 14973 2150 15025 2202
rect 15037 2150 15089 2202
rect 15101 2150 15153 2202
rect 15165 2150 15217 2202
rect 15229 2150 15281 2202
<< metal2 >>
rect 2226 18856 2282 19656
rect 6550 18856 6606 19656
rect 10874 18986 10930 19656
rect 15198 18986 15254 19656
rect 10874 18958 11008 18986
rect 10874 18856 10930 18958
rect 2240 17270 2268 18856
rect 3519 17436 3827 17445
rect 3519 17434 3525 17436
rect 3581 17434 3605 17436
rect 3661 17434 3685 17436
rect 3741 17434 3765 17436
rect 3821 17434 3827 17436
rect 3581 17382 3583 17434
rect 3763 17382 3765 17434
rect 3519 17380 3525 17382
rect 3581 17380 3605 17382
rect 3661 17380 3685 17382
rect 3741 17380 3765 17382
rect 3821 17380 3827 17382
rect 3519 17371 3827 17380
rect 2228 17264 2280 17270
rect 2228 17206 2280 17212
rect 2504 16992 2556 16998
rect 2504 16934 2556 16940
rect 2516 3602 2544 16934
rect 2859 16892 3167 16901
rect 2859 16890 2865 16892
rect 2921 16890 2945 16892
rect 3001 16890 3025 16892
rect 3081 16890 3105 16892
rect 3161 16890 3167 16892
rect 2921 16838 2923 16890
rect 3103 16838 3105 16890
rect 2859 16836 2865 16838
rect 2921 16836 2945 16838
rect 3001 16836 3025 16838
rect 3081 16836 3105 16838
rect 3161 16836 3167 16838
rect 2859 16827 3167 16836
rect 3519 16348 3827 16357
rect 3519 16346 3525 16348
rect 3581 16346 3605 16348
rect 3661 16346 3685 16348
rect 3741 16346 3765 16348
rect 3821 16346 3827 16348
rect 3581 16294 3583 16346
rect 3763 16294 3765 16346
rect 3519 16292 3525 16294
rect 3581 16292 3605 16294
rect 3661 16292 3685 16294
rect 3741 16292 3765 16294
rect 3821 16292 3827 16294
rect 3519 16283 3827 16292
rect 2859 15804 3167 15813
rect 2859 15802 2865 15804
rect 2921 15802 2945 15804
rect 3001 15802 3025 15804
rect 3081 15802 3105 15804
rect 3161 15802 3167 15804
rect 2921 15750 2923 15802
rect 3103 15750 3105 15802
rect 2859 15748 2865 15750
rect 2921 15748 2945 15750
rect 3001 15748 3025 15750
rect 3081 15748 3105 15750
rect 3161 15748 3167 15750
rect 2859 15739 3167 15748
rect 6564 15366 6592 18856
rect 7337 17436 7645 17445
rect 7337 17434 7343 17436
rect 7399 17434 7423 17436
rect 7479 17434 7503 17436
rect 7559 17434 7583 17436
rect 7639 17434 7645 17436
rect 7399 17382 7401 17434
rect 7581 17382 7583 17434
rect 7337 17380 7343 17382
rect 7399 17380 7423 17382
rect 7479 17380 7503 17382
rect 7559 17380 7583 17382
rect 7639 17380 7645 17382
rect 7337 17371 7645 17380
rect 10980 17354 11008 18958
rect 15198 18958 15424 18986
rect 15198 18856 15254 18958
rect 11155 17436 11463 17445
rect 11155 17434 11161 17436
rect 11217 17434 11241 17436
rect 11297 17434 11321 17436
rect 11377 17434 11401 17436
rect 11457 17434 11463 17436
rect 11217 17382 11219 17434
rect 11399 17382 11401 17434
rect 11155 17380 11161 17382
rect 11217 17380 11241 17382
rect 11297 17380 11321 17382
rect 11377 17380 11401 17382
rect 11457 17380 11463 17382
rect 11155 17371 11463 17380
rect 14973 17436 15281 17445
rect 14973 17434 14979 17436
rect 15035 17434 15059 17436
rect 15115 17434 15139 17436
rect 15195 17434 15219 17436
rect 15275 17434 15281 17436
rect 15035 17382 15037 17434
rect 15217 17382 15219 17434
rect 14973 17380 14979 17382
rect 15035 17380 15059 17382
rect 15115 17380 15139 17382
rect 15195 17380 15219 17382
rect 15275 17380 15281 17382
rect 14973 17371 15281 17380
rect 10980 17338 11100 17354
rect 10980 17332 11112 17338
rect 10980 17326 11060 17332
rect 11060 17274 11112 17280
rect 15396 17270 15424 18958
rect 15384 17264 15436 17270
rect 15384 17206 15436 17212
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 6677 16892 6985 16901
rect 6677 16890 6683 16892
rect 6739 16890 6763 16892
rect 6819 16890 6843 16892
rect 6899 16890 6923 16892
rect 6979 16890 6985 16892
rect 6739 16838 6741 16890
rect 6921 16838 6923 16890
rect 6677 16836 6683 16838
rect 6739 16836 6763 16838
rect 6819 16836 6843 16838
rect 6899 16836 6923 16838
rect 6979 16836 6985 16838
rect 6677 16827 6985 16836
rect 7337 16348 7645 16357
rect 7337 16346 7343 16348
rect 7399 16346 7423 16348
rect 7479 16346 7503 16348
rect 7559 16346 7583 16348
rect 7639 16346 7645 16348
rect 7399 16294 7401 16346
rect 7581 16294 7583 16346
rect 7337 16292 7343 16294
rect 7399 16292 7423 16294
rect 7479 16292 7503 16294
rect 7559 16292 7583 16294
rect 7639 16292 7645 16294
rect 7337 16283 7645 16292
rect 6677 15804 6985 15813
rect 6677 15802 6683 15804
rect 6739 15802 6763 15804
rect 6819 15802 6843 15804
rect 6899 15802 6923 15804
rect 6979 15802 6985 15804
rect 6739 15750 6741 15802
rect 6921 15750 6923 15802
rect 6677 15748 6683 15750
rect 6739 15748 6763 15750
rect 6819 15748 6843 15750
rect 6899 15748 6923 15750
rect 6979 15748 6985 15750
rect 6677 15739 6985 15748
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 3519 15260 3827 15269
rect 3519 15258 3525 15260
rect 3581 15258 3605 15260
rect 3661 15258 3685 15260
rect 3741 15258 3765 15260
rect 3821 15258 3827 15260
rect 3581 15206 3583 15258
rect 3763 15206 3765 15258
rect 3519 15204 3525 15206
rect 3581 15204 3605 15206
rect 3661 15204 3685 15206
rect 3741 15204 3765 15206
rect 3821 15204 3827 15206
rect 3519 15195 3827 15204
rect 2859 14716 3167 14725
rect 2859 14714 2865 14716
rect 2921 14714 2945 14716
rect 3001 14714 3025 14716
rect 3081 14714 3105 14716
rect 3161 14714 3167 14716
rect 2921 14662 2923 14714
rect 3103 14662 3105 14714
rect 2859 14660 2865 14662
rect 2921 14660 2945 14662
rect 3001 14660 3025 14662
rect 3081 14660 3105 14662
rect 3161 14660 3167 14662
rect 2859 14651 3167 14660
rect 6677 14716 6985 14725
rect 6677 14714 6683 14716
rect 6739 14714 6763 14716
rect 6819 14714 6843 14716
rect 6899 14714 6923 14716
rect 6979 14714 6985 14716
rect 6739 14662 6741 14714
rect 6921 14662 6923 14714
rect 6677 14660 6683 14662
rect 6739 14660 6763 14662
rect 6819 14660 6843 14662
rect 6899 14660 6923 14662
rect 6979 14660 6985 14662
rect 6677 14651 6985 14660
rect 3519 14172 3827 14181
rect 3519 14170 3525 14172
rect 3581 14170 3605 14172
rect 3661 14170 3685 14172
rect 3741 14170 3765 14172
rect 3821 14170 3827 14172
rect 3581 14118 3583 14170
rect 3763 14118 3765 14170
rect 3519 14116 3525 14118
rect 3581 14116 3605 14118
rect 3661 14116 3685 14118
rect 3741 14116 3765 14118
rect 3821 14116 3827 14118
rect 3519 14107 3827 14116
rect 2859 13628 3167 13637
rect 2859 13626 2865 13628
rect 2921 13626 2945 13628
rect 3001 13626 3025 13628
rect 3081 13626 3105 13628
rect 3161 13626 3167 13628
rect 2921 13574 2923 13626
rect 3103 13574 3105 13626
rect 2859 13572 2865 13574
rect 2921 13572 2945 13574
rect 3001 13572 3025 13574
rect 3081 13572 3105 13574
rect 3161 13572 3167 13574
rect 2859 13563 3167 13572
rect 6677 13628 6985 13637
rect 6677 13626 6683 13628
rect 6739 13626 6763 13628
rect 6819 13626 6843 13628
rect 6899 13626 6923 13628
rect 6979 13626 6985 13628
rect 6739 13574 6741 13626
rect 6921 13574 6923 13626
rect 6677 13572 6683 13574
rect 6739 13572 6763 13574
rect 6819 13572 6843 13574
rect 6899 13572 6923 13574
rect 6979 13572 6985 13574
rect 6677 13563 6985 13572
rect 3519 13084 3827 13093
rect 3519 13082 3525 13084
rect 3581 13082 3605 13084
rect 3661 13082 3685 13084
rect 3741 13082 3765 13084
rect 3821 13082 3827 13084
rect 3581 13030 3583 13082
rect 3763 13030 3765 13082
rect 3519 13028 3525 13030
rect 3581 13028 3605 13030
rect 3661 13028 3685 13030
rect 3741 13028 3765 13030
rect 3821 13028 3827 13030
rect 3519 13019 3827 13028
rect 2859 12540 3167 12549
rect 2859 12538 2865 12540
rect 2921 12538 2945 12540
rect 3001 12538 3025 12540
rect 3081 12538 3105 12540
rect 3161 12538 3167 12540
rect 2921 12486 2923 12538
rect 3103 12486 3105 12538
rect 2859 12484 2865 12486
rect 2921 12484 2945 12486
rect 3001 12484 3025 12486
rect 3081 12484 3105 12486
rect 3161 12484 3167 12486
rect 2859 12475 3167 12484
rect 6677 12540 6985 12549
rect 6677 12538 6683 12540
rect 6739 12538 6763 12540
rect 6819 12538 6843 12540
rect 6899 12538 6923 12540
rect 6979 12538 6985 12540
rect 6739 12486 6741 12538
rect 6921 12486 6923 12538
rect 6677 12484 6683 12486
rect 6739 12484 6763 12486
rect 6819 12484 6843 12486
rect 6899 12484 6923 12486
rect 6979 12484 6985 12486
rect 6677 12475 6985 12484
rect 3519 11996 3827 12005
rect 3519 11994 3525 11996
rect 3581 11994 3605 11996
rect 3661 11994 3685 11996
rect 3741 11994 3765 11996
rect 3821 11994 3827 11996
rect 3581 11942 3583 11994
rect 3763 11942 3765 11994
rect 3519 11940 3525 11942
rect 3581 11940 3605 11942
rect 3661 11940 3685 11942
rect 3741 11940 3765 11942
rect 3821 11940 3827 11942
rect 3519 11931 3827 11940
rect 2859 11452 3167 11461
rect 2859 11450 2865 11452
rect 2921 11450 2945 11452
rect 3001 11450 3025 11452
rect 3081 11450 3105 11452
rect 3161 11450 3167 11452
rect 2921 11398 2923 11450
rect 3103 11398 3105 11450
rect 2859 11396 2865 11398
rect 2921 11396 2945 11398
rect 3001 11396 3025 11398
rect 3081 11396 3105 11398
rect 3161 11396 3167 11398
rect 2859 11387 3167 11396
rect 6677 11452 6985 11461
rect 6677 11450 6683 11452
rect 6739 11450 6763 11452
rect 6819 11450 6843 11452
rect 6899 11450 6923 11452
rect 6979 11450 6985 11452
rect 6739 11398 6741 11450
rect 6921 11398 6923 11450
rect 6677 11396 6683 11398
rect 6739 11396 6763 11398
rect 6819 11396 6843 11398
rect 6899 11396 6923 11398
rect 6979 11396 6985 11398
rect 6677 11387 6985 11396
rect 3519 10908 3827 10917
rect 3519 10906 3525 10908
rect 3581 10906 3605 10908
rect 3661 10906 3685 10908
rect 3741 10906 3765 10908
rect 3821 10906 3827 10908
rect 3581 10854 3583 10906
rect 3763 10854 3765 10906
rect 3519 10852 3525 10854
rect 3581 10852 3605 10854
rect 3661 10852 3685 10854
rect 3741 10852 3765 10854
rect 3821 10852 3827 10854
rect 3519 10843 3827 10852
rect 2859 10364 3167 10373
rect 2859 10362 2865 10364
rect 2921 10362 2945 10364
rect 3001 10362 3025 10364
rect 3081 10362 3105 10364
rect 3161 10362 3167 10364
rect 2921 10310 2923 10362
rect 3103 10310 3105 10362
rect 2859 10308 2865 10310
rect 2921 10308 2945 10310
rect 3001 10308 3025 10310
rect 3081 10308 3105 10310
rect 3161 10308 3167 10310
rect 2859 10299 3167 10308
rect 6677 10364 6985 10373
rect 6677 10362 6683 10364
rect 6739 10362 6763 10364
rect 6819 10362 6843 10364
rect 6899 10362 6923 10364
rect 6979 10362 6985 10364
rect 6739 10310 6741 10362
rect 6921 10310 6923 10362
rect 6677 10308 6683 10310
rect 6739 10308 6763 10310
rect 6819 10308 6843 10310
rect 6899 10308 6923 10310
rect 6979 10308 6985 10310
rect 6677 10299 6985 10308
rect 3519 9820 3827 9829
rect 3519 9818 3525 9820
rect 3581 9818 3605 9820
rect 3661 9818 3685 9820
rect 3741 9818 3765 9820
rect 3821 9818 3827 9820
rect 3581 9766 3583 9818
rect 3763 9766 3765 9818
rect 3519 9764 3525 9766
rect 3581 9764 3605 9766
rect 3661 9764 3685 9766
rect 3741 9764 3765 9766
rect 3821 9764 3827 9766
rect 3519 9755 3827 9764
rect 2859 9276 3167 9285
rect 2859 9274 2865 9276
rect 2921 9274 2945 9276
rect 3001 9274 3025 9276
rect 3081 9274 3105 9276
rect 3161 9274 3167 9276
rect 2921 9222 2923 9274
rect 3103 9222 3105 9274
rect 2859 9220 2865 9222
rect 2921 9220 2945 9222
rect 3001 9220 3025 9222
rect 3081 9220 3105 9222
rect 3161 9220 3167 9222
rect 2859 9211 3167 9220
rect 6677 9276 6985 9285
rect 6677 9274 6683 9276
rect 6739 9274 6763 9276
rect 6819 9274 6843 9276
rect 6899 9274 6923 9276
rect 6979 9274 6985 9276
rect 6739 9222 6741 9274
rect 6921 9222 6923 9274
rect 6677 9220 6683 9222
rect 6739 9220 6763 9222
rect 6819 9220 6843 9222
rect 6899 9220 6923 9222
rect 6979 9220 6985 9222
rect 6677 9211 6985 9220
rect 3519 8732 3827 8741
rect 3519 8730 3525 8732
rect 3581 8730 3605 8732
rect 3661 8730 3685 8732
rect 3741 8730 3765 8732
rect 3821 8730 3827 8732
rect 3581 8678 3583 8730
rect 3763 8678 3765 8730
rect 3519 8676 3525 8678
rect 3581 8676 3605 8678
rect 3661 8676 3685 8678
rect 3741 8676 3765 8678
rect 3821 8676 3827 8678
rect 3519 8667 3827 8676
rect 2859 8188 3167 8197
rect 2859 8186 2865 8188
rect 2921 8186 2945 8188
rect 3001 8186 3025 8188
rect 3081 8186 3105 8188
rect 3161 8186 3167 8188
rect 2921 8134 2923 8186
rect 3103 8134 3105 8186
rect 2859 8132 2865 8134
rect 2921 8132 2945 8134
rect 3001 8132 3025 8134
rect 3081 8132 3105 8134
rect 3161 8132 3167 8134
rect 2859 8123 3167 8132
rect 6677 8188 6985 8197
rect 6677 8186 6683 8188
rect 6739 8186 6763 8188
rect 6819 8186 6843 8188
rect 6899 8186 6923 8188
rect 6979 8186 6985 8188
rect 6739 8134 6741 8186
rect 6921 8134 6923 8186
rect 6677 8132 6683 8134
rect 6739 8132 6763 8134
rect 6819 8132 6843 8134
rect 6899 8132 6923 8134
rect 6979 8132 6985 8134
rect 6677 8123 6985 8132
rect 3519 7644 3827 7653
rect 3519 7642 3525 7644
rect 3581 7642 3605 7644
rect 3661 7642 3685 7644
rect 3741 7642 3765 7644
rect 3821 7642 3827 7644
rect 3581 7590 3583 7642
rect 3763 7590 3765 7642
rect 3519 7588 3525 7590
rect 3581 7588 3605 7590
rect 3661 7588 3685 7590
rect 3741 7588 3765 7590
rect 3821 7588 3827 7590
rect 3519 7579 3827 7588
rect 2859 7100 3167 7109
rect 2859 7098 2865 7100
rect 2921 7098 2945 7100
rect 3001 7098 3025 7100
rect 3081 7098 3105 7100
rect 3161 7098 3167 7100
rect 2921 7046 2923 7098
rect 3103 7046 3105 7098
rect 2859 7044 2865 7046
rect 2921 7044 2945 7046
rect 3001 7044 3025 7046
rect 3081 7044 3105 7046
rect 3161 7044 3167 7046
rect 2859 7035 3167 7044
rect 6677 7100 6985 7109
rect 6677 7098 6683 7100
rect 6739 7098 6763 7100
rect 6819 7098 6843 7100
rect 6899 7098 6923 7100
rect 6979 7098 6985 7100
rect 6739 7046 6741 7098
rect 6921 7046 6923 7098
rect 6677 7044 6683 7046
rect 6739 7044 6763 7046
rect 6819 7044 6843 7046
rect 6899 7044 6923 7046
rect 6979 7044 6985 7046
rect 6677 7035 6985 7044
rect 3519 6556 3827 6565
rect 3519 6554 3525 6556
rect 3581 6554 3605 6556
rect 3661 6554 3685 6556
rect 3741 6554 3765 6556
rect 3821 6554 3827 6556
rect 3581 6502 3583 6554
rect 3763 6502 3765 6554
rect 3519 6500 3525 6502
rect 3581 6500 3605 6502
rect 3661 6500 3685 6502
rect 3741 6500 3765 6502
rect 3821 6500 3827 6502
rect 3519 6491 3827 6500
rect 2859 6012 3167 6021
rect 2859 6010 2865 6012
rect 2921 6010 2945 6012
rect 3001 6010 3025 6012
rect 3081 6010 3105 6012
rect 3161 6010 3167 6012
rect 2921 5958 2923 6010
rect 3103 5958 3105 6010
rect 2859 5956 2865 5958
rect 2921 5956 2945 5958
rect 3001 5956 3025 5958
rect 3081 5956 3105 5958
rect 3161 5956 3167 5958
rect 2859 5947 3167 5956
rect 6677 6012 6985 6021
rect 6677 6010 6683 6012
rect 6739 6010 6763 6012
rect 6819 6010 6843 6012
rect 6899 6010 6923 6012
rect 6979 6010 6985 6012
rect 6739 5958 6741 6010
rect 6921 5958 6923 6010
rect 6677 5956 6683 5958
rect 6739 5956 6763 5958
rect 6819 5956 6843 5958
rect 6899 5956 6923 5958
rect 6979 5956 6985 5958
rect 6677 5947 6985 5956
rect 3519 5468 3827 5477
rect 3519 5466 3525 5468
rect 3581 5466 3605 5468
rect 3661 5466 3685 5468
rect 3741 5466 3765 5468
rect 3821 5466 3827 5468
rect 3581 5414 3583 5466
rect 3763 5414 3765 5466
rect 3519 5412 3525 5414
rect 3581 5412 3605 5414
rect 3661 5412 3685 5414
rect 3741 5412 3765 5414
rect 3821 5412 3827 5414
rect 3519 5403 3827 5412
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 2859 4924 3167 4933
rect 2859 4922 2865 4924
rect 2921 4922 2945 4924
rect 3001 4922 3025 4924
rect 3081 4922 3105 4924
rect 3161 4922 3167 4924
rect 2921 4870 2923 4922
rect 3103 4870 3105 4922
rect 2859 4868 2865 4870
rect 2921 4868 2945 4870
rect 3001 4868 3025 4870
rect 3081 4868 3105 4870
rect 3161 4868 3167 4870
rect 2859 4859 3167 4868
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 3519 4380 3827 4389
rect 3519 4378 3525 4380
rect 3581 4378 3605 4380
rect 3661 4378 3685 4380
rect 3741 4378 3765 4380
rect 3821 4378 3827 4380
rect 3581 4326 3583 4378
rect 3763 4326 3765 4378
rect 3519 4324 3525 4326
rect 3581 4324 3605 4326
rect 3661 4324 3685 4326
rect 3741 4324 3765 4326
rect 3821 4324 3827 4326
rect 3519 4315 3827 4324
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 2859 3836 3167 3845
rect 2859 3834 2865 3836
rect 2921 3834 2945 3836
rect 3001 3834 3025 3836
rect 3081 3834 3105 3836
rect 3161 3834 3167 3836
rect 2921 3782 2923 3834
rect 3103 3782 3105 3834
rect 2859 3780 2865 3782
rect 2921 3780 2945 3782
rect 3001 3780 3025 3782
rect 3081 3780 3105 3782
rect 3161 3780 3167 3782
rect 2859 3771 3167 3780
rect 4172 3602 4200 3878
rect 4816 3738 4844 4082
rect 5000 3738 5028 4558
rect 5184 4282 5212 4966
rect 5264 4548 5316 4554
rect 5264 4490 5316 4496
rect 5724 4548 5776 4554
rect 5724 4490 5776 4496
rect 5276 4282 5304 4490
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5644 4282 5672 4422
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 5264 4276 5316 4282
rect 5264 4218 5316 4224
rect 5632 4276 5684 4282
rect 5632 4218 5684 4224
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 2504 3596 2556 3602
rect 2504 3538 2556 3544
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 4344 3528 4396 3534
rect 4344 3470 4396 3476
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 3519 3292 3827 3301
rect 3519 3290 3525 3292
rect 3581 3290 3605 3292
rect 3661 3290 3685 3292
rect 3741 3290 3765 3292
rect 3821 3290 3827 3292
rect 3581 3238 3583 3290
rect 3763 3238 3765 3290
rect 3519 3236 3525 3238
rect 3581 3236 3605 3238
rect 3661 3236 3685 3238
rect 3741 3236 3765 3238
rect 3821 3236 3827 3238
rect 3519 3227 3827 3236
rect 4264 3194 4292 3334
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 3700 2984 3752 2990
rect 3700 2926 3752 2932
rect 2859 2748 3167 2757
rect 2859 2746 2865 2748
rect 2921 2746 2945 2748
rect 3001 2746 3025 2748
rect 3081 2746 3105 2748
rect 3161 2746 3167 2748
rect 2921 2694 2923 2746
rect 3103 2694 3105 2746
rect 2859 2692 2865 2694
rect 2921 2692 2945 2694
rect 3001 2692 3025 2694
rect 3081 2692 3105 2694
rect 3161 2692 3167 2694
rect 2859 2683 3167 2692
rect 3712 2446 3740 2926
rect 4356 2446 4384 3470
rect 5000 3194 5028 3674
rect 4988 3188 5040 3194
rect 4988 3130 5040 3136
rect 5552 2514 5580 3878
rect 5644 3534 5672 4218
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5736 3058 5764 4490
rect 5920 4282 5948 5102
rect 6677 4924 6985 4933
rect 6677 4922 6683 4924
rect 6739 4922 6763 4924
rect 6819 4922 6843 4924
rect 6899 4922 6923 4924
rect 6979 4922 6985 4924
rect 6739 4870 6741 4922
rect 6921 4870 6923 4922
rect 6677 4868 6683 4870
rect 6739 4868 6763 4870
rect 6819 4868 6843 4870
rect 6899 4868 6923 4870
rect 6979 4868 6985 4870
rect 6677 4859 6985 4868
rect 6276 4752 6328 4758
rect 6276 4694 6328 4700
rect 5908 4276 5960 4282
rect 5908 4218 5960 4224
rect 6184 3596 6236 3602
rect 6184 3538 6236 3544
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 3700 2440 3752 2446
rect 3700 2382 3752 2388
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 1308 2372 1360 2378
rect 1308 2314 1360 2320
rect 3424 2372 3476 2378
rect 3424 2314 3476 2320
rect 5632 2372 5684 2378
rect 5632 2314 5684 2320
rect 1320 800 1348 2314
rect 3436 800 3464 2314
rect 3519 2204 3827 2213
rect 3519 2202 3525 2204
rect 3581 2202 3605 2204
rect 3661 2202 3685 2204
rect 3741 2202 3765 2204
rect 3821 2202 3827 2204
rect 3581 2150 3583 2202
rect 3763 2150 3765 2202
rect 3519 2148 3525 2150
rect 3581 2148 3605 2150
rect 3661 2148 3685 2150
rect 3741 2148 3765 2150
rect 3821 2148 3827 2150
rect 3519 2139 3827 2148
rect 5644 1170 5672 2314
rect 5736 2310 5764 2994
rect 6196 2514 6224 3538
rect 6288 3126 6316 4694
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 6932 4078 6960 4422
rect 6460 4072 6512 4078
rect 6460 4014 6512 4020
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 6472 3126 6500 4014
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6564 3534 6592 3878
rect 6677 3836 6985 3845
rect 6677 3834 6683 3836
rect 6739 3834 6763 3836
rect 6819 3834 6843 3836
rect 6899 3834 6923 3836
rect 6979 3834 6985 3836
rect 6739 3782 6741 3834
rect 6921 3782 6923 3834
rect 6677 3780 6683 3782
rect 6739 3780 6763 3782
rect 6819 3780 6843 3782
rect 6899 3780 6923 3782
rect 6979 3780 6985 3782
rect 6677 3771 6985 3780
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6840 3194 6868 3334
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6276 3120 6328 3126
rect 6276 3062 6328 3068
rect 6460 3120 6512 3126
rect 6460 3062 6512 3068
rect 6552 3120 6604 3126
rect 6552 3062 6604 3068
rect 6564 2650 6592 3062
rect 7024 2922 7052 4558
rect 7208 4162 7236 15302
rect 7337 15260 7645 15269
rect 7337 15258 7343 15260
rect 7399 15258 7423 15260
rect 7479 15258 7503 15260
rect 7559 15258 7583 15260
rect 7639 15258 7645 15260
rect 7399 15206 7401 15258
rect 7581 15206 7583 15258
rect 7337 15204 7343 15206
rect 7399 15204 7423 15206
rect 7479 15204 7503 15206
rect 7559 15204 7583 15206
rect 7639 15204 7645 15206
rect 7337 15195 7645 15204
rect 7337 14172 7645 14181
rect 7337 14170 7343 14172
rect 7399 14170 7423 14172
rect 7479 14170 7503 14172
rect 7559 14170 7583 14172
rect 7639 14170 7645 14172
rect 7399 14118 7401 14170
rect 7581 14118 7583 14170
rect 7337 14116 7343 14118
rect 7399 14116 7423 14118
rect 7479 14116 7503 14118
rect 7559 14116 7583 14118
rect 7639 14116 7645 14118
rect 7337 14107 7645 14116
rect 7337 13084 7645 13093
rect 7337 13082 7343 13084
rect 7399 13082 7423 13084
rect 7479 13082 7503 13084
rect 7559 13082 7583 13084
rect 7639 13082 7645 13084
rect 7399 13030 7401 13082
rect 7581 13030 7583 13082
rect 7337 13028 7343 13030
rect 7399 13028 7423 13030
rect 7479 13028 7503 13030
rect 7559 13028 7583 13030
rect 7639 13028 7645 13030
rect 7337 13019 7645 13028
rect 7337 11996 7645 12005
rect 7337 11994 7343 11996
rect 7399 11994 7423 11996
rect 7479 11994 7503 11996
rect 7559 11994 7583 11996
rect 7639 11994 7645 11996
rect 7399 11942 7401 11994
rect 7581 11942 7583 11994
rect 7337 11940 7343 11942
rect 7399 11940 7423 11942
rect 7479 11940 7503 11942
rect 7559 11940 7583 11942
rect 7639 11940 7645 11942
rect 7337 11931 7645 11940
rect 7337 10908 7645 10917
rect 7337 10906 7343 10908
rect 7399 10906 7423 10908
rect 7479 10906 7503 10908
rect 7559 10906 7583 10908
rect 7639 10906 7645 10908
rect 7399 10854 7401 10906
rect 7581 10854 7583 10906
rect 7337 10852 7343 10854
rect 7399 10852 7423 10854
rect 7479 10852 7503 10854
rect 7559 10852 7583 10854
rect 7639 10852 7645 10854
rect 7337 10843 7645 10852
rect 7337 9820 7645 9829
rect 7337 9818 7343 9820
rect 7399 9818 7423 9820
rect 7479 9818 7503 9820
rect 7559 9818 7583 9820
rect 7639 9818 7645 9820
rect 7399 9766 7401 9818
rect 7581 9766 7583 9818
rect 7337 9764 7343 9766
rect 7399 9764 7423 9766
rect 7479 9764 7503 9766
rect 7559 9764 7583 9766
rect 7639 9764 7645 9766
rect 7337 9755 7645 9764
rect 7337 8732 7645 8741
rect 7337 8730 7343 8732
rect 7399 8730 7423 8732
rect 7479 8730 7503 8732
rect 7559 8730 7583 8732
rect 7639 8730 7645 8732
rect 7399 8678 7401 8730
rect 7581 8678 7583 8730
rect 7337 8676 7343 8678
rect 7399 8676 7423 8678
rect 7479 8676 7503 8678
rect 7559 8676 7583 8678
rect 7639 8676 7645 8678
rect 7337 8667 7645 8676
rect 7337 7644 7645 7653
rect 7337 7642 7343 7644
rect 7399 7642 7423 7644
rect 7479 7642 7503 7644
rect 7559 7642 7583 7644
rect 7639 7642 7645 7644
rect 7399 7590 7401 7642
rect 7581 7590 7583 7642
rect 7337 7588 7343 7590
rect 7399 7588 7423 7590
rect 7479 7588 7503 7590
rect 7559 7588 7583 7590
rect 7639 7588 7645 7590
rect 7337 7579 7645 7588
rect 7337 6556 7645 6565
rect 7337 6554 7343 6556
rect 7399 6554 7423 6556
rect 7479 6554 7503 6556
rect 7559 6554 7583 6556
rect 7639 6554 7645 6556
rect 7399 6502 7401 6554
rect 7581 6502 7583 6554
rect 7337 6500 7343 6502
rect 7399 6500 7423 6502
rect 7479 6500 7503 6502
rect 7559 6500 7583 6502
rect 7639 6500 7645 6502
rect 7337 6491 7645 6500
rect 7337 5468 7645 5477
rect 7337 5466 7343 5468
rect 7399 5466 7423 5468
rect 7479 5466 7503 5468
rect 7559 5466 7583 5468
rect 7639 5466 7645 5468
rect 7399 5414 7401 5466
rect 7581 5414 7583 5466
rect 7337 5412 7343 5414
rect 7399 5412 7423 5414
rect 7479 5412 7503 5414
rect 7559 5412 7583 5414
rect 7639 5412 7645 5414
rect 7337 5403 7645 5412
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 7852 4826 7880 4966
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 7337 4380 7645 4389
rect 7337 4378 7343 4380
rect 7399 4378 7423 4380
rect 7479 4378 7503 4380
rect 7559 4378 7583 4380
rect 7639 4378 7645 4380
rect 7399 4326 7401 4378
rect 7581 4326 7583 4378
rect 7337 4324 7343 4326
rect 7399 4324 7423 4326
rect 7479 4324 7503 4326
rect 7559 4324 7583 4326
rect 7639 4324 7645 4326
rect 7337 4315 7645 4324
rect 7288 4208 7340 4214
rect 7208 4156 7288 4162
rect 7208 4150 7340 4156
rect 7208 4134 7328 4150
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 7012 2916 7064 2922
rect 7012 2858 7064 2864
rect 7116 2854 7144 4014
rect 7196 3460 7248 3466
rect 7196 3402 7248 3408
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 6677 2748 6985 2757
rect 6677 2746 6683 2748
rect 6739 2746 6763 2748
rect 6819 2746 6843 2748
rect 6899 2746 6923 2748
rect 6979 2746 6985 2748
rect 6739 2694 6741 2746
rect 6921 2694 6923 2746
rect 6677 2692 6683 2694
rect 6739 2692 6763 2694
rect 6819 2692 6843 2694
rect 6899 2692 6923 2694
rect 6979 2692 6985 2694
rect 6677 2683 6985 2692
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 7116 2514 7144 2790
rect 7208 2650 7236 3402
rect 7337 3292 7645 3301
rect 7337 3290 7343 3292
rect 7399 3290 7423 3292
rect 7479 3290 7503 3292
rect 7559 3290 7583 3292
rect 7639 3290 7645 3292
rect 7399 3238 7401 3290
rect 7581 3238 7583 3290
rect 7337 3236 7343 3238
rect 7399 3236 7423 3238
rect 7479 3236 7503 3238
rect 7559 3236 7583 3238
rect 7639 3236 7645 3238
rect 7337 3227 7645 3236
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 7852 2446 7880 4422
rect 8220 3738 8248 4422
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8220 2990 8248 3674
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 8220 2530 8248 2926
rect 8404 2854 8432 5102
rect 9588 4684 9640 4690
rect 9588 4626 9640 4632
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8588 3738 8616 3878
rect 9416 3738 9444 4014
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 8128 2502 8248 2530
rect 8128 2446 8156 2502
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 8404 2310 8432 2790
rect 8588 2650 8616 3470
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8772 2990 8800 3334
rect 9416 3194 9444 3674
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 9600 2514 9628 4626
rect 10244 4622 10272 16934
rect 10495 16892 10803 16901
rect 10495 16890 10501 16892
rect 10557 16890 10581 16892
rect 10637 16890 10661 16892
rect 10717 16890 10741 16892
rect 10797 16890 10803 16892
rect 10557 16838 10559 16890
rect 10739 16838 10741 16890
rect 10495 16836 10501 16838
rect 10557 16836 10581 16838
rect 10637 16836 10661 16838
rect 10717 16836 10741 16838
rect 10797 16836 10803 16838
rect 10495 16827 10803 16836
rect 14313 16892 14621 16901
rect 14313 16890 14319 16892
rect 14375 16890 14399 16892
rect 14455 16890 14479 16892
rect 14535 16890 14559 16892
rect 14615 16890 14621 16892
rect 14375 16838 14377 16890
rect 14557 16838 14559 16890
rect 14313 16836 14319 16838
rect 14375 16836 14399 16838
rect 14455 16836 14479 16838
rect 14535 16836 14559 16838
rect 14615 16836 14621 16838
rect 14313 16827 14621 16836
rect 11155 16348 11463 16357
rect 11155 16346 11161 16348
rect 11217 16346 11241 16348
rect 11297 16346 11321 16348
rect 11377 16346 11401 16348
rect 11457 16346 11463 16348
rect 11217 16294 11219 16346
rect 11399 16294 11401 16346
rect 11155 16292 11161 16294
rect 11217 16292 11241 16294
rect 11297 16292 11321 16294
rect 11377 16292 11401 16294
rect 11457 16292 11463 16294
rect 11155 16283 11463 16292
rect 14973 16348 15281 16357
rect 14973 16346 14979 16348
rect 15035 16346 15059 16348
rect 15115 16346 15139 16348
rect 15195 16346 15219 16348
rect 15275 16346 15281 16348
rect 15035 16294 15037 16346
rect 15217 16294 15219 16346
rect 14973 16292 14979 16294
rect 15035 16292 15059 16294
rect 15115 16292 15139 16294
rect 15195 16292 15219 16294
rect 15275 16292 15281 16294
rect 14973 16283 15281 16292
rect 10495 15804 10803 15813
rect 10495 15802 10501 15804
rect 10557 15802 10581 15804
rect 10637 15802 10661 15804
rect 10717 15802 10741 15804
rect 10797 15802 10803 15804
rect 10557 15750 10559 15802
rect 10739 15750 10741 15802
rect 10495 15748 10501 15750
rect 10557 15748 10581 15750
rect 10637 15748 10661 15750
rect 10717 15748 10741 15750
rect 10797 15748 10803 15750
rect 10495 15739 10803 15748
rect 14313 15804 14621 15813
rect 14313 15802 14319 15804
rect 14375 15802 14399 15804
rect 14455 15802 14479 15804
rect 14535 15802 14559 15804
rect 14615 15802 14621 15804
rect 14375 15750 14377 15802
rect 14557 15750 14559 15802
rect 14313 15748 14319 15750
rect 14375 15748 14399 15750
rect 14455 15748 14479 15750
rect 14535 15748 14559 15750
rect 14615 15748 14621 15750
rect 14313 15739 14621 15748
rect 11155 15260 11463 15269
rect 11155 15258 11161 15260
rect 11217 15258 11241 15260
rect 11297 15258 11321 15260
rect 11377 15258 11401 15260
rect 11457 15258 11463 15260
rect 11217 15206 11219 15258
rect 11399 15206 11401 15258
rect 11155 15204 11161 15206
rect 11217 15204 11241 15206
rect 11297 15204 11321 15206
rect 11377 15204 11401 15206
rect 11457 15204 11463 15206
rect 11155 15195 11463 15204
rect 14973 15260 15281 15269
rect 14973 15258 14979 15260
rect 15035 15258 15059 15260
rect 15115 15258 15139 15260
rect 15195 15258 15219 15260
rect 15275 15258 15281 15260
rect 15035 15206 15037 15258
rect 15217 15206 15219 15258
rect 14973 15204 14979 15206
rect 15035 15204 15059 15206
rect 15115 15204 15139 15206
rect 15195 15204 15219 15206
rect 15275 15204 15281 15206
rect 14973 15195 15281 15204
rect 10495 14716 10803 14725
rect 10495 14714 10501 14716
rect 10557 14714 10581 14716
rect 10637 14714 10661 14716
rect 10717 14714 10741 14716
rect 10797 14714 10803 14716
rect 10557 14662 10559 14714
rect 10739 14662 10741 14714
rect 10495 14660 10501 14662
rect 10557 14660 10581 14662
rect 10637 14660 10661 14662
rect 10717 14660 10741 14662
rect 10797 14660 10803 14662
rect 10495 14651 10803 14660
rect 14313 14716 14621 14725
rect 14313 14714 14319 14716
rect 14375 14714 14399 14716
rect 14455 14714 14479 14716
rect 14535 14714 14559 14716
rect 14615 14714 14621 14716
rect 14375 14662 14377 14714
rect 14557 14662 14559 14714
rect 14313 14660 14319 14662
rect 14375 14660 14399 14662
rect 14455 14660 14479 14662
rect 14535 14660 14559 14662
rect 14615 14660 14621 14662
rect 14313 14651 14621 14660
rect 11155 14172 11463 14181
rect 11155 14170 11161 14172
rect 11217 14170 11241 14172
rect 11297 14170 11321 14172
rect 11377 14170 11401 14172
rect 11457 14170 11463 14172
rect 11217 14118 11219 14170
rect 11399 14118 11401 14170
rect 11155 14116 11161 14118
rect 11217 14116 11241 14118
rect 11297 14116 11321 14118
rect 11377 14116 11401 14118
rect 11457 14116 11463 14118
rect 11155 14107 11463 14116
rect 14973 14172 15281 14181
rect 14973 14170 14979 14172
rect 15035 14170 15059 14172
rect 15115 14170 15139 14172
rect 15195 14170 15219 14172
rect 15275 14170 15281 14172
rect 15035 14118 15037 14170
rect 15217 14118 15219 14170
rect 14973 14116 14979 14118
rect 15035 14116 15059 14118
rect 15115 14116 15139 14118
rect 15195 14116 15219 14118
rect 15275 14116 15281 14118
rect 14973 14107 15281 14116
rect 10495 13628 10803 13637
rect 10495 13626 10501 13628
rect 10557 13626 10581 13628
rect 10637 13626 10661 13628
rect 10717 13626 10741 13628
rect 10797 13626 10803 13628
rect 10557 13574 10559 13626
rect 10739 13574 10741 13626
rect 10495 13572 10501 13574
rect 10557 13572 10581 13574
rect 10637 13572 10661 13574
rect 10717 13572 10741 13574
rect 10797 13572 10803 13574
rect 10495 13563 10803 13572
rect 14313 13628 14621 13637
rect 14313 13626 14319 13628
rect 14375 13626 14399 13628
rect 14455 13626 14479 13628
rect 14535 13626 14559 13628
rect 14615 13626 14621 13628
rect 14375 13574 14377 13626
rect 14557 13574 14559 13626
rect 14313 13572 14319 13574
rect 14375 13572 14399 13574
rect 14455 13572 14479 13574
rect 14535 13572 14559 13574
rect 14615 13572 14621 13574
rect 14313 13563 14621 13572
rect 11155 13084 11463 13093
rect 11155 13082 11161 13084
rect 11217 13082 11241 13084
rect 11297 13082 11321 13084
rect 11377 13082 11401 13084
rect 11457 13082 11463 13084
rect 11217 13030 11219 13082
rect 11399 13030 11401 13082
rect 11155 13028 11161 13030
rect 11217 13028 11241 13030
rect 11297 13028 11321 13030
rect 11377 13028 11401 13030
rect 11457 13028 11463 13030
rect 11155 13019 11463 13028
rect 14973 13084 15281 13093
rect 14973 13082 14979 13084
rect 15035 13082 15059 13084
rect 15115 13082 15139 13084
rect 15195 13082 15219 13084
rect 15275 13082 15281 13084
rect 15035 13030 15037 13082
rect 15217 13030 15219 13082
rect 14973 13028 14979 13030
rect 15035 13028 15059 13030
rect 15115 13028 15139 13030
rect 15195 13028 15219 13030
rect 15275 13028 15281 13030
rect 14973 13019 15281 13028
rect 10495 12540 10803 12549
rect 10495 12538 10501 12540
rect 10557 12538 10581 12540
rect 10637 12538 10661 12540
rect 10717 12538 10741 12540
rect 10797 12538 10803 12540
rect 10557 12486 10559 12538
rect 10739 12486 10741 12538
rect 10495 12484 10501 12486
rect 10557 12484 10581 12486
rect 10637 12484 10661 12486
rect 10717 12484 10741 12486
rect 10797 12484 10803 12486
rect 10495 12475 10803 12484
rect 14313 12540 14621 12549
rect 14313 12538 14319 12540
rect 14375 12538 14399 12540
rect 14455 12538 14479 12540
rect 14535 12538 14559 12540
rect 14615 12538 14621 12540
rect 14375 12486 14377 12538
rect 14557 12486 14559 12538
rect 14313 12484 14319 12486
rect 14375 12484 14399 12486
rect 14455 12484 14479 12486
rect 14535 12484 14559 12486
rect 14615 12484 14621 12486
rect 14313 12475 14621 12484
rect 11155 11996 11463 12005
rect 11155 11994 11161 11996
rect 11217 11994 11241 11996
rect 11297 11994 11321 11996
rect 11377 11994 11401 11996
rect 11457 11994 11463 11996
rect 11217 11942 11219 11994
rect 11399 11942 11401 11994
rect 11155 11940 11161 11942
rect 11217 11940 11241 11942
rect 11297 11940 11321 11942
rect 11377 11940 11401 11942
rect 11457 11940 11463 11942
rect 11155 11931 11463 11940
rect 14973 11996 15281 12005
rect 14973 11994 14979 11996
rect 15035 11994 15059 11996
rect 15115 11994 15139 11996
rect 15195 11994 15219 11996
rect 15275 11994 15281 11996
rect 15035 11942 15037 11994
rect 15217 11942 15219 11994
rect 14973 11940 14979 11942
rect 15035 11940 15059 11942
rect 15115 11940 15139 11942
rect 15195 11940 15219 11942
rect 15275 11940 15281 11942
rect 14973 11931 15281 11940
rect 10495 11452 10803 11461
rect 10495 11450 10501 11452
rect 10557 11450 10581 11452
rect 10637 11450 10661 11452
rect 10717 11450 10741 11452
rect 10797 11450 10803 11452
rect 10557 11398 10559 11450
rect 10739 11398 10741 11450
rect 10495 11396 10501 11398
rect 10557 11396 10581 11398
rect 10637 11396 10661 11398
rect 10717 11396 10741 11398
rect 10797 11396 10803 11398
rect 10495 11387 10803 11396
rect 14313 11452 14621 11461
rect 14313 11450 14319 11452
rect 14375 11450 14399 11452
rect 14455 11450 14479 11452
rect 14535 11450 14559 11452
rect 14615 11450 14621 11452
rect 14375 11398 14377 11450
rect 14557 11398 14559 11450
rect 14313 11396 14319 11398
rect 14375 11396 14399 11398
rect 14455 11396 14479 11398
rect 14535 11396 14559 11398
rect 14615 11396 14621 11398
rect 14313 11387 14621 11396
rect 11155 10908 11463 10917
rect 11155 10906 11161 10908
rect 11217 10906 11241 10908
rect 11297 10906 11321 10908
rect 11377 10906 11401 10908
rect 11457 10906 11463 10908
rect 11217 10854 11219 10906
rect 11399 10854 11401 10906
rect 11155 10852 11161 10854
rect 11217 10852 11241 10854
rect 11297 10852 11321 10854
rect 11377 10852 11401 10854
rect 11457 10852 11463 10854
rect 11155 10843 11463 10852
rect 14973 10908 15281 10917
rect 14973 10906 14979 10908
rect 15035 10906 15059 10908
rect 15115 10906 15139 10908
rect 15195 10906 15219 10908
rect 15275 10906 15281 10908
rect 15035 10854 15037 10906
rect 15217 10854 15219 10906
rect 14973 10852 14979 10854
rect 15035 10852 15059 10854
rect 15115 10852 15139 10854
rect 15195 10852 15219 10854
rect 15275 10852 15281 10854
rect 14973 10843 15281 10852
rect 10495 10364 10803 10373
rect 10495 10362 10501 10364
rect 10557 10362 10581 10364
rect 10637 10362 10661 10364
rect 10717 10362 10741 10364
rect 10797 10362 10803 10364
rect 10557 10310 10559 10362
rect 10739 10310 10741 10362
rect 10495 10308 10501 10310
rect 10557 10308 10581 10310
rect 10637 10308 10661 10310
rect 10717 10308 10741 10310
rect 10797 10308 10803 10310
rect 10495 10299 10803 10308
rect 14313 10364 14621 10373
rect 14313 10362 14319 10364
rect 14375 10362 14399 10364
rect 14455 10362 14479 10364
rect 14535 10362 14559 10364
rect 14615 10362 14621 10364
rect 14375 10310 14377 10362
rect 14557 10310 14559 10362
rect 14313 10308 14319 10310
rect 14375 10308 14399 10310
rect 14455 10308 14479 10310
rect 14535 10308 14559 10310
rect 14615 10308 14621 10310
rect 14313 10299 14621 10308
rect 11155 9820 11463 9829
rect 11155 9818 11161 9820
rect 11217 9818 11241 9820
rect 11297 9818 11321 9820
rect 11377 9818 11401 9820
rect 11457 9818 11463 9820
rect 11217 9766 11219 9818
rect 11399 9766 11401 9818
rect 11155 9764 11161 9766
rect 11217 9764 11241 9766
rect 11297 9764 11321 9766
rect 11377 9764 11401 9766
rect 11457 9764 11463 9766
rect 11155 9755 11463 9764
rect 14973 9820 15281 9829
rect 14973 9818 14979 9820
rect 15035 9818 15059 9820
rect 15115 9818 15139 9820
rect 15195 9818 15219 9820
rect 15275 9818 15281 9820
rect 15035 9766 15037 9818
rect 15217 9766 15219 9818
rect 14973 9764 14979 9766
rect 15035 9764 15059 9766
rect 15115 9764 15139 9766
rect 15195 9764 15219 9766
rect 15275 9764 15281 9766
rect 14973 9755 15281 9764
rect 10495 9276 10803 9285
rect 10495 9274 10501 9276
rect 10557 9274 10581 9276
rect 10637 9274 10661 9276
rect 10717 9274 10741 9276
rect 10797 9274 10803 9276
rect 10557 9222 10559 9274
rect 10739 9222 10741 9274
rect 10495 9220 10501 9222
rect 10557 9220 10581 9222
rect 10637 9220 10661 9222
rect 10717 9220 10741 9222
rect 10797 9220 10803 9222
rect 10495 9211 10803 9220
rect 14313 9276 14621 9285
rect 14313 9274 14319 9276
rect 14375 9274 14399 9276
rect 14455 9274 14479 9276
rect 14535 9274 14559 9276
rect 14615 9274 14621 9276
rect 14375 9222 14377 9274
rect 14557 9222 14559 9274
rect 14313 9220 14319 9222
rect 14375 9220 14399 9222
rect 14455 9220 14479 9222
rect 14535 9220 14559 9222
rect 14615 9220 14621 9222
rect 14313 9211 14621 9220
rect 11155 8732 11463 8741
rect 11155 8730 11161 8732
rect 11217 8730 11241 8732
rect 11297 8730 11321 8732
rect 11377 8730 11401 8732
rect 11457 8730 11463 8732
rect 11217 8678 11219 8730
rect 11399 8678 11401 8730
rect 11155 8676 11161 8678
rect 11217 8676 11241 8678
rect 11297 8676 11321 8678
rect 11377 8676 11401 8678
rect 11457 8676 11463 8678
rect 11155 8667 11463 8676
rect 14973 8732 15281 8741
rect 14973 8730 14979 8732
rect 15035 8730 15059 8732
rect 15115 8730 15139 8732
rect 15195 8730 15219 8732
rect 15275 8730 15281 8732
rect 15035 8678 15037 8730
rect 15217 8678 15219 8730
rect 14973 8676 14979 8678
rect 15035 8676 15059 8678
rect 15115 8676 15139 8678
rect 15195 8676 15219 8678
rect 15275 8676 15281 8678
rect 14973 8667 15281 8676
rect 10495 8188 10803 8197
rect 10495 8186 10501 8188
rect 10557 8186 10581 8188
rect 10637 8186 10661 8188
rect 10717 8186 10741 8188
rect 10797 8186 10803 8188
rect 10557 8134 10559 8186
rect 10739 8134 10741 8186
rect 10495 8132 10501 8134
rect 10557 8132 10581 8134
rect 10637 8132 10661 8134
rect 10717 8132 10741 8134
rect 10797 8132 10803 8134
rect 10495 8123 10803 8132
rect 14313 8188 14621 8197
rect 14313 8186 14319 8188
rect 14375 8186 14399 8188
rect 14455 8186 14479 8188
rect 14535 8186 14559 8188
rect 14615 8186 14621 8188
rect 14375 8134 14377 8186
rect 14557 8134 14559 8186
rect 14313 8132 14319 8134
rect 14375 8132 14399 8134
rect 14455 8132 14479 8134
rect 14535 8132 14559 8134
rect 14615 8132 14621 8134
rect 14313 8123 14621 8132
rect 11155 7644 11463 7653
rect 11155 7642 11161 7644
rect 11217 7642 11241 7644
rect 11297 7642 11321 7644
rect 11377 7642 11401 7644
rect 11457 7642 11463 7644
rect 11217 7590 11219 7642
rect 11399 7590 11401 7642
rect 11155 7588 11161 7590
rect 11217 7588 11241 7590
rect 11297 7588 11321 7590
rect 11377 7588 11401 7590
rect 11457 7588 11463 7590
rect 11155 7579 11463 7588
rect 14973 7644 15281 7653
rect 14973 7642 14979 7644
rect 15035 7642 15059 7644
rect 15115 7642 15139 7644
rect 15195 7642 15219 7644
rect 15275 7642 15281 7644
rect 15035 7590 15037 7642
rect 15217 7590 15219 7642
rect 14973 7588 14979 7590
rect 15035 7588 15059 7590
rect 15115 7588 15139 7590
rect 15195 7588 15219 7590
rect 15275 7588 15281 7590
rect 14973 7579 15281 7588
rect 10495 7100 10803 7109
rect 10495 7098 10501 7100
rect 10557 7098 10581 7100
rect 10637 7098 10661 7100
rect 10717 7098 10741 7100
rect 10797 7098 10803 7100
rect 10557 7046 10559 7098
rect 10739 7046 10741 7098
rect 10495 7044 10501 7046
rect 10557 7044 10581 7046
rect 10637 7044 10661 7046
rect 10717 7044 10741 7046
rect 10797 7044 10803 7046
rect 10495 7035 10803 7044
rect 14313 7100 14621 7109
rect 14313 7098 14319 7100
rect 14375 7098 14399 7100
rect 14455 7098 14479 7100
rect 14535 7098 14559 7100
rect 14615 7098 14621 7100
rect 14375 7046 14377 7098
rect 14557 7046 14559 7098
rect 14313 7044 14319 7046
rect 14375 7044 14399 7046
rect 14455 7044 14479 7046
rect 14535 7044 14559 7046
rect 14615 7044 14621 7046
rect 14313 7035 14621 7044
rect 11155 6556 11463 6565
rect 11155 6554 11161 6556
rect 11217 6554 11241 6556
rect 11297 6554 11321 6556
rect 11377 6554 11401 6556
rect 11457 6554 11463 6556
rect 11217 6502 11219 6554
rect 11399 6502 11401 6554
rect 11155 6500 11161 6502
rect 11217 6500 11241 6502
rect 11297 6500 11321 6502
rect 11377 6500 11401 6502
rect 11457 6500 11463 6502
rect 11155 6491 11463 6500
rect 14973 6556 15281 6565
rect 14973 6554 14979 6556
rect 15035 6554 15059 6556
rect 15115 6554 15139 6556
rect 15195 6554 15219 6556
rect 15275 6554 15281 6556
rect 15035 6502 15037 6554
rect 15217 6502 15219 6554
rect 14973 6500 14979 6502
rect 15035 6500 15059 6502
rect 15115 6500 15139 6502
rect 15195 6500 15219 6502
rect 15275 6500 15281 6502
rect 14973 6491 15281 6500
rect 10495 6012 10803 6021
rect 10495 6010 10501 6012
rect 10557 6010 10581 6012
rect 10637 6010 10661 6012
rect 10717 6010 10741 6012
rect 10797 6010 10803 6012
rect 10557 5958 10559 6010
rect 10739 5958 10741 6010
rect 10495 5956 10501 5958
rect 10557 5956 10581 5958
rect 10637 5956 10661 5958
rect 10717 5956 10741 5958
rect 10797 5956 10803 5958
rect 10495 5947 10803 5956
rect 14313 6012 14621 6021
rect 14313 6010 14319 6012
rect 14375 6010 14399 6012
rect 14455 6010 14479 6012
rect 14535 6010 14559 6012
rect 14615 6010 14621 6012
rect 14375 5958 14377 6010
rect 14557 5958 14559 6010
rect 14313 5956 14319 5958
rect 14375 5956 14399 5958
rect 14455 5956 14479 5958
rect 14535 5956 14559 5958
rect 14615 5956 14621 5958
rect 14313 5947 14621 5956
rect 11155 5468 11463 5477
rect 11155 5466 11161 5468
rect 11217 5466 11241 5468
rect 11297 5466 11321 5468
rect 11377 5466 11401 5468
rect 11457 5466 11463 5468
rect 11217 5414 11219 5466
rect 11399 5414 11401 5466
rect 11155 5412 11161 5414
rect 11217 5412 11241 5414
rect 11297 5412 11321 5414
rect 11377 5412 11401 5414
rect 11457 5412 11463 5414
rect 11155 5403 11463 5412
rect 14973 5468 15281 5477
rect 14973 5466 14979 5468
rect 15035 5466 15059 5468
rect 15115 5466 15139 5468
rect 15195 5466 15219 5468
rect 15275 5466 15281 5468
rect 15035 5414 15037 5466
rect 15217 5414 15219 5466
rect 14973 5412 14979 5414
rect 15035 5412 15059 5414
rect 15115 5412 15139 5414
rect 15195 5412 15219 5414
rect 15275 5412 15281 5414
rect 14973 5403 15281 5412
rect 10495 4924 10803 4933
rect 10495 4922 10501 4924
rect 10557 4922 10581 4924
rect 10637 4922 10661 4924
rect 10717 4922 10741 4924
rect 10797 4922 10803 4924
rect 10557 4870 10559 4922
rect 10739 4870 10741 4922
rect 10495 4868 10501 4870
rect 10557 4868 10581 4870
rect 10637 4868 10661 4870
rect 10717 4868 10741 4870
rect 10797 4868 10803 4870
rect 10495 4859 10803 4868
rect 14313 4924 14621 4933
rect 14313 4922 14319 4924
rect 14375 4922 14399 4924
rect 14455 4922 14479 4924
rect 14535 4922 14559 4924
rect 14615 4922 14621 4924
rect 14375 4870 14377 4922
rect 14557 4870 14559 4922
rect 14313 4868 14319 4870
rect 14375 4868 14399 4870
rect 14455 4868 14479 4870
rect 14535 4868 14559 4870
rect 14615 4868 14621 4870
rect 14313 4859 14621 4868
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 9864 4480 9916 4486
rect 9864 4422 9916 4428
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 9876 4282 9904 4422
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10428 3534 10456 4014
rect 11072 3942 11100 4422
rect 11155 4380 11463 4389
rect 11155 4378 11161 4380
rect 11217 4378 11241 4380
rect 11297 4378 11321 4380
rect 11377 4378 11401 4380
rect 11457 4378 11463 4380
rect 11217 4326 11219 4378
rect 11399 4326 11401 4378
rect 11155 4324 11161 4326
rect 11217 4324 11241 4326
rect 11297 4324 11321 4326
rect 11377 4324 11401 4326
rect 11457 4324 11463 4326
rect 11155 4315 11463 4324
rect 14973 4380 15281 4389
rect 14973 4378 14979 4380
rect 15035 4378 15059 4380
rect 15115 4378 15139 4380
rect 15195 4378 15219 4380
rect 15275 4378 15281 4380
rect 15035 4326 15037 4378
rect 15217 4326 15219 4378
rect 14973 4324 14979 4326
rect 15035 4324 15059 4326
rect 15115 4324 15139 4326
rect 15195 4324 15219 4326
rect 15275 4324 15281 4326
rect 14973 4315 15281 4324
rect 15488 4214 15516 16934
rect 15476 4208 15528 4214
rect 15476 4150 15528 4156
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 10495 3836 10803 3845
rect 10495 3834 10501 3836
rect 10557 3834 10581 3836
rect 10637 3834 10661 3836
rect 10717 3834 10741 3836
rect 10797 3834 10803 3836
rect 10557 3782 10559 3834
rect 10739 3782 10741 3834
rect 10495 3780 10501 3782
rect 10557 3780 10581 3782
rect 10637 3780 10661 3782
rect 10717 3780 10741 3782
rect 10797 3780 10803 3782
rect 10495 3771 10803 3780
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 10428 3126 10456 3470
rect 10692 3392 10744 3398
rect 10692 3334 10744 3340
rect 10704 3194 10732 3334
rect 10692 3188 10744 3194
rect 11072 3176 11100 3878
rect 14313 3836 14621 3845
rect 14313 3834 14319 3836
rect 14375 3834 14399 3836
rect 14455 3834 14479 3836
rect 14535 3834 14559 3836
rect 14615 3834 14621 3836
rect 14375 3782 14377 3834
rect 14557 3782 14559 3834
rect 14313 3780 14319 3782
rect 14375 3780 14399 3782
rect 14455 3780 14479 3782
rect 14535 3780 14559 3782
rect 14615 3780 14621 3782
rect 14313 3771 14621 3780
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11155 3292 11463 3301
rect 11155 3290 11161 3292
rect 11217 3290 11241 3292
rect 11297 3290 11321 3292
rect 11377 3290 11401 3292
rect 11457 3290 11463 3292
rect 11217 3238 11219 3290
rect 11399 3238 11401 3290
rect 11155 3236 11161 3238
rect 11217 3236 11241 3238
rect 11297 3236 11321 3238
rect 11377 3236 11401 3238
rect 11457 3236 11463 3238
rect 11155 3227 11463 3236
rect 11072 3148 11192 3176
rect 10692 3130 10744 3136
rect 10416 3120 10468 3126
rect 10416 3062 10468 3068
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 9588 2508 9640 2514
rect 9588 2450 9640 2456
rect 5724 2304 5776 2310
rect 5724 2246 5776 2252
rect 7656 2304 7708 2310
rect 8392 2304 8444 2310
rect 7708 2252 7788 2258
rect 7656 2246 7788 2252
rect 8392 2246 8444 2252
rect 7668 2230 7788 2246
rect 7337 2204 7645 2213
rect 7337 2202 7343 2204
rect 7399 2202 7423 2204
rect 7479 2202 7503 2204
rect 7559 2202 7583 2204
rect 7639 2202 7645 2204
rect 7399 2150 7401 2202
rect 7581 2150 7583 2202
rect 7337 2148 7343 2150
rect 7399 2148 7423 2150
rect 7479 2148 7503 2150
rect 7559 2148 7583 2150
rect 7639 2148 7645 2150
rect 7337 2139 7645 2148
rect 7760 1170 7788 2230
rect 5552 1142 5672 1170
rect 7668 1142 7788 1170
rect 5552 800 5580 1142
rect 7668 800 7696 1142
rect 9784 800 9812 2790
rect 10495 2748 10803 2757
rect 10495 2746 10501 2748
rect 10557 2746 10581 2748
rect 10637 2746 10661 2748
rect 10717 2746 10741 2748
rect 10797 2746 10803 2748
rect 10557 2694 10559 2746
rect 10739 2694 10741 2746
rect 10495 2692 10501 2694
rect 10557 2692 10581 2694
rect 10637 2692 10661 2694
rect 10717 2692 10741 2694
rect 10797 2692 10803 2694
rect 10495 2683 10803 2692
rect 11072 2650 11100 2790
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11164 2446 11192 3148
rect 11520 2848 11572 2854
rect 11520 2790 11572 2796
rect 11532 2514 11560 2790
rect 11624 2650 11652 3470
rect 14973 3292 15281 3301
rect 14973 3290 14979 3292
rect 15035 3290 15059 3292
rect 15115 3290 15139 3292
rect 15195 3290 15219 3292
rect 15275 3290 15281 3292
rect 15035 3238 15037 3290
rect 15217 3238 15219 3290
rect 14973 3236 14979 3238
rect 15035 3236 15059 3238
rect 15115 3236 15139 3238
rect 15195 3236 15219 3238
rect 15275 3236 15281 3238
rect 14973 3227 15281 3236
rect 12072 2984 12124 2990
rect 12072 2926 12124 2932
rect 11612 2644 11664 2650
rect 11612 2586 11664 2592
rect 11520 2508 11572 2514
rect 11520 2450 11572 2456
rect 12084 2446 12112 2926
rect 14313 2748 14621 2757
rect 14313 2746 14319 2748
rect 14375 2746 14399 2748
rect 14455 2746 14479 2748
rect 14535 2746 14559 2748
rect 14615 2746 14621 2748
rect 14375 2694 14377 2746
rect 14557 2694 14559 2746
rect 14313 2692 14319 2694
rect 14375 2692 14399 2694
rect 14455 2692 14479 2694
rect 14535 2692 14559 2694
rect 14615 2692 14621 2694
rect 14313 2683 14621 2692
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 12072 2440 12124 2446
rect 12072 2382 12124 2388
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 14004 2304 14056 2310
rect 14004 2246 14056 2252
rect 11155 2204 11463 2213
rect 11155 2202 11161 2204
rect 11217 2202 11241 2204
rect 11297 2202 11321 2204
rect 11377 2202 11401 2204
rect 11457 2202 11463 2204
rect 11217 2150 11219 2202
rect 11399 2150 11401 2202
rect 11155 2148 11161 2150
rect 11217 2148 11241 2150
rect 11297 2148 11321 2150
rect 11377 2148 11401 2150
rect 11457 2148 11463 2150
rect 11155 2139 11463 2148
rect 11900 800 11928 2246
rect 14016 800 14044 2246
rect 14973 2204 15281 2213
rect 14973 2202 14979 2204
rect 15035 2202 15059 2204
rect 15115 2202 15139 2204
rect 15195 2202 15219 2204
rect 15275 2202 15281 2204
rect 15035 2150 15037 2202
rect 15217 2150 15219 2202
rect 14973 2148 14979 2150
rect 15035 2148 15059 2150
rect 15115 2148 15139 2150
rect 15195 2148 15219 2150
rect 15275 2148 15281 2150
rect 14973 2139 15281 2148
rect 16040 1306 16068 2382
rect 16040 1278 16160 1306
rect 16132 800 16160 1278
rect 1306 0 1362 800
rect 3422 0 3478 800
rect 5538 0 5594 800
rect 7654 0 7710 800
rect 9770 0 9826 800
rect 11886 0 11942 800
rect 14002 0 14058 800
rect 16118 0 16174 800
<< via2 >>
rect 3525 17434 3581 17436
rect 3605 17434 3661 17436
rect 3685 17434 3741 17436
rect 3765 17434 3821 17436
rect 3525 17382 3571 17434
rect 3571 17382 3581 17434
rect 3605 17382 3635 17434
rect 3635 17382 3647 17434
rect 3647 17382 3661 17434
rect 3685 17382 3699 17434
rect 3699 17382 3711 17434
rect 3711 17382 3741 17434
rect 3765 17382 3775 17434
rect 3775 17382 3821 17434
rect 3525 17380 3581 17382
rect 3605 17380 3661 17382
rect 3685 17380 3741 17382
rect 3765 17380 3821 17382
rect 2865 16890 2921 16892
rect 2945 16890 3001 16892
rect 3025 16890 3081 16892
rect 3105 16890 3161 16892
rect 2865 16838 2911 16890
rect 2911 16838 2921 16890
rect 2945 16838 2975 16890
rect 2975 16838 2987 16890
rect 2987 16838 3001 16890
rect 3025 16838 3039 16890
rect 3039 16838 3051 16890
rect 3051 16838 3081 16890
rect 3105 16838 3115 16890
rect 3115 16838 3161 16890
rect 2865 16836 2921 16838
rect 2945 16836 3001 16838
rect 3025 16836 3081 16838
rect 3105 16836 3161 16838
rect 3525 16346 3581 16348
rect 3605 16346 3661 16348
rect 3685 16346 3741 16348
rect 3765 16346 3821 16348
rect 3525 16294 3571 16346
rect 3571 16294 3581 16346
rect 3605 16294 3635 16346
rect 3635 16294 3647 16346
rect 3647 16294 3661 16346
rect 3685 16294 3699 16346
rect 3699 16294 3711 16346
rect 3711 16294 3741 16346
rect 3765 16294 3775 16346
rect 3775 16294 3821 16346
rect 3525 16292 3581 16294
rect 3605 16292 3661 16294
rect 3685 16292 3741 16294
rect 3765 16292 3821 16294
rect 2865 15802 2921 15804
rect 2945 15802 3001 15804
rect 3025 15802 3081 15804
rect 3105 15802 3161 15804
rect 2865 15750 2911 15802
rect 2911 15750 2921 15802
rect 2945 15750 2975 15802
rect 2975 15750 2987 15802
rect 2987 15750 3001 15802
rect 3025 15750 3039 15802
rect 3039 15750 3051 15802
rect 3051 15750 3081 15802
rect 3105 15750 3115 15802
rect 3115 15750 3161 15802
rect 2865 15748 2921 15750
rect 2945 15748 3001 15750
rect 3025 15748 3081 15750
rect 3105 15748 3161 15750
rect 7343 17434 7399 17436
rect 7423 17434 7479 17436
rect 7503 17434 7559 17436
rect 7583 17434 7639 17436
rect 7343 17382 7389 17434
rect 7389 17382 7399 17434
rect 7423 17382 7453 17434
rect 7453 17382 7465 17434
rect 7465 17382 7479 17434
rect 7503 17382 7517 17434
rect 7517 17382 7529 17434
rect 7529 17382 7559 17434
rect 7583 17382 7593 17434
rect 7593 17382 7639 17434
rect 7343 17380 7399 17382
rect 7423 17380 7479 17382
rect 7503 17380 7559 17382
rect 7583 17380 7639 17382
rect 11161 17434 11217 17436
rect 11241 17434 11297 17436
rect 11321 17434 11377 17436
rect 11401 17434 11457 17436
rect 11161 17382 11207 17434
rect 11207 17382 11217 17434
rect 11241 17382 11271 17434
rect 11271 17382 11283 17434
rect 11283 17382 11297 17434
rect 11321 17382 11335 17434
rect 11335 17382 11347 17434
rect 11347 17382 11377 17434
rect 11401 17382 11411 17434
rect 11411 17382 11457 17434
rect 11161 17380 11217 17382
rect 11241 17380 11297 17382
rect 11321 17380 11377 17382
rect 11401 17380 11457 17382
rect 14979 17434 15035 17436
rect 15059 17434 15115 17436
rect 15139 17434 15195 17436
rect 15219 17434 15275 17436
rect 14979 17382 15025 17434
rect 15025 17382 15035 17434
rect 15059 17382 15089 17434
rect 15089 17382 15101 17434
rect 15101 17382 15115 17434
rect 15139 17382 15153 17434
rect 15153 17382 15165 17434
rect 15165 17382 15195 17434
rect 15219 17382 15229 17434
rect 15229 17382 15275 17434
rect 14979 17380 15035 17382
rect 15059 17380 15115 17382
rect 15139 17380 15195 17382
rect 15219 17380 15275 17382
rect 6683 16890 6739 16892
rect 6763 16890 6819 16892
rect 6843 16890 6899 16892
rect 6923 16890 6979 16892
rect 6683 16838 6729 16890
rect 6729 16838 6739 16890
rect 6763 16838 6793 16890
rect 6793 16838 6805 16890
rect 6805 16838 6819 16890
rect 6843 16838 6857 16890
rect 6857 16838 6869 16890
rect 6869 16838 6899 16890
rect 6923 16838 6933 16890
rect 6933 16838 6979 16890
rect 6683 16836 6739 16838
rect 6763 16836 6819 16838
rect 6843 16836 6899 16838
rect 6923 16836 6979 16838
rect 7343 16346 7399 16348
rect 7423 16346 7479 16348
rect 7503 16346 7559 16348
rect 7583 16346 7639 16348
rect 7343 16294 7389 16346
rect 7389 16294 7399 16346
rect 7423 16294 7453 16346
rect 7453 16294 7465 16346
rect 7465 16294 7479 16346
rect 7503 16294 7517 16346
rect 7517 16294 7529 16346
rect 7529 16294 7559 16346
rect 7583 16294 7593 16346
rect 7593 16294 7639 16346
rect 7343 16292 7399 16294
rect 7423 16292 7479 16294
rect 7503 16292 7559 16294
rect 7583 16292 7639 16294
rect 6683 15802 6739 15804
rect 6763 15802 6819 15804
rect 6843 15802 6899 15804
rect 6923 15802 6979 15804
rect 6683 15750 6729 15802
rect 6729 15750 6739 15802
rect 6763 15750 6793 15802
rect 6793 15750 6805 15802
rect 6805 15750 6819 15802
rect 6843 15750 6857 15802
rect 6857 15750 6869 15802
rect 6869 15750 6899 15802
rect 6923 15750 6933 15802
rect 6933 15750 6979 15802
rect 6683 15748 6739 15750
rect 6763 15748 6819 15750
rect 6843 15748 6899 15750
rect 6923 15748 6979 15750
rect 3525 15258 3581 15260
rect 3605 15258 3661 15260
rect 3685 15258 3741 15260
rect 3765 15258 3821 15260
rect 3525 15206 3571 15258
rect 3571 15206 3581 15258
rect 3605 15206 3635 15258
rect 3635 15206 3647 15258
rect 3647 15206 3661 15258
rect 3685 15206 3699 15258
rect 3699 15206 3711 15258
rect 3711 15206 3741 15258
rect 3765 15206 3775 15258
rect 3775 15206 3821 15258
rect 3525 15204 3581 15206
rect 3605 15204 3661 15206
rect 3685 15204 3741 15206
rect 3765 15204 3821 15206
rect 2865 14714 2921 14716
rect 2945 14714 3001 14716
rect 3025 14714 3081 14716
rect 3105 14714 3161 14716
rect 2865 14662 2911 14714
rect 2911 14662 2921 14714
rect 2945 14662 2975 14714
rect 2975 14662 2987 14714
rect 2987 14662 3001 14714
rect 3025 14662 3039 14714
rect 3039 14662 3051 14714
rect 3051 14662 3081 14714
rect 3105 14662 3115 14714
rect 3115 14662 3161 14714
rect 2865 14660 2921 14662
rect 2945 14660 3001 14662
rect 3025 14660 3081 14662
rect 3105 14660 3161 14662
rect 6683 14714 6739 14716
rect 6763 14714 6819 14716
rect 6843 14714 6899 14716
rect 6923 14714 6979 14716
rect 6683 14662 6729 14714
rect 6729 14662 6739 14714
rect 6763 14662 6793 14714
rect 6793 14662 6805 14714
rect 6805 14662 6819 14714
rect 6843 14662 6857 14714
rect 6857 14662 6869 14714
rect 6869 14662 6899 14714
rect 6923 14662 6933 14714
rect 6933 14662 6979 14714
rect 6683 14660 6739 14662
rect 6763 14660 6819 14662
rect 6843 14660 6899 14662
rect 6923 14660 6979 14662
rect 3525 14170 3581 14172
rect 3605 14170 3661 14172
rect 3685 14170 3741 14172
rect 3765 14170 3821 14172
rect 3525 14118 3571 14170
rect 3571 14118 3581 14170
rect 3605 14118 3635 14170
rect 3635 14118 3647 14170
rect 3647 14118 3661 14170
rect 3685 14118 3699 14170
rect 3699 14118 3711 14170
rect 3711 14118 3741 14170
rect 3765 14118 3775 14170
rect 3775 14118 3821 14170
rect 3525 14116 3581 14118
rect 3605 14116 3661 14118
rect 3685 14116 3741 14118
rect 3765 14116 3821 14118
rect 2865 13626 2921 13628
rect 2945 13626 3001 13628
rect 3025 13626 3081 13628
rect 3105 13626 3161 13628
rect 2865 13574 2911 13626
rect 2911 13574 2921 13626
rect 2945 13574 2975 13626
rect 2975 13574 2987 13626
rect 2987 13574 3001 13626
rect 3025 13574 3039 13626
rect 3039 13574 3051 13626
rect 3051 13574 3081 13626
rect 3105 13574 3115 13626
rect 3115 13574 3161 13626
rect 2865 13572 2921 13574
rect 2945 13572 3001 13574
rect 3025 13572 3081 13574
rect 3105 13572 3161 13574
rect 6683 13626 6739 13628
rect 6763 13626 6819 13628
rect 6843 13626 6899 13628
rect 6923 13626 6979 13628
rect 6683 13574 6729 13626
rect 6729 13574 6739 13626
rect 6763 13574 6793 13626
rect 6793 13574 6805 13626
rect 6805 13574 6819 13626
rect 6843 13574 6857 13626
rect 6857 13574 6869 13626
rect 6869 13574 6899 13626
rect 6923 13574 6933 13626
rect 6933 13574 6979 13626
rect 6683 13572 6739 13574
rect 6763 13572 6819 13574
rect 6843 13572 6899 13574
rect 6923 13572 6979 13574
rect 3525 13082 3581 13084
rect 3605 13082 3661 13084
rect 3685 13082 3741 13084
rect 3765 13082 3821 13084
rect 3525 13030 3571 13082
rect 3571 13030 3581 13082
rect 3605 13030 3635 13082
rect 3635 13030 3647 13082
rect 3647 13030 3661 13082
rect 3685 13030 3699 13082
rect 3699 13030 3711 13082
rect 3711 13030 3741 13082
rect 3765 13030 3775 13082
rect 3775 13030 3821 13082
rect 3525 13028 3581 13030
rect 3605 13028 3661 13030
rect 3685 13028 3741 13030
rect 3765 13028 3821 13030
rect 2865 12538 2921 12540
rect 2945 12538 3001 12540
rect 3025 12538 3081 12540
rect 3105 12538 3161 12540
rect 2865 12486 2911 12538
rect 2911 12486 2921 12538
rect 2945 12486 2975 12538
rect 2975 12486 2987 12538
rect 2987 12486 3001 12538
rect 3025 12486 3039 12538
rect 3039 12486 3051 12538
rect 3051 12486 3081 12538
rect 3105 12486 3115 12538
rect 3115 12486 3161 12538
rect 2865 12484 2921 12486
rect 2945 12484 3001 12486
rect 3025 12484 3081 12486
rect 3105 12484 3161 12486
rect 6683 12538 6739 12540
rect 6763 12538 6819 12540
rect 6843 12538 6899 12540
rect 6923 12538 6979 12540
rect 6683 12486 6729 12538
rect 6729 12486 6739 12538
rect 6763 12486 6793 12538
rect 6793 12486 6805 12538
rect 6805 12486 6819 12538
rect 6843 12486 6857 12538
rect 6857 12486 6869 12538
rect 6869 12486 6899 12538
rect 6923 12486 6933 12538
rect 6933 12486 6979 12538
rect 6683 12484 6739 12486
rect 6763 12484 6819 12486
rect 6843 12484 6899 12486
rect 6923 12484 6979 12486
rect 3525 11994 3581 11996
rect 3605 11994 3661 11996
rect 3685 11994 3741 11996
rect 3765 11994 3821 11996
rect 3525 11942 3571 11994
rect 3571 11942 3581 11994
rect 3605 11942 3635 11994
rect 3635 11942 3647 11994
rect 3647 11942 3661 11994
rect 3685 11942 3699 11994
rect 3699 11942 3711 11994
rect 3711 11942 3741 11994
rect 3765 11942 3775 11994
rect 3775 11942 3821 11994
rect 3525 11940 3581 11942
rect 3605 11940 3661 11942
rect 3685 11940 3741 11942
rect 3765 11940 3821 11942
rect 2865 11450 2921 11452
rect 2945 11450 3001 11452
rect 3025 11450 3081 11452
rect 3105 11450 3161 11452
rect 2865 11398 2911 11450
rect 2911 11398 2921 11450
rect 2945 11398 2975 11450
rect 2975 11398 2987 11450
rect 2987 11398 3001 11450
rect 3025 11398 3039 11450
rect 3039 11398 3051 11450
rect 3051 11398 3081 11450
rect 3105 11398 3115 11450
rect 3115 11398 3161 11450
rect 2865 11396 2921 11398
rect 2945 11396 3001 11398
rect 3025 11396 3081 11398
rect 3105 11396 3161 11398
rect 6683 11450 6739 11452
rect 6763 11450 6819 11452
rect 6843 11450 6899 11452
rect 6923 11450 6979 11452
rect 6683 11398 6729 11450
rect 6729 11398 6739 11450
rect 6763 11398 6793 11450
rect 6793 11398 6805 11450
rect 6805 11398 6819 11450
rect 6843 11398 6857 11450
rect 6857 11398 6869 11450
rect 6869 11398 6899 11450
rect 6923 11398 6933 11450
rect 6933 11398 6979 11450
rect 6683 11396 6739 11398
rect 6763 11396 6819 11398
rect 6843 11396 6899 11398
rect 6923 11396 6979 11398
rect 3525 10906 3581 10908
rect 3605 10906 3661 10908
rect 3685 10906 3741 10908
rect 3765 10906 3821 10908
rect 3525 10854 3571 10906
rect 3571 10854 3581 10906
rect 3605 10854 3635 10906
rect 3635 10854 3647 10906
rect 3647 10854 3661 10906
rect 3685 10854 3699 10906
rect 3699 10854 3711 10906
rect 3711 10854 3741 10906
rect 3765 10854 3775 10906
rect 3775 10854 3821 10906
rect 3525 10852 3581 10854
rect 3605 10852 3661 10854
rect 3685 10852 3741 10854
rect 3765 10852 3821 10854
rect 2865 10362 2921 10364
rect 2945 10362 3001 10364
rect 3025 10362 3081 10364
rect 3105 10362 3161 10364
rect 2865 10310 2911 10362
rect 2911 10310 2921 10362
rect 2945 10310 2975 10362
rect 2975 10310 2987 10362
rect 2987 10310 3001 10362
rect 3025 10310 3039 10362
rect 3039 10310 3051 10362
rect 3051 10310 3081 10362
rect 3105 10310 3115 10362
rect 3115 10310 3161 10362
rect 2865 10308 2921 10310
rect 2945 10308 3001 10310
rect 3025 10308 3081 10310
rect 3105 10308 3161 10310
rect 6683 10362 6739 10364
rect 6763 10362 6819 10364
rect 6843 10362 6899 10364
rect 6923 10362 6979 10364
rect 6683 10310 6729 10362
rect 6729 10310 6739 10362
rect 6763 10310 6793 10362
rect 6793 10310 6805 10362
rect 6805 10310 6819 10362
rect 6843 10310 6857 10362
rect 6857 10310 6869 10362
rect 6869 10310 6899 10362
rect 6923 10310 6933 10362
rect 6933 10310 6979 10362
rect 6683 10308 6739 10310
rect 6763 10308 6819 10310
rect 6843 10308 6899 10310
rect 6923 10308 6979 10310
rect 3525 9818 3581 9820
rect 3605 9818 3661 9820
rect 3685 9818 3741 9820
rect 3765 9818 3821 9820
rect 3525 9766 3571 9818
rect 3571 9766 3581 9818
rect 3605 9766 3635 9818
rect 3635 9766 3647 9818
rect 3647 9766 3661 9818
rect 3685 9766 3699 9818
rect 3699 9766 3711 9818
rect 3711 9766 3741 9818
rect 3765 9766 3775 9818
rect 3775 9766 3821 9818
rect 3525 9764 3581 9766
rect 3605 9764 3661 9766
rect 3685 9764 3741 9766
rect 3765 9764 3821 9766
rect 2865 9274 2921 9276
rect 2945 9274 3001 9276
rect 3025 9274 3081 9276
rect 3105 9274 3161 9276
rect 2865 9222 2911 9274
rect 2911 9222 2921 9274
rect 2945 9222 2975 9274
rect 2975 9222 2987 9274
rect 2987 9222 3001 9274
rect 3025 9222 3039 9274
rect 3039 9222 3051 9274
rect 3051 9222 3081 9274
rect 3105 9222 3115 9274
rect 3115 9222 3161 9274
rect 2865 9220 2921 9222
rect 2945 9220 3001 9222
rect 3025 9220 3081 9222
rect 3105 9220 3161 9222
rect 6683 9274 6739 9276
rect 6763 9274 6819 9276
rect 6843 9274 6899 9276
rect 6923 9274 6979 9276
rect 6683 9222 6729 9274
rect 6729 9222 6739 9274
rect 6763 9222 6793 9274
rect 6793 9222 6805 9274
rect 6805 9222 6819 9274
rect 6843 9222 6857 9274
rect 6857 9222 6869 9274
rect 6869 9222 6899 9274
rect 6923 9222 6933 9274
rect 6933 9222 6979 9274
rect 6683 9220 6739 9222
rect 6763 9220 6819 9222
rect 6843 9220 6899 9222
rect 6923 9220 6979 9222
rect 3525 8730 3581 8732
rect 3605 8730 3661 8732
rect 3685 8730 3741 8732
rect 3765 8730 3821 8732
rect 3525 8678 3571 8730
rect 3571 8678 3581 8730
rect 3605 8678 3635 8730
rect 3635 8678 3647 8730
rect 3647 8678 3661 8730
rect 3685 8678 3699 8730
rect 3699 8678 3711 8730
rect 3711 8678 3741 8730
rect 3765 8678 3775 8730
rect 3775 8678 3821 8730
rect 3525 8676 3581 8678
rect 3605 8676 3661 8678
rect 3685 8676 3741 8678
rect 3765 8676 3821 8678
rect 2865 8186 2921 8188
rect 2945 8186 3001 8188
rect 3025 8186 3081 8188
rect 3105 8186 3161 8188
rect 2865 8134 2911 8186
rect 2911 8134 2921 8186
rect 2945 8134 2975 8186
rect 2975 8134 2987 8186
rect 2987 8134 3001 8186
rect 3025 8134 3039 8186
rect 3039 8134 3051 8186
rect 3051 8134 3081 8186
rect 3105 8134 3115 8186
rect 3115 8134 3161 8186
rect 2865 8132 2921 8134
rect 2945 8132 3001 8134
rect 3025 8132 3081 8134
rect 3105 8132 3161 8134
rect 6683 8186 6739 8188
rect 6763 8186 6819 8188
rect 6843 8186 6899 8188
rect 6923 8186 6979 8188
rect 6683 8134 6729 8186
rect 6729 8134 6739 8186
rect 6763 8134 6793 8186
rect 6793 8134 6805 8186
rect 6805 8134 6819 8186
rect 6843 8134 6857 8186
rect 6857 8134 6869 8186
rect 6869 8134 6899 8186
rect 6923 8134 6933 8186
rect 6933 8134 6979 8186
rect 6683 8132 6739 8134
rect 6763 8132 6819 8134
rect 6843 8132 6899 8134
rect 6923 8132 6979 8134
rect 3525 7642 3581 7644
rect 3605 7642 3661 7644
rect 3685 7642 3741 7644
rect 3765 7642 3821 7644
rect 3525 7590 3571 7642
rect 3571 7590 3581 7642
rect 3605 7590 3635 7642
rect 3635 7590 3647 7642
rect 3647 7590 3661 7642
rect 3685 7590 3699 7642
rect 3699 7590 3711 7642
rect 3711 7590 3741 7642
rect 3765 7590 3775 7642
rect 3775 7590 3821 7642
rect 3525 7588 3581 7590
rect 3605 7588 3661 7590
rect 3685 7588 3741 7590
rect 3765 7588 3821 7590
rect 2865 7098 2921 7100
rect 2945 7098 3001 7100
rect 3025 7098 3081 7100
rect 3105 7098 3161 7100
rect 2865 7046 2911 7098
rect 2911 7046 2921 7098
rect 2945 7046 2975 7098
rect 2975 7046 2987 7098
rect 2987 7046 3001 7098
rect 3025 7046 3039 7098
rect 3039 7046 3051 7098
rect 3051 7046 3081 7098
rect 3105 7046 3115 7098
rect 3115 7046 3161 7098
rect 2865 7044 2921 7046
rect 2945 7044 3001 7046
rect 3025 7044 3081 7046
rect 3105 7044 3161 7046
rect 6683 7098 6739 7100
rect 6763 7098 6819 7100
rect 6843 7098 6899 7100
rect 6923 7098 6979 7100
rect 6683 7046 6729 7098
rect 6729 7046 6739 7098
rect 6763 7046 6793 7098
rect 6793 7046 6805 7098
rect 6805 7046 6819 7098
rect 6843 7046 6857 7098
rect 6857 7046 6869 7098
rect 6869 7046 6899 7098
rect 6923 7046 6933 7098
rect 6933 7046 6979 7098
rect 6683 7044 6739 7046
rect 6763 7044 6819 7046
rect 6843 7044 6899 7046
rect 6923 7044 6979 7046
rect 3525 6554 3581 6556
rect 3605 6554 3661 6556
rect 3685 6554 3741 6556
rect 3765 6554 3821 6556
rect 3525 6502 3571 6554
rect 3571 6502 3581 6554
rect 3605 6502 3635 6554
rect 3635 6502 3647 6554
rect 3647 6502 3661 6554
rect 3685 6502 3699 6554
rect 3699 6502 3711 6554
rect 3711 6502 3741 6554
rect 3765 6502 3775 6554
rect 3775 6502 3821 6554
rect 3525 6500 3581 6502
rect 3605 6500 3661 6502
rect 3685 6500 3741 6502
rect 3765 6500 3821 6502
rect 2865 6010 2921 6012
rect 2945 6010 3001 6012
rect 3025 6010 3081 6012
rect 3105 6010 3161 6012
rect 2865 5958 2911 6010
rect 2911 5958 2921 6010
rect 2945 5958 2975 6010
rect 2975 5958 2987 6010
rect 2987 5958 3001 6010
rect 3025 5958 3039 6010
rect 3039 5958 3051 6010
rect 3051 5958 3081 6010
rect 3105 5958 3115 6010
rect 3115 5958 3161 6010
rect 2865 5956 2921 5958
rect 2945 5956 3001 5958
rect 3025 5956 3081 5958
rect 3105 5956 3161 5958
rect 6683 6010 6739 6012
rect 6763 6010 6819 6012
rect 6843 6010 6899 6012
rect 6923 6010 6979 6012
rect 6683 5958 6729 6010
rect 6729 5958 6739 6010
rect 6763 5958 6793 6010
rect 6793 5958 6805 6010
rect 6805 5958 6819 6010
rect 6843 5958 6857 6010
rect 6857 5958 6869 6010
rect 6869 5958 6899 6010
rect 6923 5958 6933 6010
rect 6933 5958 6979 6010
rect 6683 5956 6739 5958
rect 6763 5956 6819 5958
rect 6843 5956 6899 5958
rect 6923 5956 6979 5958
rect 3525 5466 3581 5468
rect 3605 5466 3661 5468
rect 3685 5466 3741 5468
rect 3765 5466 3821 5468
rect 3525 5414 3571 5466
rect 3571 5414 3581 5466
rect 3605 5414 3635 5466
rect 3635 5414 3647 5466
rect 3647 5414 3661 5466
rect 3685 5414 3699 5466
rect 3699 5414 3711 5466
rect 3711 5414 3741 5466
rect 3765 5414 3775 5466
rect 3775 5414 3821 5466
rect 3525 5412 3581 5414
rect 3605 5412 3661 5414
rect 3685 5412 3741 5414
rect 3765 5412 3821 5414
rect 2865 4922 2921 4924
rect 2945 4922 3001 4924
rect 3025 4922 3081 4924
rect 3105 4922 3161 4924
rect 2865 4870 2911 4922
rect 2911 4870 2921 4922
rect 2945 4870 2975 4922
rect 2975 4870 2987 4922
rect 2987 4870 3001 4922
rect 3025 4870 3039 4922
rect 3039 4870 3051 4922
rect 3051 4870 3081 4922
rect 3105 4870 3115 4922
rect 3115 4870 3161 4922
rect 2865 4868 2921 4870
rect 2945 4868 3001 4870
rect 3025 4868 3081 4870
rect 3105 4868 3161 4870
rect 3525 4378 3581 4380
rect 3605 4378 3661 4380
rect 3685 4378 3741 4380
rect 3765 4378 3821 4380
rect 3525 4326 3571 4378
rect 3571 4326 3581 4378
rect 3605 4326 3635 4378
rect 3635 4326 3647 4378
rect 3647 4326 3661 4378
rect 3685 4326 3699 4378
rect 3699 4326 3711 4378
rect 3711 4326 3741 4378
rect 3765 4326 3775 4378
rect 3775 4326 3821 4378
rect 3525 4324 3581 4326
rect 3605 4324 3661 4326
rect 3685 4324 3741 4326
rect 3765 4324 3821 4326
rect 2865 3834 2921 3836
rect 2945 3834 3001 3836
rect 3025 3834 3081 3836
rect 3105 3834 3161 3836
rect 2865 3782 2911 3834
rect 2911 3782 2921 3834
rect 2945 3782 2975 3834
rect 2975 3782 2987 3834
rect 2987 3782 3001 3834
rect 3025 3782 3039 3834
rect 3039 3782 3051 3834
rect 3051 3782 3081 3834
rect 3105 3782 3115 3834
rect 3115 3782 3161 3834
rect 2865 3780 2921 3782
rect 2945 3780 3001 3782
rect 3025 3780 3081 3782
rect 3105 3780 3161 3782
rect 3525 3290 3581 3292
rect 3605 3290 3661 3292
rect 3685 3290 3741 3292
rect 3765 3290 3821 3292
rect 3525 3238 3571 3290
rect 3571 3238 3581 3290
rect 3605 3238 3635 3290
rect 3635 3238 3647 3290
rect 3647 3238 3661 3290
rect 3685 3238 3699 3290
rect 3699 3238 3711 3290
rect 3711 3238 3741 3290
rect 3765 3238 3775 3290
rect 3775 3238 3821 3290
rect 3525 3236 3581 3238
rect 3605 3236 3661 3238
rect 3685 3236 3741 3238
rect 3765 3236 3821 3238
rect 2865 2746 2921 2748
rect 2945 2746 3001 2748
rect 3025 2746 3081 2748
rect 3105 2746 3161 2748
rect 2865 2694 2911 2746
rect 2911 2694 2921 2746
rect 2945 2694 2975 2746
rect 2975 2694 2987 2746
rect 2987 2694 3001 2746
rect 3025 2694 3039 2746
rect 3039 2694 3051 2746
rect 3051 2694 3081 2746
rect 3105 2694 3115 2746
rect 3115 2694 3161 2746
rect 2865 2692 2921 2694
rect 2945 2692 3001 2694
rect 3025 2692 3081 2694
rect 3105 2692 3161 2694
rect 6683 4922 6739 4924
rect 6763 4922 6819 4924
rect 6843 4922 6899 4924
rect 6923 4922 6979 4924
rect 6683 4870 6729 4922
rect 6729 4870 6739 4922
rect 6763 4870 6793 4922
rect 6793 4870 6805 4922
rect 6805 4870 6819 4922
rect 6843 4870 6857 4922
rect 6857 4870 6869 4922
rect 6869 4870 6899 4922
rect 6923 4870 6933 4922
rect 6933 4870 6979 4922
rect 6683 4868 6739 4870
rect 6763 4868 6819 4870
rect 6843 4868 6899 4870
rect 6923 4868 6979 4870
rect 3525 2202 3581 2204
rect 3605 2202 3661 2204
rect 3685 2202 3741 2204
rect 3765 2202 3821 2204
rect 3525 2150 3571 2202
rect 3571 2150 3581 2202
rect 3605 2150 3635 2202
rect 3635 2150 3647 2202
rect 3647 2150 3661 2202
rect 3685 2150 3699 2202
rect 3699 2150 3711 2202
rect 3711 2150 3741 2202
rect 3765 2150 3775 2202
rect 3775 2150 3821 2202
rect 3525 2148 3581 2150
rect 3605 2148 3661 2150
rect 3685 2148 3741 2150
rect 3765 2148 3821 2150
rect 6683 3834 6739 3836
rect 6763 3834 6819 3836
rect 6843 3834 6899 3836
rect 6923 3834 6979 3836
rect 6683 3782 6729 3834
rect 6729 3782 6739 3834
rect 6763 3782 6793 3834
rect 6793 3782 6805 3834
rect 6805 3782 6819 3834
rect 6843 3782 6857 3834
rect 6857 3782 6869 3834
rect 6869 3782 6899 3834
rect 6923 3782 6933 3834
rect 6933 3782 6979 3834
rect 6683 3780 6739 3782
rect 6763 3780 6819 3782
rect 6843 3780 6899 3782
rect 6923 3780 6979 3782
rect 7343 15258 7399 15260
rect 7423 15258 7479 15260
rect 7503 15258 7559 15260
rect 7583 15258 7639 15260
rect 7343 15206 7389 15258
rect 7389 15206 7399 15258
rect 7423 15206 7453 15258
rect 7453 15206 7465 15258
rect 7465 15206 7479 15258
rect 7503 15206 7517 15258
rect 7517 15206 7529 15258
rect 7529 15206 7559 15258
rect 7583 15206 7593 15258
rect 7593 15206 7639 15258
rect 7343 15204 7399 15206
rect 7423 15204 7479 15206
rect 7503 15204 7559 15206
rect 7583 15204 7639 15206
rect 7343 14170 7399 14172
rect 7423 14170 7479 14172
rect 7503 14170 7559 14172
rect 7583 14170 7639 14172
rect 7343 14118 7389 14170
rect 7389 14118 7399 14170
rect 7423 14118 7453 14170
rect 7453 14118 7465 14170
rect 7465 14118 7479 14170
rect 7503 14118 7517 14170
rect 7517 14118 7529 14170
rect 7529 14118 7559 14170
rect 7583 14118 7593 14170
rect 7593 14118 7639 14170
rect 7343 14116 7399 14118
rect 7423 14116 7479 14118
rect 7503 14116 7559 14118
rect 7583 14116 7639 14118
rect 7343 13082 7399 13084
rect 7423 13082 7479 13084
rect 7503 13082 7559 13084
rect 7583 13082 7639 13084
rect 7343 13030 7389 13082
rect 7389 13030 7399 13082
rect 7423 13030 7453 13082
rect 7453 13030 7465 13082
rect 7465 13030 7479 13082
rect 7503 13030 7517 13082
rect 7517 13030 7529 13082
rect 7529 13030 7559 13082
rect 7583 13030 7593 13082
rect 7593 13030 7639 13082
rect 7343 13028 7399 13030
rect 7423 13028 7479 13030
rect 7503 13028 7559 13030
rect 7583 13028 7639 13030
rect 7343 11994 7399 11996
rect 7423 11994 7479 11996
rect 7503 11994 7559 11996
rect 7583 11994 7639 11996
rect 7343 11942 7389 11994
rect 7389 11942 7399 11994
rect 7423 11942 7453 11994
rect 7453 11942 7465 11994
rect 7465 11942 7479 11994
rect 7503 11942 7517 11994
rect 7517 11942 7529 11994
rect 7529 11942 7559 11994
rect 7583 11942 7593 11994
rect 7593 11942 7639 11994
rect 7343 11940 7399 11942
rect 7423 11940 7479 11942
rect 7503 11940 7559 11942
rect 7583 11940 7639 11942
rect 7343 10906 7399 10908
rect 7423 10906 7479 10908
rect 7503 10906 7559 10908
rect 7583 10906 7639 10908
rect 7343 10854 7389 10906
rect 7389 10854 7399 10906
rect 7423 10854 7453 10906
rect 7453 10854 7465 10906
rect 7465 10854 7479 10906
rect 7503 10854 7517 10906
rect 7517 10854 7529 10906
rect 7529 10854 7559 10906
rect 7583 10854 7593 10906
rect 7593 10854 7639 10906
rect 7343 10852 7399 10854
rect 7423 10852 7479 10854
rect 7503 10852 7559 10854
rect 7583 10852 7639 10854
rect 7343 9818 7399 9820
rect 7423 9818 7479 9820
rect 7503 9818 7559 9820
rect 7583 9818 7639 9820
rect 7343 9766 7389 9818
rect 7389 9766 7399 9818
rect 7423 9766 7453 9818
rect 7453 9766 7465 9818
rect 7465 9766 7479 9818
rect 7503 9766 7517 9818
rect 7517 9766 7529 9818
rect 7529 9766 7559 9818
rect 7583 9766 7593 9818
rect 7593 9766 7639 9818
rect 7343 9764 7399 9766
rect 7423 9764 7479 9766
rect 7503 9764 7559 9766
rect 7583 9764 7639 9766
rect 7343 8730 7399 8732
rect 7423 8730 7479 8732
rect 7503 8730 7559 8732
rect 7583 8730 7639 8732
rect 7343 8678 7389 8730
rect 7389 8678 7399 8730
rect 7423 8678 7453 8730
rect 7453 8678 7465 8730
rect 7465 8678 7479 8730
rect 7503 8678 7517 8730
rect 7517 8678 7529 8730
rect 7529 8678 7559 8730
rect 7583 8678 7593 8730
rect 7593 8678 7639 8730
rect 7343 8676 7399 8678
rect 7423 8676 7479 8678
rect 7503 8676 7559 8678
rect 7583 8676 7639 8678
rect 7343 7642 7399 7644
rect 7423 7642 7479 7644
rect 7503 7642 7559 7644
rect 7583 7642 7639 7644
rect 7343 7590 7389 7642
rect 7389 7590 7399 7642
rect 7423 7590 7453 7642
rect 7453 7590 7465 7642
rect 7465 7590 7479 7642
rect 7503 7590 7517 7642
rect 7517 7590 7529 7642
rect 7529 7590 7559 7642
rect 7583 7590 7593 7642
rect 7593 7590 7639 7642
rect 7343 7588 7399 7590
rect 7423 7588 7479 7590
rect 7503 7588 7559 7590
rect 7583 7588 7639 7590
rect 7343 6554 7399 6556
rect 7423 6554 7479 6556
rect 7503 6554 7559 6556
rect 7583 6554 7639 6556
rect 7343 6502 7389 6554
rect 7389 6502 7399 6554
rect 7423 6502 7453 6554
rect 7453 6502 7465 6554
rect 7465 6502 7479 6554
rect 7503 6502 7517 6554
rect 7517 6502 7529 6554
rect 7529 6502 7559 6554
rect 7583 6502 7593 6554
rect 7593 6502 7639 6554
rect 7343 6500 7399 6502
rect 7423 6500 7479 6502
rect 7503 6500 7559 6502
rect 7583 6500 7639 6502
rect 7343 5466 7399 5468
rect 7423 5466 7479 5468
rect 7503 5466 7559 5468
rect 7583 5466 7639 5468
rect 7343 5414 7389 5466
rect 7389 5414 7399 5466
rect 7423 5414 7453 5466
rect 7453 5414 7465 5466
rect 7465 5414 7479 5466
rect 7503 5414 7517 5466
rect 7517 5414 7529 5466
rect 7529 5414 7559 5466
rect 7583 5414 7593 5466
rect 7593 5414 7639 5466
rect 7343 5412 7399 5414
rect 7423 5412 7479 5414
rect 7503 5412 7559 5414
rect 7583 5412 7639 5414
rect 7343 4378 7399 4380
rect 7423 4378 7479 4380
rect 7503 4378 7559 4380
rect 7583 4378 7639 4380
rect 7343 4326 7389 4378
rect 7389 4326 7399 4378
rect 7423 4326 7453 4378
rect 7453 4326 7465 4378
rect 7465 4326 7479 4378
rect 7503 4326 7517 4378
rect 7517 4326 7529 4378
rect 7529 4326 7559 4378
rect 7583 4326 7593 4378
rect 7593 4326 7639 4378
rect 7343 4324 7399 4326
rect 7423 4324 7479 4326
rect 7503 4324 7559 4326
rect 7583 4324 7639 4326
rect 6683 2746 6739 2748
rect 6763 2746 6819 2748
rect 6843 2746 6899 2748
rect 6923 2746 6979 2748
rect 6683 2694 6729 2746
rect 6729 2694 6739 2746
rect 6763 2694 6793 2746
rect 6793 2694 6805 2746
rect 6805 2694 6819 2746
rect 6843 2694 6857 2746
rect 6857 2694 6869 2746
rect 6869 2694 6899 2746
rect 6923 2694 6933 2746
rect 6933 2694 6979 2746
rect 6683 2692 6739 2694
rect 6763 2692 6819 2694
rect 6843 2692 6899 2694
rect 6923 2692 6979 2694
rect 7343 3290 7399 3292
rect 7423 3290 7479 3292
rect 7503 3290 7559 3292
rect 7583 3290 7639 3292
rect 7343 3238 7389 3290
rect 7389 3238 7399 3290
rect 7423 3238 7453 3290
rect 7453 3238 7465 3290
rect 7465 3238 7479 3290
rect 7503 3238 7517 3290
rect 7517 3238 7529 3290
rect 7529 3238 7559 3290
rect 7583 3238 7593 3290
rect 7593 3238 7639 3290
rect 7343 3236 7399 3238
rect 7423 3236 7479 3238
rect 7503 3236 7559 3238
rect 7583 3236 7639 3238
rect 10501 16890 10557 16892
rect 10581 16890 10637 16892
rect 10661 16890 10717 16892
rect 10741 16890 10797 16892
rect 10501 16838 10547 16890
rect 10547 16838 10557 16890
rect 10581 16838 10611 16890
rect 10611 16838 10623 16890
rect 10623 16838 10637 16890
rect 10661 16838 10675 16890
rect 10675 16838 10687 16890
rect 10687 16838 10717 16890
rect 10741 16838 10751 16890
rect 10751 16838 10797 16890
rect 10501 16836 10557 16838
rect 10581 16836 10637 16838
rect 10661 16836 10717 16838
rect 10741 16836 10797 16838
rect 14319 16890 14375 16892
rect 14399 16890 14455 16892
rect 14479 16890 14535 16892
rect 14559 16890 14615 16892
rect 14319 16838 14365 16890
rect 14365 16838 14375 16890
rect 14399 16838 14429 16890
rect 14429 16838 14441 16890
rect 14441 16838 14455 16890
rect 14479 16838 14493 16890
rect 14493 16838 14505 16890
rect 14505 16838 14535 16890
rect 14559 16838 14569 16890
rect 14569 16838 14615 16890
rect 14319 16836 14375 16838
rect 14399 16836 14455 16838
rect 14479 16836 14535 16838
rect 14559 16836 14615 16838
rect 11161 16346 11217 16348
rect 11241 16346 11297 16348
rect 11321 16346 11377 16348
rect 11401 16346 11457 16348
rect 11161 16294 11207 16346
rect 11207 16294 11217 16346
rect 11241 16294 11271 16346
rect 11271 16294 11283 16346
rect 11283 16294 11297 16346
rect 11321 16294 11335 16346
rect 11335 16294 11347 16346
rect 11347 16294 11377 16346
rect 11401 16294 11411 16346
rect 11411 16294 11457 16346
rect 11161 16292 11217 16294
rect 11241 16292 11297 16294
rect 11321 16292 11377 16294
rect 11401 16292 11457 16294
rect 14979 16346 15035 16348
rect 15059 16346 15115 16348
rect 15139 16346 15195 16348
rect 15219 16346 15275 16348
rect 14979 16294 15025 16346
rect 15025 16294 15035 16346
rect 15059 16294 15089 16346
rect 15089 16294 15101 16346
rect 15101 16294 15115 16346
rect 15139 16294 15153 16346
rect 15153 16294 15165 16346
rect 15165 16294 15195 16346
rect 15219 16294 15229 16346
rect 15229 16294 15275 16346
rect 14979 16292 15035 16294
rect 15059 16292 15115 16294
rect 15139 16292 15195 16294
rect 15219 16292 15275 16294
rect 10501 15802 10557 15804
rect 10581 15802 10637 15804
rect 10661 15802 10717 15804
rect 10741 15802 10797 15804
rect 10501 15750 10547 15802
rect 10547 15750 10557 15802
rect 10581 15750 10611 15802
rect 10611 15750 10623 15802
rect 10623 15750 10637 15802
rect 10661 15750 10675 15802
rect 10675 15750 10687 15802
rect 10687 15750 10717 15802
rect 10741 15750 10751 15802
rect 10751 15750 10797 15802
rect 10501 15748 10557 15750
rect 10581 15748 10637 15750
rect 10661 15748 10717 15750
rect 10741 15748 10797 15750
rect 14319 15802 14375 15804
rect 14399 15802 14455 15804
rect 14479 15802 14535 15804
rect 14559 15802 14615 15804
rect 14319 15750 14365 15802
rect 14365 15750 14375 15802
rect 14399 15750 14429 15802
rect 14429 15750 14441 15802
rect 14441 15750 14455 15802
rect 14479 15750 14493 15802
rect 14493 15750 14505 15802
rect 14505 15750 14535 15802
rect 14559 15750 14569 15802
rect 14569 15750 14615 15802
rect 14319 15748 14375 15750
rect 14399 15748 14455 15750
rect 14479 15748 14535 15750
rect 14559 15748 14615 15750
rect 11161 15258 11217 15260
rect 11241 15258 11297 15260
rect 11321 15258 11377 15260
rect 11401 15258 11457 15260
rect 11161 15206 11207 15258
rect 11207 15206 11217 15258
rect 11241 15206 11271 15258
rect 11271 15206 11283 15258
rect 11283 15206 11297 15258
rect 11321 15206 11335 15258
rect 11335 15206 11347 15258
rect 11347 15206 11377 15258
rect 11401 15206 11411 15258
rect 11411 15206 11457 15258
rect 11161 15204 11217 15206
rect 11241 15204 11297 15206
rect 11321 15204 11377 15206
rect 11401 15204 11457 15206
rect 14979 15258 15035 15260
rect 15059 15258 15115 15260
rect 15139 15258 15195 15260
rect 15219 15258 15275 15260
rect 14979 15206 15025 15258
rect 15025 15206 15035 15258
rect 15059 15206 15089 15258
rect 15089 15206 15101 15258
rect 15101 15206 15115 15258
rect 15139 15206 15153 15258
rect 15153 15206 15165 15258
rect 15165 15206 15195 15258
rect 15219 15206 15229 15258
rect 15229 15206 15275 15258
rect 14979 15204 15035 15206
rect 15059 15204 15115 15206
rect 15139 15204 15195 15206
rect 15219 15204 15275 15206
rect 10501 14714 10557 14716
rect 10581 14714 10637 14716
rect 10661 14714 10717 14716
rect 10741 14714 10797 14716
rect 10501 14662 10547 14714
rect 10547 14662 10557 14714
rect 10581 14662 10611 14714
rect 10611 14662 10623 14714
rect 10623 14662 10637 14714
rect 10661 14662 10675 14714
rect 10675 14662 10687 14714
rect 10687 14662 10717 14714
rect 10741 14662 10751 14714
rect 10751 14662 10797 14714
rect 10501 14660 10557 14662
rect 10581 14660 10637 14662
rect 10661 14660 10717 14662
rect 10741 14660 10797 14662
rect 14319 14714 14375 14716
rect 14399 14714 14455 14716
rect 14479 14714 14535 14716
rect 14559 14714 14615 14716
rect 14319 14662 14365 14714
rect 14365 14662 14375 14714
rect 14399 14662 14429 14714
rect 14429 14662 14441 14714
rect 14441 14662 14455 14714
rect 14479 14662 14493 14714
rect 14493 14662 14505 14714
rect 14505 14662 14535 14714
rect 14559 14662 14569 14714
rect 14569 14662 14615 14714
rect 14319 14660 14375 14662
rect 14399 14660 14455 14662
rect 14479 14660 14535 14662
rect 14559 14660 14615 14662
rect 11161 14170 11217 14172
rect 11241 14170 11297 14172
rect 11321 14170 11377 14172
rect 11401 14170 11457 14172
rect 11161 14118 11207 14170
rect 11207 14118 11217 14170
rect 11241 14118 11271 14170
rect 11271 14118 11283 14170
rect 11283 14118 11297 14170
rect 11321 14118 11335 14170
rect 11335 14118 11347 14170
rect 11347 14118 11377 14170
rect 11401 14118 11411 14170
rect 11411 14118 11457 14170
rect 11161 14116 11217 14118
rect 11241 14116 11297 14118
rect 11321 14116 11377 14118
rect 11401 14116 11457 14118
rect 14979 14170 15035 14172
rect 15059 14170 15115 14172
rect 15139 14170 15195 14172
rect 15219 14170 15275 14172
rect 14979 14118 15025 14170
rect 15025 14118 15035 14170
rect 15059 14118 15089 14170
rect 15089 14118 15101 14170
rect 15101 14118 15115 14170
rect 15139 14118 15153 14170
rect 15153 14118 15165 14170
rect 15165 14118 15195 14170
rect 15219 14118 15229 14170
rect 15229 14118 15275 14170
rect 14979 14116 15035 14118
rect 15059 14116 15115 14118
rect 15139 14116 15195 14118
rect 15219 14116 15275 14118
rect 10501 13626 10557 13628
rect 10581 13626 10637 13628
rect 10661 13626 10717 13628
rect 10741 13626 10797 13628
rect 10501 13574 10547 13626
rect 10547 13574 10557 13626
rect 10581 13574 10611 13626
rect 10611 13574 10623 13626
rect 10623 13574 10637 13626
rect 10661 13574 10675 13626
rect 10675 13574 10687 13626
rect 10687 13574 10717 13626
rect 10741 13574 10751 13626
rect 10751 13574 10797 13626
rect 10501 13572 10557 13574
rect 10581 13572 10637 13574
rect 10661 13572 10717 13574
rect 10741 13572 10797 13574
rect 14319 13626 14375 13628
rect 14399 13626 14455 13628
rect 14479 13626 14535 13628
rect 14559 13626 14615 13628
rect 14319 13574 14365 13626
rect 14365 13574 14375 13626
rect 14399 13574 14429 13626
rect 14429 13574 14441 13626
rect 14441 13574 14455 13626
rect 14479 13574 14493 13626
rect 14493 13574 14505 13626
rect 14505 13574 14535 13626
rect 14559 13574 14569 13626
rect 14569 13574 14615 13626
rect 14319 13572 14375 13574
rect 14399 13572 14455 13574
rect 14479 13572 14535 13574
rect 14559 13572 14615 13574
rect 11161 13082 11217 13084
rect 11241 13082 11297 13084
rect 11321 13082 11377 13084
rect 11401 13082 11457 13084
rect 11161 13030 11207 13082
rect 11207 13030 11217 13082
rect 11241 13030 11271 13082
rect 11271 13030 11283 13082
rect 11283 13030 11297 13082
rect 11321 13030 11335 13082
rect 11335 13030 11347 13082
rect 11347 13030 11377 13082
rect 11401 13030 11411 13082
rect 11411 13030 11457 13082
rect 11161 13028 11217 13030
rect 11241 13028 11297 13030
rect 11321 13028 11377 13030
rect 11401 13028 11457 13030
rect 14979 13082 15035 13084
rect 15059 13082 15115 13084
rect 15139 13082 15195 13084
rect 15219 13082 15275 13084
rect 14979 13030 15025 13082
rect 15025 13030 15035 13082
rect 15059 13030 15089 13082
rect 15089 13030 15101 13082
rect 15101 13030 15115 13082
rect 15139 13030 15153 13082
rect 15153 13030 15165 13082
rect 15165 13030 15195 13082
rect 15219 13030 15229 13082
rect 15229 13030 15275 13082
rect 14979 13028 15035 13030
rect 15059 13028 15115 13030
rect 15139 13028 15195 13030
rect 15219 13028 15275 13030
rect 10501 12538 10557 12540
rect 10581 12538 10637 12540
rect 10661 12538 10717 12540
rect 10741 12538 10797 12540
rect 10501 12486 10547 12538
rect 10547 12486 10557 12538
rect 10581 12486 10611 12538
rect 10611 12486 10623 12538
rect 10623 12486 10637 12538
rect 10661 12486 10675 12538
rect 10675 12486 10687 12538
rect 10687 12486 10717 12538
rect 10741 12486 10751 12538
rect 10751 12486 10797 12538
rect 10501 12484 10557 12486
rect 10581 12484 10637 12486
rect 10661 12484 10717 12486
rect 10741 12484 10797 12486
rect 14319 12538 14375 12540
rect 14399 12538 14455 12540
rect 14479 12538 14535 12540
rect 14559 12538 14615 12540
rect 14319 12486 14365 12538
rect 14365 12486 14375 12538
rect 14399 12486 14429 12538
rect 14429 12486 14441 12538
rect 14441 12486 14455 12538
rect 14479 12486 14493 12538
rect 14493 12486 14505 12538
rect 14505 12486 14535 12538
rect 14559 12486 14569 12538
rect 14569 12486 14615 12538
rect 14319 12484 14375 12486
rect 14399 12484 14455 12486
rect 14479 12484 14535 12486
rect 14559 12484 14615 12486
rect 11161 11994 11217 11996
rect 11241 11994 11297 11996
rect 11321 11994 11377 11996
rect 11401 11994 11457 11996
rect 11161 11942 11207 11994
rect 11207 11942 11217 11994
rect 11241 11942 11271 11994
rect 11271 11942 11283 11994
rect 11283 11942 11297 11994
rect 11321 11942 11335 11994
rect 11335 11942 11347 11994
rect 11347 11942 11377 11994
rect 11401 11942 11411 11994
rect 11411 11942 11457 11994
rect 11161 11940 11217 11942
rect 11241 11940 11297 11942
rect 11321 11940 11377 11942
rect 11401 11940 11457 11942
rect 14979 11994 15035 11996
rect 15059 11994 15115 11996
rect 15139 11994 15195 11996
rect 15219 11994 15275 11996
rect 14979 11942 15025 11994
rect 15025 11942 15035 11994
rect 15059 11942 15089 11994
rect 15089 11942 15101 11994
rect 15101 11942 15115 11994
rect 15139 11942 15153 11994
rect 15153 11942 15165 11994
rect 15165 11942 15195 11994
rect 15219 11942 15229 11994
rect 15229 11942 15275 11994
rect 14979 11940 15035 11942
rect 15059 11940 15115 11942
rect 15139 11940 15195 11942
rect 15219 11940 15275 11942
rect 10501 11450 10557 11452
rect 10581 11450 10637 11452
rect 10661 11450 10717 11452
rect 10741 11450 10797 11452
rect 10501 11398 10547 11450
rect 10547 11398 10557 11450
rect 10581 11398 10611 11450
rect 10611 11398 10623 11450
rect 10623 11398 10637 11450
rect 10661 11398 10675 11450
rect 10675 11398 10687 11450
rect 10687 11398 10717 11450
rect 10741 11398 10751 11450
rect 10751 11398 10797 11450
rect 10501 11396 10557 11398
rect 10581 11396 10637 11398
rect 10661 11396 10717 11398
rect 10741 11396 10797 11398
rect 14319 11450 14375 11452
rect 14399 11450 14455 11452
rect 14479 11450 14535 11452
rect 14559 11450 14615 11452
rect 14319 11398 14365 11450
rect 14365 11398 14375 11450
rect 14399 11398 14429 11450
rect 14429 11398 14441 11450
rect 14441 11398 14455 11450
rect 14479 11398 14493 11450
rect 14493 11398 14505 11450
rect 14505 11398 14535 11450
rect 14559 11398 14569 11450
rect 14569 11398 14615 11450
rect 14319 11396 14375 11398
rect 14399 11396 14455 11398
rect 14479 11396 14535 11398
rect 14559 11396 14615 11398
rect 11161 10906 11217 10908
rect 11241 10906 11297 10908
rect 11321 10906 11377 10908
rect 11401 10906 11457 10908
rect 11161 10854 11207 10906
rect 11207 10854 11217 10906
rect 11241 10854 11271 10906
rect 11271 10854 11283 10906
rect 11283 10854 11297 10906
rect 11321 10854 11335 10906
rect 11335 10854 11347 10906
rect 11347 10854 11377 10906
rect 11401 10854 11411 10906
rect 11411 10854 11457 10906
rect 11161 10852 11217 10854
rect 11241 10852 11297 10854
rect 11321 10852 11377 10854
rect 11401 10852 11457 10854
rect 14979 10906 15035 10908
rect 15059 10906 15115 10908
rect 15139 10906 15195 10908
rect 15219 10906 15275 10908
rect 14979 10854 15025 10906
rect 15025 10854 15035 10906
rect 15059 10854 15089 10906
rect 15089 10854 15101 10906
rect 15101 10854 15115 10906
rect 15139 10854 15153 10906
rect 15153 10854 15165 10906
rect 15165 10854 15195 10906
rect 15219 10854 15229 10906
rect 15229 10854 15275 10906
rect 14979 10852 15035 10854
rect 15059 10852 15115 10854
rect 15139 10852 15195 10854
rect 15219 10852 15275 10854
rect 10501 10362 10557 10364
rect 10581 10362 10637 10364
rect 10661 10362 10717 10364
rect 10741 10362 10797 10364
rect 10501 10310 10547 10362
rect 10547 10310 10557 10362
rect 10581 10310 10611 10362
rect 10611 10310 10623 10362
rect 10623 10310 10637 10362
rect 10661 10310 10675 10362
rect 10675 10310 10687 10362
rect 10687 10310 10717 10362
rect 10741 10310 10751 10362
rect 10751 10310 10797 10362
rect 10501 10308 10557 10310
rect 10581 10308 10637 10310
rect 10661 10308 10717 10310
rect 10741 10308 10797 10310
rect 14319 10362 14375 10364
rect 14399 10362 14455 10364
rect 14479 10362 14535 10364
rect 14559 10362 14615 10364
rect 14319 10310 14365 10362
rect 14365 10310 14375 10362
rect 14399 10310 14429 10362
rect 14429 10310 14441 10362
rect 14441 10310 14455 10362
rect 14479 10310 14493 10362
rect 14493 10310 14505 10362
rect 14505 10310 14535 10362
rect 14559 10310 14569 10362
rect 14569 10310 14615 10362
rect 14319 10308 14375 10310
rect 14399 10308 14455 10310
rect 14479 10308 14535 10310
rect 14559 10308 14615 10310
rect 11161 9818 11217 9820
rect 11241 9818 11297 9820
rect 11321 9818 11377 9820
rect 11401 9818 11457 9820
rect 11161 9766 11207 9818
rect 11207 9766 11217 9818
rect 11241 9766 11271 9818
rect 11271 9766 11283 9818
rect 11283 9766 11297 9818
rect 11321 9766 11335 9818
rect 11335 9766 11347 9818
rect 11347 9766 11377 9818
rect 11401 9766 11411 9818
rect 11411 9766 11457 9818
rect 11161 9764 11217 9766
rect 11241 9764 11297 9766
rect 11321 9764 11377 9766
rect 11401 9764 11457 9766
rect 14979 9818 15035 9820
rect 15059 9818 15115 9820
rect 15139 9818 15195 9820
rect 15219 9818 15275 9820
rect 14979 9766 15025 9818
rect 15025 9766 15035 9818
rect 15059 9766 15089 9818
rect 15089 9766 15101 9818
rect 15101 9766 15115 9818
rect 15139 9766 15153 9818
rect 15153 9766 15165 9818
rect 15165 9766 15195 9818
rect 15219 9766 15229 9818
rect 15229 9766 15275 9818
rect 14979 9764 15035 9766
rect 15059 9764 15115 9766
rect 15139 9764 15195 9766
rect 15219 9764 15275 9766
rect 10501 9274 10557 9276
rect 10581 9274 10637 9276
rect 10661 9274 10717 9276
rect 10741 9274 10797 9276
rect 10501 9222 10547 9274
rect 10547 9222 10557 9274
rect 10581 9222 10611 9274
rect 10611 9222 10623 9274
rect 10623 9222 10637 9274
rect 10661 9222 10675 9274
rect 10675 9222 10687 9274
rect 10687 9222 10717 9274
rect 10741 9222 10751 9274
rect 10751 9222 10797 9274
rect 10501 9220 10557 9222
rect 10581 9220 10637 9222
rect 10661 9220 10717 9222
rect 10741 9220 10797 9222
rect 14319 9274 14375 9276
rect 14399 9274 14455 9276
rect 14479 9274 14535 9276
rect 14559 9274 14615 9276
rect 14319 9222 14365 9274
rect 14365 9222 14375 9274
rect 14399 9222 14429 9274
rect 14429 9222 14441 9274
rect 14441 9222 14455 9274
rect 14479 9222 14493 9274
rect 14493 9222 14505 9274
rect 14505 9222 14535 9274
rect 14559 9222 14569 9274
rect 14569 9222 14615 9274
rect 14319 9220 14375 9222
rect 14399 9220 14455 9222
rect 14479 9220 14535 9222
rect 14559 9220 14615 9222
rect 11161 8730 11217 8732
rect 11241 8730 11297 8732
rect 11321 8730 11377 8732
rect 11401 8730 11457 8732
rect 11161 8678 11207 8730
rect 11207 8678 11217 8730
rect 11241 8678 11271 8730
rect 11271 8678 11283 8730
rect 11283 8678 11297 8730
rect 11321 8678 11335 8730
rect 11335 8678 11347 8730
rect 11347 8678 11377 8730
rect 11401 8678 11411 8730
rect 11411 8678 11457 8730
rect 11161 8676 11217 8678
rect 11241 8676 11297 8678
rect 11321 8676 11377 8678
rect 11401 8676 11457 8678
rect 14979 8730 15035 8732
rect 15059 8730 15115 8732
rect 15139 8730 15195 8732
rect 15219 8730 15275 8732
rect 14979 8678 15025 8730
rect 15025 8678 15035 8730
rect 15059 8678 15089 8730
rect 15089 8678 15101 8730
rect 15101 8678 15115 8730
rect 15139 8678 15153 8730
rect 15153 8678 15165 8730
rect 15165 8678 15195 8730
rect 15219 8678 15229 8730
rect 15229 8678 15275 8730
rect 14979 8676 15035 8678
rect 15059 8676 15115 8678
rect 15139 8676 15195 8678
rect 15219 8676 15275 8678
rect 10501 8186 10557 8188
rect 10581 8186 10637 8188
rect 10661 8186 10717 8188
rect 10741 8186 10797 8188
rect 10501 8134 10547 8186
rect 10547 8134 10557 8186
rect 10581 8134 10611 8186
rect 10611 8134 10623 8186
rect 10623 8134 10637 8186
rect 10661 8134 10675 8186
rect 10675 8134 10687 8186
rect 10687 8134 10717 8186
rect 10741 8134 10751 8186
rect 10751 8134 10797 8186
rect 10501 8132 10557 8134
rect 10581 8132 10637 8134
rect 10661 8132 10717 8134
rect 10741 8132 10797 8134
rect 14319 8186 14375 8188
rect 14399 8186 14455 8188
rect 14479 8186 14535 8188
rect 14559 8186 14615 8188
rect 14319 8134 14365 8186
rect 14365 8134 14375 8186
rect 14399 8134 14429 8186
rect 14429 8134 14441 8186
rect 14441 8134 14455 8186
rect 14479 8134 14493 8186
rect 14493 8134 14505 8186
rect 14505 8134 14535 8186
rect 14559 8134 14569 8186
rect 14569 8134 14615 8186
rect 14319 8132 14375 8134
rect 14399 8132 14455 8134
rect 14479 8132 14535 8134
rect 14559 8132 14615 8134
rect 11161 7642 11217 7644
rect 11241 7642 11297 7644
rect 11321 7642 11377 7644
rect 11401 7642 11457 7644
rect 11161 7590 11207 7642
rect 11207 7590 11217 7642
rect 11241 7590 11271 7642
rect 11271 7590 11283 7642
rect 11283 7590 11297 7642
rect 11321 7590 11335 7642
rect 11335 7590 11347 7642
rect 11347 7590 11377 7642
rect 11401 7590 11411 7642
rect 11411 7590 11457 7642
rect 11161 7588 11217 7590
rect 11241 7588 11297 7590
rect 11321 7588 11377 7590
rect 11401 7588 11457 7590
rect 14979 7642 15035 7644
rect 15059 7642 15115 7644
rect 15139 7642 15195 7644
rect 15219 7642 15275 7644
rect 14979 7590 15025 7642
rect 15025 7590 15035 7642
rect 15059 7590 15089 7642
rect 15089 7590 15101 7642
rect 15101 7590 15115 7642
rect 15139 7590 15153 7642
rect 15153 7590 15165 7642
rect 15165 7590 15195 7642
rect 15219 7590 15229 7642
rect 15229 7590 15275 7642
rect 14979 7588 15035 7590
rect 15059 7588 15115 7590
rect 15139 7588 15195 7590
rect 15219 7588 15275 7590
rect 10501 7098 10557 7100
rect 10581 7098 10637 7100
rect 10661 7098 10717 7100
rect 10741 7098 10797 7100
rect 10501 7046 10547 7098
rect 10547 7046 10557 7098
rect 10581 7046 10611 7098
rect 10611 7046 10623 7098
rect 10623 7046 10637 7098
rect 10661 7046 10675 7098
rect 10675 7046 10687 7098
rect 10687 7046 10717 7098
rect 10741 7046 10751 7098
rect 10751 7046 10797 7098
rect 10501 7044 10557 7046
rect 10581 7044 10637 7046
rect 10661 7044 10717 7046
rect 10741 7044 10797 7046
rect 14319 7098 14375 7100
rect 14399 7098 14455 7100
rect 14479 7098 14535 7100
rect 14559 7098 14615 7100
rect 14319 7046 14365 7098
rect 14365 7046 14375 7098
rect 14399 7046 14429 7098
rect 14429 7046 14441 7098
rect 14441 7046 14455 7098
rect 14479 7046 14493 7098
rect 14493 7046 14505 7098
rect 14505 7046 14535 7098
rect 14559 7046 14569 7098
rect 14569 7046 14615 7098
rect 14319 7044 14375 7046
rect 14399 7044 14455 7046
rect 14479 7044 14535 7046
rect 14559 7044 14615 7046
rect 11161 6554 11217 6556
rect 11241 6554 11297 6556
rect 11321 6554 11377 6556
rect 11401 6554 11457 6556
rect 11161 6502 11207 6554
rect 11207 6502 11217 6554
rect 11241 6502 11271 6554
rect 11271 6502 11283 6554
rect 11283 6502 11297 6554
rect 11321 6502 11335 6554
rect 11335 6502 11347 6554
rect 11347 6502 11377 6554
rect 11401 6502 11411 6554
rect 11411 6502 11457 6554
rect 11161 6500 11217 6502
rect 11241 6500 11297 6502
rect 11321 6500 11377 6502
rect 11401 6500 11457 6502
rect 14979 6554 15035 6556
rect 15059 6554 15115 6556
rect 15139 6554 15195 6556
rect 15219 6554 15275 6556
rect 14979 6502 15025 6554
rect 15025 6502 15035 6554
rect 15059 6502 15089 6554
rect 15089 6502 15101 6554
rect 15101 6502 15115 6554
rect 15139 6502 15153 6554
rect 15153 6502 15165 6554
rect 15165 6502 15195 6554
rect 15219 6502 15229 6554
rect 15229 6502 15275 6554
rect 14979 6500 15035 6502
rect 15059 6500 15115 6502
rect 15139 6500 15195 6502
rect 15219 6500 15275 6502
rect 10501 6010 10557 6012
rect 10581 6010 10637 6012
rect 10661 6010 10717 6012
rect 10741 6010 10797 6012
rect 10501 5958 10547 6010
rect 10547 5958 10557 6010
rect 10581 5958 10611 6010
rect 10611 5958 10623 6010
rect 10623 5958 10637 6010
rect 10661 5958 10675 6010
rect 10675 5958 10687 6010
rect 10687 5958 10717 6010
rect 10741 5958 10751 6010
rect 10751 5958 10797 6010
rect 10501 5956 10557 5958
rect 10581 5956 10637 5958
rect 10661 5956 10717 5958
rect 10741 5956 10797 5958
rect 14319 6010 14375 6012
rect 14399 6010 14455 6012
rect 14479 6010 14535 6012
rect 14559 6010 14615 6012
rect 14319 5958 14365 6010
rect 14365 5958 14375 6010
rect 14399 5958 14429 6010
rect 14429 5958 14441 6010
rect 14441 5958 14455 6010
rect 14479 5958 14493 6010
rect 14493 5958 14505 6010
rect 14505 5958 14535 6010
rect 14559 5958 14569 6010
rect 14569 5958 14615 6010
rect 14319 5956 14375 5958
rect 14399 5956 14455 5958
rect 14479 5956 14535 5958
rect 14559 5956 14615 5958
rect 11161 5466 11217 5468
rect 11241 5466 11297 5468
rect 11321 5466 11377 5468
rect 11401 5466 11457 5468
rect 11161 5414 11207 5466
rect 11207 5414 11217 5466
rect 11241 5414 11271 5466
rect 11271 5414 11283 5466
rect 11283 5414 11297 5466
rect 11321 5414 11335 5466
rect 11335 5414 11347 5466
rect 11347 5414 11377 5466
rect 11401 5414 11411 5466
rect 11411 5414 11457 5466
rect 11161 5412 11217 5414
rect 11241 5412 11297 5414
rect 11321 5412 11377 5414
rect 11401 5412 11457 5414
rect 14979 5466 15035 5468
rect 15059 5466 15115 5468
rect 15139 5466 15195 5468
rect 15219 5466 15275 5468
rect 14979 5414 15025 5466
rect 15025 5414 15035 5466
rect 15059 5414 15089 5466
rect 15089 5414 15101 5466
rect 15101 5414 15115 5466
rect 15139 5414 15153 5466
rect 15153 5414 15165 5466
rect 15165 5414 15195 5466
rect 15219 5414 15229 5466
rect 15229 5414 15275 5466
rect 14979 5412 15035 5414
rect 15059 5412 15115 5414
rect 15139 5412 15195 5414
rect 15219 5412 15275 5414
rect 10501 4922 10557 4924
rect 10581 4922 10637 4924
rect 10661 4922 10717 4924
rect 10741 4922 10797 4924
rect 10501 4870 10547 4922
rect 10547 4870 10557 4922
rect 10581 4870 10611 4922
rect 10611 4870 10623 4922
rect 10623 4870 10637 4922
rect 10661 4870 10675 4922
rect 10675 4870 10687 4922
rect 10687 4870 10717 4922
rect 10741 4870 10751 4922
rect 10751 4870 10797 4922
rect 10501 4868 10557 4870
rect 10581 4868 10637 4870
rect 10661 4868 10717 4870
rect 10741 4868 10797 4870
rect 14319 4922 14375 4924
rect 14399 4922 14455 4924
rect 14479 4922 14535 4924
rect 14559 4922 14615 4924
rect 14319 4870 14365 4922
rect 14365 4870 14375 4922
rect 14399 4870 14429 4922
rect 14429 4870 14441 4922
rect 14441 4870 14455 4922
rect 14479 4870 14493 4922
rect 14493 4870 14505 4922
rect 14505 4870 14535 4922
rect 14559 4870 14569 4922
rect 14569 4870 14615 4922
rect 14319 4868 14375 4870
rect 14399 4868 14455 4870
rect 14479 4868 14535 4870
rect 14559 4868 14615 4870
rect 11161 4378 11217 4380
rect 11241 4378 11297 4380
rect 11321 4378 11377 4380
rect 11401 4378 11457 4380
rect 11161 4326 11207 4378
rect 11207 4326 11217 4378
rect 11241 4326 11271 4378
rect 11271 4326 11283 4378
rect 11283 4326 11297 4378
rect 11321 4326 11335 4378
rect 11335 4326 11347 4378
rect 11347 4326 11377 4378
rect 11401 4326 11411 4378
rect 11411 4326 11457 4378
rect 11161 4324 11217 4326
rect 11241 4324 11297 4326
rect 11321 4324 11377 4326
rect 11401 4324 11457 4326
rect 14979 4378 15035 4380
rect 15059 4378 15115 4380
rect 15139 4378 15195 4380
rect 15219 4378 15275 4380
rect 14979 4326 15025 4378
rect 15025 4326 15035 4378
rect 15059 4326 15089 4378
rect 15089 4326 15101 4378
rect 15101 4326 15115 4378
rect 15139 4326 15153 4378
rect 15153 4326 15165 4378
rect 15165 4326 15195 4378
rect 15219 4326 15229 4378
rect 15229 4326 15275 4378
rect 14979 4324 15035 4326
rect 15059 4324 15115 4326
rect 15139 4324 15195 4326
rect 15219 4324 15275 4326
rect 10501 3834 10557 3836
rect 10581 3834 10637 3836
rect 10661 3834 10717 3836
rect 10741 3834 10797 3836
rect 10501 3782 10547 3834
rect 10547 3782 10557 3834
rect 10581 3782 10611 3834
rect 10611 3782 10623 3834
rect 10623 3782 10637 3834
rect 10661 3782 10675 3834
rect 10675 3782 10687 3834
rect 10687 3782 10717 3834
rect 10741 3782 10751 3834
rect 10751 3782 10797 3834
rect 10501 3780 10557 3782
rect 10581 3780 10637 3782
rect 10661 3780 10717 3782
rect 10741 3780 10797 3782
rect 14319 3834 14375 3836
rect 14399 3834 14455 3836
rect 14479 3834 14535 3836
rect 14559 3834 14615 3836
rect 14319 3782 14365 3834
rect 14365 3782 14375 3834
rect 14399 3782 14429 3834
rect 14429 3782 14441 3834
rect 14441 3782 14455 3834
rect 14479 3782 14493 3834
rect 14493 3782 14505 3834
rect 14505 3782 14535 3834
rect 14559 3782 14569 3834
rect 14569 3782 14615 3834
rect 14319 3780 14375 3782
rect 14399 3780 14455 3782
rect 14479 3780 14535 3782
rect 14559 3780 14615 3782
rect 11161 3290 11217 3292
rect 11241 3290 11297 3292
rect 11321 3290 11377 3292
rect 11401 3290 11457 3292
rect 11161 3238 11207 3290
rect 11207 3238 11217 3290
rect 11241 3238 11271 3290
rect 11271 3238 11283 3290
rect 11283 3238 11297 3290
rect 11321 3238 11335 3290
rect 11335 3238 11347 3290
rect 11347 3238 11377 3290
rect 11401 3238 11411 3290
rect 11411 3238 11457 3290
rect 11161 3236 11217 3238
rect 11241 3236 11297 3238
rect 11321 3236 11377 3238
rect 11401 3236 11457 3238
rect 7343 2202 7399 2204
rect 7423 2202 7479 2204
rect 7503 2202 7559 2204
rect 7583 2202 7639 2204
rect 7343 2150 7389 2202
rect 7389 2150 7399 2202
rect 7423 2150 7453 2202
rect 7453 2150 7465 2202
rect 7465 2150 7479 2202
rect 7503 2150 7517 2202
rect 7517 2150 7529 2202
rect 7529 2150 7559 2202
rect 7583 2150 7593 2202
rect 7593 2150 7639 2202
rect 7343 2148 7399 2150
rect 7423 2148 7479 2150
rect 7503 2148 7559 2150
rect 7583 2148 7639 2150
rect 10501 2746 10557 2748
rect 10581 2746 10637 2748
rect 10661 2746 10717 2748
rect 10741 2746 10797 2748
rect 10501 2694 10547 2746
rect 10547 2694 10557 2746
rect 10581 2694 10611 2746
rect 10611 2694 10623 2746
rect 10623 2694 10637 2746
rect 10661 2694 10675 2746
rect 10675 2694 10687 2746
rect 10687 2694 10717 2746
rect 10741 2694 10751 2746
rect 10751 2694 10797 2746
rect 10501 2692 10557 2694
rect 10581 2692 10637 2694
rect 10661 2692 10717 2694
rect 10741 2692 10797 2694
rect 14979 3290 15035 3292
rect 15059 3290 15115 3292
rect 15139 3290 15195 3292
rect 15219 3290 15275 3292
rect 14979 3238 15025 3290
rect 15025 3238 15035 3290
rect 15059 3238 15089 3290
rect 15089 3238 15101 3290
rect 15101 3238 15115 3290
rect 15139 3238 15153 3290
rect 15153 3238 15165 3290
rect 15165 3238 15195 3290
rect 15219 3238 15229 3290
rect 15229 3238 15275 3290
rect 14979 3236 15035 3238
rect 15059 3236 15115 3238
rect 15139 3236 15195 3238
rect 15219 3236 15275 3238
rect 14319 2746 14375 2748
rect 14399 2746 14455 2748
rect 14479 2746 14535 2748
rect 14559 2746 14615 2748
rect 14319 2694 14365 2746
rect 14365 2694 14375 2746
rect 14399 2694 14429 2746
rect 14429 2694 14441 2746
rect 14441 2694 14455 2746
rect 14479 2694 14493 2746
rect 14493 2694 14505 2746
rect 14505 2694 14535 2746
rect 14559 2694 14569 2746
rect 14569 2694 14615 2746
rect 14319 2692 14375 2694
rect 14399 2692 14455 2694
rect 14479 2692 14535 2694
rect 14559 2692 14615 2694
rect 11161 2202 11217 2204
rect 11241 2202 11297 2204
rect 11321 2202 11377 2204
rect 11401 2202 11457 2204
rect 11161 2150 11207 2202
rect 11207 2150 11217 2202
rect 11241 2150 11271 2202
rect 11271 2150 11283 2202
rect 11283 2150 11297 2202
rect 11321 2150 11335 2202
rect 11335 2150 11347 2202
rect 11347 2150 11377 2202
rect 11401 2150 11411 2202
rect 11411 2150 11457 2202
rect 11161 2148 11217 2150
rect 11241 2148 11297 2150
rect 11321 2148 11377 2150
rect 11401 2148 11457 2150
rect 14979 2202 15035 2204
rect 15059 2202 15115 2204
rect 15139 2202 15195 2204
rect 15219 2202 15275 2204
rect 14979 2150 15025 2202
rect 15025 2150 15035 2202
rect 15059 2150 15089 2202
rect 15089 2150 15101 2202
rect 15101 2150 15115 2202
rect 15139 2150 15153 2202
rect 15153 2150 15165 2202
rect 15165 2150 15195 2202
rect 15219 2150 15229 2202
rect 15229 2150 15275 2202
rect 14979 2148 15035 2150
rect 15059 2148 15115 2150
rect 15139 2148 15195 2150
rect 15219 2148 15275 2150
<< metal3 >>
rect 3515 17440 3831 17441
rect 3515 17376 3521 17440
rect 3585 17376 3601 17440
rect 3665 17376 3681 17440
rect 3745 17376 3761 17440
rect 3825 17376 3831 17440
rect 3515 17375 3831 17376
rect 7333 17440 7649 17441
rect 7333 17376 7339 17440
rect 7403 17376 7419 17440
rect 7483 17376 7499 17440
rect 7563 17376 7579 17440
rect 7643 17376 7649 17440
rect 7333 17375 7649 17376
rect 11151 17440 11467 17441
rect 11151 17376 11157 17440
rect 11221 17376 11237 17440
rect 11301 17376 11317 17440
rect 11381 17376 11397 17440
rect 11461 17376 11467 17440
rect 11151 17375 11467 17376
rect 14969 17440 15285 17441
rect 14969 17376 14975 17440
rect 15039 17376 15055 17440
rect 15119 17376 15135 17440
rect 15199 17376 15215 17440
rect 15279 17376 15285 17440
rect 14969 17375 15285 17376
rect 2855 16896 3171 16897
rect 2855 16832 2861 16896
rect 2925 16832 2941 16896
rect 3005 16832 3021 16896
rect 3085 16832 3101 16896
rect 3165 16832 3171 16896
rect 2855 16831 3171 16832
rect 6673 16896 6989 16897
rect 6673 16832 6679 16896
rect 6743 16832 6759 16896
rect 6823 16832 6839 16896
rect 6903 16832 6919 16896
rect 6983 16832 6989 16896
rect 6673 16831 6989 16832
rect 10491 16896 10807 16897
rect 10491 16832 10497 16896
rect 10561 16832 10577 16896
rect 10641 16832 10657 16896
rect 10721 16832 10737 16896
rect 10801 16832 10807 16896
rect 10491 16831 10807 16832
rect 14309 16896 14625 16897
rect 14309 16832 14315 16896
rect 14379 16832 14395 16896
rect 14459 16832 14475 16896
rect 14539 16832 14555 16896
rect 14619 16832 14625 16896
rect 14309 16831 14625 16832
rect 3515 16352 3831 16353
rect 3515 16288 3521 16352
rect 3585 16288 3601 16352
rect 3665 16288 3681 16352
rect 3745 16288 3761 16352
rect 3825 16288 3831 16352
rect 3515 16287 3831 16288
rect 7333 16352 7649 16353
rect 7333 16288 7339 16352
rect 7403 16288 7419 16352
rect 7483 16288 7499 16352
rect 7563 16288 7579 16352
rect 7643 16288 7649 16352
rect 7333 16287 7649 16288
rect 11151 16352 11467 16353
rect 11151 16288 11157 16352
rect 11221 16288 11237 16352
rect 11301 16288 11317 16352
rect 11381 16288 11397 16352
rect 11461 16288 11467 16352
rect 11151 16287 11467 16288
rect 14969 16352 15285 16353
rect 14969 16288 14975 16352
rect 15039 16288 15055 16352
rect 15119 16288 15135 16352
rect 15199 16288 15215 16352
rect 15279 16288 15285 16352
rect 14969 16287 15285 16288
rect 2855 15808 3171 15809
rect 2855 15744 2861 15808
rect 2925 15744 2941 15808
rect 3005 15744 3021 15808
rect 3085 15744 3101 15808
rect 3165 15744 3171 15808
rect 2855 15743 3171 15744
rect 6673 15808 6989 15809
rect 6673 15744 6679 15808
rect 6743 15744 6759 15808
rect 6823 15744 6839 15808
rect 6903 15744 6919 15808
rect 6983 15744 6989 15808
rect 6673 15743 6989 15744
rect 10491 15808 10807 15809
rect 10491 15744 10497 15808
rect 10561 15744 10577 15808
rect 10641 15744 10657 15808
rect 10721 15744 10737 15808
rect 10801 15744 10807 15808
rect 10491 15743 10807 15744
rect 14309 15808 14625 15809
rect 14309 15744 14315 15808
rect 14379 15744 14395 15808
rect 14459 15744 14475 15808
rect 14539 15744 14555 15808
rect 14619 15744 14625 15808
rect 14309 15743 14625 15744
rect 3515 15264 3831 15265
rect 3515 15200 3521 15264
rect 3585 15200 3601 15264
rect 3665 15200 3681 15264
rect 3745 15200 3761 15264
rect 3825 15200 3831 15264
rect 3515 15199 3831 15200
rect 7333 15264 7649 15265
rect 7333 15200 7339 15264
rect 7403 15200 7419 15264
rect 7483 15200 7499 15264
rect 7563 15200 7579 15264
rect 7643 15200 7649 15264
rect 7333 15199 7649 15200
rect 11151 15264 11467 15265
rect 11151 15200 11157 15264
rect 11221 15200 11237 15264
rect 11301 15200 11317 15264
rect 11381 15200 11397 15264
rect 11461 15200 11467 15264
rect 11151 15199 11467 15200
rect 14969 15264 15285 15265
rect 14969 15200 14975 15264
rect 15039 15200 15055 15264
rect 15119 15200 15135 15264
rect 15199 15200 15215 15264
rect 15279 15200 15285 15264
rect 14969 15199 15285 15200
rect 2855 14720 3171 14721
rect 2855 14656 2861 14720
rect 2925 14656 2941 14720
rect 3005 14656 3021 14720
rect 3085 14656 3101 14720
rect 3165 14656 3171 14720
rect 2855 14655 3171 14656
rect 6673 14720 6989 14721
rect 6673 14656 6679 14720
rect 6743 14656 6759 14720
rect 6823 14656 6839 14720
rect 6903 14656 6919 14720
rect 6983 14656 6989 14720
rect 6673 14655 6989 14656
rect 10491 14720 10807 14721
rect 10491 14656 10497 14720
rect 10561 14656 10577 14720
rect 10641 14656 10657 14720
rect 10721 14656 10737 14720
rect 10801 14656 10807 14720
rect 10491 14655 10807 14656
rect 14309 14720 14625 14721
rect 14309 14656 14315 14720
rect 14379 14656 14395 14720
rect 14459 14656 14475 14720
rect 14539 14656 14555 14720
rect 14619 14656 14625 14720
rect 14309 14655 14625 14656
rect 3515 14176 3831 14177
rect 3515 14112 3521 14176
rect 3585 14112 3601 14176
rect 3665 14112 3681 14176
rect 3745 14112 3761 14176
rect 3825 14112 3831 14176
rect 3515 14111 3831 14112
rect 7333 14176 7649 14177
rect 7333 14112 7339 14176
rect 7403 14112 7419 14176
rect 7483 14112 7499 14176
rect 7563 14112 7579 14176
rect 7643 14112 7649 14176
rect 7333 14111 7649 14112
rect 11151 14176 11467 14177
rect 11151 14112 11157 14176
rect 11221 14112 11237 14176
rect 11301 14112 11317 14176
rect 11381 14112 11397 14176
rect 11461 14112 11467 14176
rect 11151 14111 11467 14112
rect 14969 14176 15285 14177
rect 14969 14112 14975 14176
rect 15039 14112 15055 14176
rect 15119 14112 15135 14176
rect 15199 14112 15215 14176
rect 15279 14112 15285 14176
rect 14969 14111 15285 14112
rect 2855 13632 3171 13633
rect 2855 13568 2861 13632
rect 2925 13568 2941 13632
rect 3005 13568 3021 13632
rect 3085 13568 3101 13632
rect 3165 13568 3171 13632
rect 2855 13567 3171 13568
rect 6673 13632 6989 13633
rect 6673 13568 6679 13632
rect 6743 13568 6759 13632
rect 6823 13568 6839 13632
rect 6903 13568 6919 13632
rect 6983 13568 6989 13632
rect 6673 13567 6989 13568
rect 10491 13632 10807 13633
rect 10491 13568 10497 13632
rect 10561 13568 10577 13632
rect 10641 13568 10657 13632
rect 10721 13568 10737 13632
rect 10801 13568 10807 13632
rect 10491 13567 10807 13568
rect 14309 13632 14625 13633
rect 14309 13568 14315 13632
rect 14379 13568 14395 13632
rect 14459 13568 14475 13632
rect 14539 13568 14555 13632
rect 14619 13568 14625 13632
rect 14309 13567 14625 13568
rect 3515 13088 3831 13089
rect 3515 13024 3521 13088
rect 3585 13024 3601 13088
rect 3665 13024 3681 13088
rect 3745 13024 3761 13088
rect 3825 13024 3831 13088
rect 3515 13023 3831 13024
rect 7333 13088 7649 13089
rect 7333 13024 7339 13088
rect 7403 13024 7419 13088
rect 7483 13024 7499 13088
rect 7563 13024 7579 13088
rect 7643 13024 7649 13088
rect 7333 13023 7649 13024
rect 11151 13088 11467 13089
rect 11151 13024 11157 13088
rect 11221 13024 11237 13088
rect 11301 13024 11317 13088
rect 11381 13024 11397 13088
rect 11461 13024 11467 13088
rect 11151 13023 11467 13024
rect 14969 13088 15285 13089
rect 14969 13024 14975 13088
rect 15039 13024 15055 13088
rect 15119 13024 15135 13088
rect 15199 13024 15215 13088
rect 15279 13024 15285 13088
rect 14969 13023 15285 13024
rect 2855 12544 3171 12545
rect 2855 12480 2861 12544
rect 2925 12480 2941 12544
rect 3005 12480 3021 12544
rect 3085 12480 3101 12544
rect 3165 12480 3171 12544
rect 2855 12479 3171 12480
rect 6673 12544 6989 12545
rect 6673 12480 6679 12544
rect 6743 12480 6759 12544
rect 6823 12480 6839 12544
rect 6903 12480 6919 12544
rect 6983 12480 6989 12544
rect 6673 12479 6989 12480
rect 10491 12544 10807 12545
rect 10491 12480 10497 12544
rect 10561 12480 10577 12544
rect 10641 12480 10657 12544
rect 10721 12480 10737 12544
rect 10801 12480 10807 12544
rect 10491 12479 10807 12480
rect 14309 12544 14625 12545
rect 14309 12480 14315 12544
rect 14379 12480 14395 12544
rect 14459 12480 14475 12544
rect 14539 12480 14555 12544
rect 14619 12480 14625 12544
rect 14309 12479 14625 12480
rect 3515 12000 3831 12001
rect 3515 11936 3521 12000
rect 3585 11936 3601 12000
rect 3665 11936 3681 12000
rect 3745 11936 3761 12000
rect 3825 11936 3831 12000
rect 3515 11935 3831 11936
rect 7333 12000 7649 12001
rect 7333 11936 7339 12000
rect 7403 11936 7419 12000
rect 7483 11936 7499 12000
rect 7563 11936 7579 12000
rect 7643 11936 7649 12000
rect 7333 11935 7649 11936
rect 11151 12000 11467 12001
rect 11151 11936 11157 12000
rect 11221 11936 11237 12000
rect 11301 11936 11317 12000
rect 11381 11936 11397 12000
rect 11461 11936 11467 12000
rect 11151 11935 11467 11936
rect 14969 12000 15285 12001
rect 14969 11936 14975 12000
rect 15039 11936 15055 12000
rect 15119 11936 15135 12000
rect 15199 11936 15215 12000
rect 15279 11936 15285 12000
rect 14969 11935 15285 11936
rect 2855 11456 3171 11457
rect 2855 11392 2861 11456
rect 2925 11392 2941 11456
rect 3005 11392 3021 11456
rect 3085 11392 3101 11456
rect 3165 11392 3171 11456
rect 2855 11391 3171 11392
rect 6673 11456 6989 11457
rect 6673 11392 6679 11456
rect 6743 11392 6759 11456
rect 6823 11392 6839 11456
rect 6903 11392 6919 11456
rect 6983 11392 6989 11456
rect 6673 11391 6989 11392
rect 10491 11456 10807 11457
rect 10491 11392 10497 11456
rect 10561 11392 10577 11456
rect 10641 11392 10657 11456
rect 10721 11392 10737 11456
rect 10801 11392 10807 11456
rect 10491 11391 10807 11392
rect 14309 11456 14625 11457
rect 14309 11392 14315 11456
rect 14379 11392 14395 11456
rect 14459 11392 14475 11456
rect 14539 11392 14555 11456
rect 14619 11392 14625 11456
rect 14309 11391 14625 11392
rect 3515 10912 3831 10913
rect 3515 10848 3521 10912
rect 3585 10848 3601 10912
rect 3665 10848 3681 10912
rect 3745 10848 3761 10912
rect 3825 10848 3831 10912
rect 3515 10847 3831 10848
rect 7333 10912 7649 10913
rect 7333 10848 7339 10912
rect 7403 10848 7419 10912
rect 7483 10848 7499 10912
rect 7563 10848 7579 10912
rect 7643 10848 7649 10912
rect 7333 10847 7649 10848
rect 11151 10912 11467 10913
rect 11151 10848 11157 10912
rect 11221 10848 11237 10912
rect 11301 10848 11317 10912
rect 11381 10848 11397 10912
rect 11461 10848 11467 10912
rect 11151 10847 11467 10848
rect 14969 10912 15285 10913
rect 14969 10848 14975 10912
rect 15039 10848 15055 10912
rect 15119 10848 15135 10912
rect 15199 10848 15215 10912
rect 15279 10848 15285 10912
rect 14969 10847 15285 10848
rect 2855 10368 3171 10369
rect 2855 10304 2861 10368
rect 2925 10304 2941 10368
rect 3005 10304 3021 10368
rect 3085 10304 3101 10368
rect 3165 10304 3171 10368
rect 2855 10303 3171 10304
rect 6673 10368 6989 10369
rect 6673 10304 6679 10368
rect 6743 10304 6759 10368
rect 6823 10304 6839 10368
rect 6903 10304 6919 10368
rect 6983 10304 6989 10368
rect 6673 10303 6989 10304
rect 10491 10368 10807 10369
rect 10491 10304 10497 10368
rect 10561 10304 10577 10368
rect 10641 10304 10657 10368
rect 10721 10304 10737 10368
rect 10801 10304 10807 10368
rect 10491 10303 10807 10304
rect 14309 10368 14625 10369
rect 14309 10304 14315 10368
rect 14379 10304 14395 10368
rect 14459 10304 14475 10368
rect 14539 10304 14555 10368
rect 14619 10304 14625 10368
rect 14309 10303 14625 10304
rect 3515 9824 3831 9825
rect 3515 9760 3521 9824
rect 3585 9760 3601 9824
rect 3665 9760 3681 9824
rect 3745 9760 3761 9824
rect 3825 9760 3831 9824
rect 3515 9759 3831 9760
rect 7333 9824 7649 9825
rect 7333 9760 7339 9824
rect 7403 9760 7419 9824
rect 7483 9760 7499 9824
rect 7563 9760 7579 9824
rect 7643 9760 7649 9824
rect 7333 9759 7649 9760
rect 11151 9824 11467 9825
rect 11151 9760 11157 9824
rect 11221 9760 11237 9824
rect 11301 9760 11317 9824
rect 11381 9760 11397 9824
rect 11461 9760 11467 9824
rect 11151 9759 11467 9760
rect 14969 9824 15285 9825
rect 14969 9760 14975 9824
rect 15039 9760 15055 9824
rect 15119 9760 15135 9824
rect 15199 9760 15215 9824
rect 15279 9760 15285 9824
rect 14969 9759 15285 9760
rect 2855 9280 3171 9281
rect 2855 9216 2861 9280
rect 2925 9216 2941 9280
rect 3005 9216 3021 9280
rect 3085 9216 3101 9280
rect 3165 9216 3171 9280
rect 2855 9215 3171 9216
rect 6673 9280 6989 9281
rect 6673 9216 6679 9280
rect 6743 9216 6759 9280
rect 6823 9216 6839 9280
rect 6903 9216 6919 9280
rect 6983 9216 6989 9280
rect 6673 9215 6989 9216
rect 10491 9280 10807 9281
rect 10491 9216 10497 9280
rect 10561 9216 10577 9280
rect 10641 9216 10657 9280
rect 10721 9216 10737 9280
rect 10801 9216 10807 9280
rect 10491 9215 10807 9216
rect 14309 9280 14625 9281
rect 14309 9216 14315 9280
rect 14379 9216 14395 9280
rect 14459 9216 14475 9280
rect 14539 9216 14555 9280
rect 14619 9216 14625 9280
rect 14309 9215 14625 9216
rect 3515 8736 3831 8737
rect 3515 8672 3521 8736
rect 3585 8672 3601 8736
rect 3665 8672 3681 8736
rect 3745 8672 3761 8736
rect 3825 8672 3831 8736
rect 3515 8671 3831 8672
rect 7333 8736 7649 8737
rect 7333 8672 7339 8736
rect 7403 8672 7419 8736
rect 7483 8672 7499 8736
rect 7563 8672 7579 8736
rect 7643 8672 7649 8736
rect 7333 8671 7649 8672
rect 11151 8736 11467 8737
rect 11151 8672 11157 8736
rect 11221 8672 11237 8736
rect 11301 8672 11317 8736
rect 11381 8672 11397 8736
rect 11461 8672 11467 8736
rect 11151 8671 11467 8672
rect 14969 8736 15285 8737
rect 14969 8672 14975 8736
rect 15039 8672 15055 8736
rect 15119 8672 15135 8736
rect 15199 8672 15215 8736
rect 15279 8672 15285 8736
rect 14969 8671 15285 8672
rect 2855 8192 3171 8193
rect 2855 8128 2861 8192
rect 2925 8128 2941 8192
rect 3005 8128 3021 8192
rect 3085 8128 3101 8192
rect 3165 8128 3171 8192
rect 2855 8127 3171 8128
rect 6673 8192 6989 8193
rect 6673 8128 6679 8192
rect 6743 8128 6759 8192
rect 6823 8128 6839 8192
rect 6903 8128 6919 8192
rect 6983 8128 6989 8192
rect 6673 8127 6989 8128
rect 10491 8192 10807 8193
rect 10491 8128 10497 8192
rect 10561 8128 10577 8192
rect 10641 8128 10657 8192
rect 10721 8128 10737 8192
rect 10801 8128 10807 8192
rect 10491 8127 10807 8128
rect 14309 8192 14625 8193
rect 14309 8128 14315 8192
rect 14379 8128 14395 8192
rect 14459 8128 14475 8192
rect 14539 8128 14555 8192
rect 14619 8128 14625 8192
rect 14309 8127 14625 8128
rect 3515 7648 3831 7649
rect 3515 7584 3521 7648
rect 3585 7584 3601 7648
rect 3665 7584 3681 7648
rect 3745 7584 3761 7648
rect 3825 7584 3831 7648
rect 3515 7583 3831 7584
rect 7333 7648 7649 7649
rect 7333 7584 7339 7648
rect 7403 7584 7419 7648
rect 7483 7584 7499 7648
rect 7563 7584 7579 7648
rect 7643 7584 7649 7648
rect 7333 7583 7649 7584
rect 11151 7648 11467 7649
rect 11151 7584 11157 7648
rect 11221 7584 11237 7648
rect 11301 7584 11317 7648
rect 11381 7584 11397 7648
rect 11461 7584 11467 7648
rect 11151 7583 11467 7584
rect 14969 7648 15285 7649
rect 14969 7584 14975 7648
rect 15039 7584 15055 7648
rect 15119 7584 15135 7648
rect 15199 7584 15215 7648
rect 15279 7584 15285 7648
rect 14969 7583 15285 7584
rect 2855 7104 3171 7105
rect 2855 7040 2861 7104
rect 2925 7040 2941 7104
rect 3005 7040 3021 7104
rect 3085 7040 3101 7104
rect 3165 7040 3171 7104
rect 2855 7039 3171 7040
rect 6673 7104 6989 7105
rect 6673 7040 6679 7104
rect 6743 7040 6759 7104
rect 6823 7040 6839 7104
rect 6903 7040 6919 7104
rect 6983 7040 6989 7104
rect 6673 7039 6989 7040
rect 10491 7104 10807 7105
rect 10491 7040 10497 7104
rect 10561 7040 10577 7104
rect 10641 7040 10657 7104
rect 10721 7040 10737 7104
rect 10801 7040 10807 7104
rect 10491 7039 10807 7040
rect 14309 7104 14625 7105
rect 14309 7040 14315 7104
rect 14379 7040 14395 7104
rect 14459 7040 14475 7104
rect 14539 7040 14555 7104
rect 14619 7040 14625 7104
rect 14309 7039 14625 7040
rect 3515 6560 3831 6561
rect 3515 6496 3521 6560
rect 3585 6496 3601 6560
rect 3665 6496 3681 6560
rect 3745 6496 3761 6560
rect 3825 6496 3831 6560
rect 3515 6495 3831 6496
rect 7333 6560 7649 6561
rect 7333 6496 7339 6560
rect 7403 6496 7419 6560
rect 7483 6496 7499 6560
rect 7563 6496 7579 6560
rect 7643 6496 7649 6560
rect 7333 6495 7649 6496
rect 11151 6560 11467 6561
rect 11151 6496 11157 6560
rect 11221 6496 11237 6560
rect 11301 6496 11317 6560
rect 11381 6496 11397 6560
rect 11461 6496 11467 6560
rect 11151 6495 11467 6496
rect 14969 6560 15285 6561
rect 14969 6496 14975 6560
rect 15039 6496 15055 6560
rect 15119 6496 15135 6560
rect 15199 6496 15215 6560
rect 15279 6496 15285 6560
rect 14969 6495 15285 6496
rect 2855 6016 3171 6017
rect 2855 5952 2861 6016
rect 2925 5952 2941 6016
rect 3005 5952 3021 6016
rect 3085 5952 3101 6016
rect 3165 5952 3171 6016
rect 2855 5951 3171 5952
rect 6673 6016 6989 6017
rect 6673 5952 6679 6016
rect 6743 5952 6759 6016
rect 6823 5952 6839 6016
rect 6903 5952 6919 6016
rect 6983 5952 6989 6016
rect 6673 5951 6989 5952
rect 10491 6016 10807 6017
rect 10491 5952 10497 6016
rect 10561 5952 10577 6016
rect 10641 5952 10657 6016
rect 10721 5952 10737 6016
rect 10801 5952 10807 6016
rect 10491 5951 10807 5952
rect 14309 6016 14625 6017
rect 14309 5952 14315 6016
rect 14379 5952 14395 6016
rect 14459 5952 14475 6016
rect 14539 5952 14555 6016
rect 14619 5952 14625 6016
rect 14309 5951 14625 5952
rect 3515 5472 3831 5473
rect 3515 5408 3521 5472
rect 3585 5408 3601 5472
rect 3665 5408 3681 5472
rect 3745 5408 3761 5472
rect 3825 5408 3831 5472
rect 3515 5407 3831 5408
rect 7333 5472 7649 5473
rect 7333 5408 7339 5472
rect 7403 5408 7419 5472
rect 7483 5408 7499 5472
rect 7563 5408 7579 5472
rect 7643 5408 7649 5472
rect 7333 5407 7649 5408
rect 11151 5472 11467 5473
rect 11151 5408 11157 5472
rect 11221 5408 11237 5472
rect 11301 5408 11317 5472
rect 11381 5408 11397 5472
rect 11461 5408 11467 5472
rect 11151 5407 11467 5408
rect 14969 5472 15285 5473
rect 14969 5408 14975 5472
rect 15039 5408 15055 5472
rect 15119 5408 15135 5472
rect 15199 5408 15215 5472
rect 15279 5408 15285 5472
rect 14969 5407 15285 5408
rect 2855 4928 3171 4929
rect 2855 4864 2861 4928
rect 2925 4864 2941 4928
rect 3005 4864 3021 4928
rect 3085 4864 3101 4928
rect 3165 4864 3171 4928
rect 2855 4863 3171 4864
rect 6673 4928 6989 4929
rect 6673 4864 6679 4928
rect 6743 4864 6759 4928
rect 6823 4864 6839 4928
rect 6903 4864 6919 4928
rect 6983 4864 6989 4928
rect 6673 4863 6989 4864
rect 10491 4928 10807 4929
rect 10491 4864 10497 4928
rect 10561 4864 10577 4928
rect 10641 4864 10657 4928
rect 10721 4864 10737 4928
rect 10801 4864 10807 4928
rect 10491 4863 10807 4864
rect 14309 4928 14625 4929
rect 14309 4864 14315 4928
rect 14379 4864 14395 4928
rect 14459 4864 14475 4928
rect 14539 4864 14555 4928
rect 14619 4864 14625 4928
rect 14309 4863 14625 4864
rect 3515 4384 3831 4385
rect 3515 4320 3521 4384
rect 3585 4320 3601 4384
rect 3665 4320 3681 4384
rect 3745 4320 3761 4384
rect 3825 4320 3831 4384
rect 3515 4319 3831 4320
rect 7333 4384 7649 4385
rect 7333 4320 7339 4384
rect 7403 4320 7419 4384
rect 7483 4320 7499 4384
rect 7563 4320 7579 4384
rect 7643 4320 7649 4384
rect 7333 4319 7649 4320
rect 11151 4384 11467 4385
rect 11151 4320 11157 4384
rect 11221 4320 11237 4384
rect 11301 4320 11317 4384
rect 11381 4320 11397 4384
rect 11461 4320 11467 4384
rect 11151 4319 11467 4320
rect 14969 4384 15285 4385
rect 14969 4320 14975 4384
rect 15039 4320 15055 4384
rect 15119 4320 15135 4384
rect 15199 4320 15215 4384
rect 15279 4320 15285 4384
rect 14969 4319 15285 4320
rect 2855 3840 3171 3841
rect 2855 3776 2861 3840
rect 2925 3776 2941 3840
rect 3005 3776 3021 3840
rect 3085 3776 3101 3840
rect 3165 3776 3171 3840
rect 2855 3775 3171 3776
rect 6673 3840 6989 3841
rect 6673 3776 6679 3840
rect 6743 3776 6759 3840
rect 6823 3776 6839 3840
rect 6903 3776 6919 3840
rect 6983 3776 6989 3840
rect 6673 3775 6989 3776
rect 10491 3840 10807 3841
rect 10491 3776 10497 3840
rect 10561 3776 10577 3840
rect 10641 3776 10657 3840
rect 10721 3776 10737 3840
rect 10801 3776 10807 3840
rect 10491 3775 10807 3776
rect 14309 3840 14625 3841
rect 14309 3776 14315 3840
rect 14379 3776 14395 3840
rect 14459 3776 14475 3840
rect 14539 3776 14555 3840
rect 14619 3776 14625 3840
rect 14309 3775 14625 3776
rect 3515 3296 3831 3297
rect 3515 3232 3521 3296
rect 3585 3232 3601 3296
rect 3665 3232 3681 3296
rect 3745 3232 3761 3296
rect 3825 3232 3831 3296
rect 3515 3231 3831 3232
rect 7333 3296 7649 3297
rect 7333 3232 7339 3296
rect 7403 3232 7419 3296
rect 7483 3232 7499 3296
rect 7563 3232 7579 3296
rect 7643 3232 7649 3296
rect 7333 3231 7649 3232
rect 11151 3296 11467 3297
rect 11151 3232 11157 3296
rect 11221 3232 11237 3296
rect 11301 3232 11317 3296
rect 11381 3232 11397 3296
rect 11461 3232 11467 3296
rect 11151 3231 11467 3232
rect 14969 3296 15285 3297
rect 14969 3232 14975 3296
rect 15039 3232 15055 3296
rect 15119 3232 15135 3296
rect 15199 3232 15215 3296
rect 15279 3232 15285 3296
rect 14969 3231 15285 3232
rect 2855 2752 3171 2753
rect 2855 2688 2861 2752
rect 2925 2688 2941 2752
rect 3005 2688 3021 2752
rect 3085 2688 3101 2752
rect 3165 2688 3171 2752
rect 2855 2687 3171 2688
rect 6673 2752 6989 2753
rect 6673 2688 6679 2752
rect 6743 2688 6759 2752
rect 6823 2688 6839 2752
rect 6903 2688 6919 2752
rect 6983 2688 6989 2752
rect 6673 2687 6989 2688
rect 10491 2752 10807 2753
rect 10491 2688 10497 2752
rect 10561 2688 10577 2752
rect 10641 2688 10657 2752
rect 10721 2688 10737 2752
rect 10801 2688 10807 2752
rect 10491 2687 10807 2688
rect 14309 2752 14625 2753
rect 14309 2688 14315 2752
rect 14379 2688 14395 2752
rect 14459 2688 14475 2752
rect 14539 2688 14555 2752
rect 14619 2688 14625 2752
rect 14309 2687 14625 2688
rect 3515 2208 3831 2209
rect 3515 2144 3521 2208
rect 3585 2144 3601 2208
rect 3665 2144 3681 2208
rect 3745 2144 3761 2208
rect 3825 2144 3831 2208
rect 3515 2143 3831 2144
rect 7333 2208 7649 2209
rect 7333 2144 7339 2208
rect 7403 2144 7419 2208
rect 7483 2144 7499 2208
rect 7563 2144 7579 2208
rect 7643 2144 7649 2208
rect 7333 2143 7649 2144
rect 11151 2208 11467 2209
rect 11151 2144 11157 2208
rect 11221 2144 11237 2208
rect 11301 2144 11317 2208
rect 11381 2144 11397 2208
rect 11461 2144 11467 2208
rect 11151 2143 11467 2144
rect 14969 2208 15285 2209
rect 14969 2144 14975 2208
rect 15039 2144 15055 2208
rect 15119 2144 15135 2208
rect 15199 2144 15215 2208
rect 15279 2144 15285 2208
rect 14969 2143 15285 2144
<< via3 >>
rect 3521 17436 3585 17440
rect 3521 17380 3525 17436
rect 3525 17380 3581 17436
rect 3581 17380 3585 17436
rect 3521 17376 3585 17380
rect 3601 17436 3665 17440
rect 3601 17380 3605 17436
rect 3605 17380 3661 17436
rect 3661 17380 3665 17436
rect 3601 17376 3665 17380
rect 3681 17436 3745 17440
rect 3681 17380 3685 17436
rect 3685 17380 3741 17436
rect 3741 17380 3745 17436
rect 3681 17376 3745 17380
rect 3761 17436 3825 17440
rect 3761 17380 3765 17436
rect 3765 17380 3821 17436
rect 3821 17380 3825 17436
rect 3761 17376 3825 17380
rect 7339 17436 7403 17440
rect 7339 17380 7343 17436
rect 7343 17380 7399 17436
rect 7399 17380 7403 17436
rect 7339 17376 7403 17380
rect 7419 17436 7483 17440
rect 7419 17380 7423 17436
rect 7423 17380 7479 17436
rect 7479 17380 7483 17436
rect 7419 17376 7483 17380
rect 7499 17436 7563 17440
rect 7499 17380 7503 17436
rect 7503 17380 7559 17436
rect 7559 17380 7563 17436
rect 7499 17376 7563 17380
rect 7579 17436 7643 17440
rect 7579 17380 7583 17436
rect 7583 17380 7639 17436
rect 7639 17380 7643 17436
rect 7579 17376 7643 17380
rect 11157 17436 11221 17440
rect 11157 17380 11161 17436
rect 11161 17380 11217 17436
rect 11217 17380 11221 17436
rect 11157 17376 11221 17380
rect 11237 17436 11301 17440
rect 11237 17380 11241 17436
rect 11241 17380 11297 17436
rect 11297 17380 11301 17436
rect 11237 17376 11301 17380
rect 11317 17436 11381 17440
rect 11317 17380 11321 17436
rect 11321 17380 11377 17436
rect 11377 17380 11381 17436
rect 11317 17376 11381 17380
rect 11397 17436 11461 17440
rect 11397 17380 11401 17436
rect 11401 17380 11457 17436
rect 11457 17380 11461 17436
rect 11397 17376 11461 17380
rect 14975 17436 15039 17440
rect 14975 17380 14979 17436
rect 14979 17380 15035 17436
rect 15035 17380 15039 17436
rect 14975 17376 15039 17380
rect 15055 17436 15119 17440
rect 15055 17380 15059 17436
rect 15059 17380 15115 17436
rect 15115 17380 15119 17436
rect 15055 17376 15119 17380
rect 15135 17436 15199 17440
rect 15135 17380 15139 17436
rect 15139 17380 15195 17436
rect 15195 17380 15199 17436
rect 15135 17376 15199 17380
rect 15215 17436 15279 17440
rect 15215 17380 15219 17436
rect 15219 17380 15275 17436
rect 15275 17380 15279 17436
rect 15215 17376 15279 17380
rect 2861 16892 2925 16896
rect 2861 16836 2865 16892
rect 2865 16836 2921 16892
rect 2921 16836 2925 16892
rect 2861 16832 2925 16836
rect 2941 16892 3005 16896
rect 2941 16836 2945 16892
rect 2945 16836 3001 16892
rect 3001 16836 3005 16892
rect 2941 16832 3005 16836
rect 3021 16892 3085 16896
rect 3021 16836 3025 16892
rect 3025 16836 3081 16892
rect 3081 16836 3085 16892
rect 3021 16832 3085 16836
rect 3101 16892 3165 16896
rect 3101 16836 3105 16892
rect 3105 16836 3161 16892
rect 3161 16836 3165 16892
rect 3101 16832 3165 16836
rect 6679 16892 6743 16896
rect 6679 16836 6683 16892
rect 6683 16836 6739 16892
rect 6739 16836 6743 16892
rect 6679 16832 6743 16836
rect 6759 16892 6823 16896
rect 6759 16836 6763 16892
rect 6763 16836 6819 16892
rect 6819 16836 6823 16892
rect 6759 16832 6823 16836
rect 6839 16892 6903 16896
rect 6839 16836 6843 16892
rect 6843 16836 6899 16892
rect 6899 16836 6903 16892
rect 6839 16832 6903 16836
rect 6919 16892 6983 16896
rect 6919 16836 6923 16892
rect 6923 16836 6979 16892
rect 6979 16836 6983 16892
rect 6919 16832 6983 16836
rect 10497 16892 10561 16896
rect 10497 16836 10501 16892
rect 10501 16836 10557 16892
rect 10557 16836 10561 16892
rect 10497 16832 10561 16836
rect 10577 16892 10641 16896
rect 10577 16836 10581 16892
rect 10581 16836 10637 16892
rect 10637 16836 10641 16892
rect 10577 16832 10641 16836
rect 10657 16892 10721 16896
rect 10657 16836 10661 16892
rect 10661 16836 10717 16892
rect 10717 16836 10721 16892
rect 10657 16832 10721 16836
rect 10737 16892 10801 16896
rect 10737 16836 10741 16892
rect 10741 16836 10797 16892
rect 10797 16836 10801 16892
rect 10737 16832 10801 16836
rect 14315 16892 14379 16896
rect 14315 16836 14319 16892
rect 14319 16836 14375 16892
rect 14375 16836 14379 16892
rect 14315 16832 14379 16836
rect 14395 16892 14459 16896
rect 14395 16836 14399 16892
rect 14399 16836 14455 16892
rect 14455 16836 14459 16892
rect 14395 16832 14459 16836
rect 14475 16892 14539 16896
rect 14475 16836 14479 16892
rect 14479 16836 14535 16892
rect 14535 16836 14539 16892
rect 14475 16832 14539 16836
rect 14555 16892 14619 16896
rect 14555 16836 14559 16892
rect 14559 16836 14615 16892
rect 14615 16836 14619 16892
rect 14555 16832 14619 16836
rect 3521 16348 3585 16352
rect 3521 16292 3525 16348
rect 3525 16292 3581 16348
rect 3581 16292 3585 16348
rect 3521 16288 3585 16292
rect 3601 16348 3665 16352
rect 3601 16292 3605 16348
rect 3605 16292 3661 16348
rect 3661 16292 3665 16348
rect 3601 16288 3665 16292
rect 3681 16348 3745 16352
rect 3681 16292 3685 16348
rect 3685 16292 3741 16348
rect 3741 16292 3745 16348
rect 3681 16288 3745 16292
rect 3761 16348 3825 16352
rect 3761 16292 3765 16348
rect 3765 16292 3821 16348
rect 3821 16292 3825 16348
rect 3761 16288 3825 16292
rect 7339 16348 7403 16352
rect 7339 16292 7343 16348
rect 7343 16292 7399 16348
rect 7399 16292 7403 16348
rect 7339 16288 7403 16292
rect 7419 16348 7483 16352
rect 7419 16292 7423 16348
rect 7423 16292 7479 16348
rect 7479 16292 7483 16348
rect 7419 16288 7483 16292
rect 7499 16348 7563 16352
rect 7499 16292 7503 16348
rect 7503 16292 7559 16348
rect 7559 16292 7563 16348
rect 7499 16288 7563 16292
rect 7579 16348 7643 16352
rect 7579 16292 7583 16348
rect 7583 16292 7639 16348
rect 7639 16292 7643 16348
rect 7579 16288 7643 16292
rect 11157 16348 11221 16352
rect 11157 16292 11161 16348
rect 11161 16292 11217 16348
rect 11217 16292 11221 16348
rect 11157 16288 11221 16292
rect 11237 16348 11301 16352
rect 11237 16292 11241 16348
rect 11241 16292 11297 16348
rect 11297 16292 11301 16348
rect 11237 16288 11301 16292
rect 11317 16348 11381 16352
rect 11317 16292 11321 16348
rect 11321 16292 11377 16348
rect 11377 16292 11381 16348
rect 11317 16288 11381 16292
rect 11397 16348 11461 16352
rect 11397 16292 11401 16348
rect 11401 16292 11457 16348
rect 11457 16292 11461 16348
rect 11397 16288 11461 16292
rect 14975 16348 15039 16352
rect 14975 16292 14979 16348
rect 14979 16292 15035 16348
rect 15035 16292 15039 16348
rect 14975 16288 15039 16292
rect 15055 16348 15119 16352
rect 15055 16292 15059 16348
rect 15059 16292 15115 16348
rect 15115 16292 15119 16348
rect 15055 16288 15119 16292
rect 15135 16348 15199 16352
rect 15135 16292 15139 16348
rect 15139 16292 15195 16348
rect 15195 16292 15199 16348
rect 15135 16288 15199 16292
rect 15215 16348 15279 16352
rect 15215 16292 15219 16348
rect 15219 16292 15275 16348
rect 15275 16292 15279 16348
rect 15215 16288 15279 16292
rect 2861 15804 2925 15808
rect 2861 15748 2865 15804
rect 2865 15748 2921 15804
rect 2921 15748 2925 15804
rect 2861 15744 2925 15748
rect 2941 15804 3005 15808
rect 2941 15748 2945 15804
rect 2945 15748 3001 15804
rect 3001 15748 3005 15804
rect 2941 15744 3005 15748
rect 3021 15804 3085 15808
rect 3021 15748 3025 15804
rect 3025 15748 3081 15804
rect 3081 15748 3085 15804
rect 3021 15744 3085 15748
rect 3101 15804 3165 15808
rect 3101 15748 3105 15804
rect 3105 15748 3161 15804
rect 3161 15748 3165 15804
rect 3101 15744 3165 15748
rect 6679 15804 6743 15808
rect 6679 15748 6683 15804
rect 6683 15748 6739 15804
rect 6739 15748 6743 15804
rect 6679 15744 6743 15748
rect 6759 15804 6823 15808
rect 6759 15748 6763 15804
rect 6763 15748 6819 15804
rect 6819 15748 6823 15804
rect 6759 15744 6823 15748
rect 6839 15804 6903 15808
rect 6839 15748 6843 15804
rect 6843 15748 6899 15804
rect 6899 15748 6903 15804
rect 6839 15744 6903 15748
rect 6919 15804 6983 15808
rect 6919 15748 6923 15804
rect 6923 15748 6979 15804
rect 6979 15748 6983 15804
rect 6919 15744 6983 15748
rect 10497 15804 10561 15808
rect 10497 15748 10501 15804
rect 10501 15748 10557 15804
rect 10557 15748 10561 15804
rect 10497 15744 10561 15748
rect 10577 15804 10641 15808
rect 10577 15748 10581 15804
rect 10581 15748 10637 15804
rect 10637 15748 10641 15804
rect 10577 15744 10641 15748
rect 10657 15804 10721 15808
rect 10657 15748 10661 15804
rect 10661 15748 10717 15804
rect 10717 15748 10721 15804
rect 10657 15744 10721 15748
rect 10737 15804 10801 15808
rect 10737 15748 10741 15804
rect 10741 15748 10797 15804
rect 10797 15748 10801 15804
rect 10737 15744 10801 15748
rect 14315 15804 14379 15808
rect 14315 15748 14319 15804
rect 14319 15748 14375 15804
rect 14375 15748 14379 15804
rect 14315 15744 14379 15748
rect 14395 15804 14459 15808
rect 14395 15748 14399 15804
rect 14399 15748 14455 15804
rect 14455 15748 14459 15804
rect 14395 15744 14459 15748
rect 14475 15804 14539 15808
rect 14475 15748 14479 15804
rect 14479 15748 14535 15804
rect 14535 15748 14539 15804
rect 14475 15744 14539 15748
rect 14555 15804 14619 15808
rect 14555 15748 14559 15804
rect 14559 15748 14615 15804
rect 14615 15748 14619 15804
rect 14555 15744 14619 15748
rect 3521 15260 3585 15264
rect 3521 15204 3525 15260
rect 3525 15204 3581 15260
rect 3581 15204 3585 15260
rect 3521 15200 3585 15204
rect 3601 15260 3665 15264
rect 3601 15204 3605 15260
rect 3605 15204 3661 15260
rect 3661 15204 3665 15260
rect 3601 15200 3665 15204
rect 3681 15260 3745 15264
rect 3681 15204 3685 15260
rect 3685 15204 3741 15260
rect 3741 15204 3745 15260
rect 3681 15200 3745 15204
rect 3761 15260 3825 15264
rect 3761 15204 3765 15260
rect 3765 15204 3821 15260
rect 3821 15204 3825 15260
rect 3761 15200 3825 15204
rect 7339 15260 7403 15264
rect 7339 15204 7343 15260
rect 7343 15204 7399 15260
rect 7399 15204 7403 15260
rect 7339 15200 7403 15204
rect 7419 15260 7483 15264
rect 7419 15204 7423 15260
rect 7423 15204 7479 15260
rect 7479 15204 7483 15260
rect 7419 15200 7483 15204
rect 7499 15260 7563 15264
rect 7499 15204 7503 15260
rect 7503 15204 7559 15260
rect 7559 15204 7563 15260
rect 7499 15200 7563 15204
rect 7579 15260 7643 15264
rect 7579 15204 7583 15260
rect 7583 15204 7639 15260
rect 7639 15204 7643 15260
rect 7579 15200 7643 15204
rect 11157 15260 11221 15264
rect 11157 15204 11161 15260
rect 11161 15204 11217 15260
rect 11217 15204 11221 15260
rect 11157 15200 11221 15204
rect 11237 15260 11301 15264
rect 11237 15204 11241 15260
rect 11241 15204 11297 15260
rect 11297 15204 11301 15260
rect 11237 15200 11301 15204
rect 11317 15260 11381 15264
rect 11317 15204 11321 15260
rect 11321 15204 11377 15260
rect 11377 15204 11381 15260
rect 11317 15200 11381 15204
rect 11397 15260 11461 15264
rect 11397 15204 11401 15260
rect 11401 15204 11457 15260
rect 11457 15204 11461 15260
rect 11397 15200 11461 15204
rect 14975 15260 15039 15264
rect 14975 15204 14979 15260
rect 14979 15204 15035 15260
rect 15035 15204 15039 15260
rect 14975 15200 15039 15204
rect 15055 15260 15119 15264
rect 15055 15204 15059 15260
rect 15059 15204 15115 15260
rect 15115 15204 15119 15260
rect 15055 15200 15119 15204
rect 15135 15260 15199 15264
rect 15135 15204 15139 15260
rect 15139 15204 15195 15260
rect 15195 15204 15199 15260
rect 15135 15200 15199 15204
rect 15215 15260 15279 15264
rect 15215 15204 15219 15260
rect 15219 15204 15275 15260
rect 15275 15204 15279 15260
rect 15215 15200 15279 15204
rect 2861 14716 2925 14720
rect 2861 14660 2865 14716
rect 2865 14660 2921 14716
rect 2921 14660 2925 14716
rect 2861 14656 2925 14660
rect 2941 14716 3005 14720
rect 2941 14660 2945 14716
rect 2945 14660 3001 14716
rect 3001 14660 3005 14716
rect 2941 14656 3005 14660
rect 3021 14716 3085 14720
rect 3021 14660 3025 14716
rect 3025 14660 3081 14716
rect 3081 14660 3085 14716
rect 3021 14656 3085 14660
rect 3101 14716 3165 14720
rect 3101 14660 3105 14716
rect 3105 14660 3161 14716
rect 3161 14660 3165 14716
rect 3101 14656 3165 14660
rect 6679 14716 6743 14720
rect 6679 14660 6683 14716
rect 6683 14660 6739 14716
rect 6739 14660 6743 14716
rect 6679 14656 6743 14660
rect 6759 14716 6823 14720
rect 6759 14660 6763 14716
rect 6763 14660 6819 14716
rect 6819 14660 6823 14716
rect 6759 14656 6823 14660
rect 6839 14716 6903 14720
rect 6839 14660 6843 14716
rect 6843 14660 6899 14716
rect 6899 14660 6903 14716
rect 6839 14656 6903 14660
rect 6919 14716 6983 14720
rect 6919 14660 6923 14716
rect 6923 14660 6979 14716
rect 6979 14660 6983 14716
rect 6919 14656 6983 14660
rect 10497 14716 10561 14720
rect 10497 14660 10501 14716
rect 10501 14660 10557 14716
rect 10557 14660 10561 14716
rect 10497 14656 10561 14660
rect 10577 14716 10641 14720
rect 10577 14660 10581 14716
rect 10581 14660 10637 14716
rect 10637 14660 10641 14716
rect 10577 14656 10641 14660
rect 10657 14716 10721 14720
rect 10657 14660 10661 14716
rect 10661 14660 10717 14716
rect 10717 14660 10721 14716
rect 10657 14656 10721 14660
rect 10737 14716 10801 14720
rect 10737 14660 10741 14716
rect 10741 14660 10797 14716
rect 10797 14660 10801 14716
rect 10737 14656 10801 14660
rect 14315 14716 14379 14720
rect 14315 14660 14319 14716
rect 14319 14660 14375 14716
rect 14375 14660 14379 14716
rect 14315 14656 14379 14660
rect 14395 14716 14459 14720
rect 14395 14660 14399 14716
rect 14399 14660 14455 14716
rect 14455 14660 14459 14716
rect 14395 14656 14459 14660
rect 14475 14716 14539 14720
rect 14475 14660 14479 14716
rect 14479 14660 14535 14716
rect 14535 14660 14539 14716
rect 14475 14656 14539 14660
rect 14555 14716 14619 14720
rect 14555 14660 14559 14716
rect 14559 14660 14615 14716
rect 14615 14660 14619 14716
rect 14555 14656 14619 14660
rect 3521 14172 3585 14176
rect 3521 14116 3525 14172
rect 3525 14116 3581 14172
rect 3581 14116 3585 14172
rect 3521 14112 3585 14116
rect 3601 14172 3665 14176
rect 3601 14116 3605 14172
rect 3605 14116 3661 14172
rect 3661 14116 3665 14172
rect 3601 14112 3665 14116
rect 3681 14172 3745 14176
rect 3681 14116 3685 14172
rect 3685 14116 3741 14172
rect 3741 14116 3745 14172
rect 3681 14112 3745 14116
rect 3761 14172 3825 14176
rect 3761 14116 3765 14172
rect 3765 14116 3821 14172
rect 3821 14116 3825 14172
rect 3761 14112 3825 14116
rect 7339 14172 7403 14176
rect 7339 14116 7343 14172
rect 7343 14116 7399 14172
rect 7399 14116 7403 14172
rect 7339 14112 7403 14116
rect 7419 14172 7483 14176
rect 7419 14116 7423 14172
rect 7423 14116 7479 14172
rect 7479 14116 7483 14172
rect 7419 14112 7483 14116
rect 7499 14172 7563 14176
rect 7499 14116 7503 14172
rect 7503 14116 7559 14172
rect 7559 14116 7563 14172
rect 7499 14112 7563 14116
rect 7579 14172 7643 14176
rect 7579 14116 7583 14172
rect 7583 14116 7639 14172
rect 7639 14116 7643 14172
rect 7579 14112 7643 14116
rect 11157 14172 11221 14176
rect 11157 14116 11161 14172
rect 11161 14116 11217 14172
rect 11217 14116 11221 14172
rect 11157 14112 11221 14116
rect 11237 14172 11301 14176
rect 11237 14116 11241 14172
rect 11241 14116 11297 14172
rect 11297 14116 11301 14172
rect 11237 14112 11301 14116
rect 11317 14172 11381 14176
rect 11317 14116 11321 14172
rect 11321 14116 11377 14172
rect 11377 14116 11381 14172
rect 11317 14112 11381 14116
rect 11397 14172 11461 14176
rect 11397 14116 11401 14172
rect 11401 14116 11457 14172
rect 11457 14116 11461 14172
rect 11397 14112 11461 14116
rect 14975 14172 15039 14176
rect 14975 14116 14979 14172
rect 14979 14116 15035 14172
rect 15035 14116 15039 14172
rect 14975 14112 15039 14116
rect 15055 14172 15119 14176
rect 15055 14116 15059 14172
rect 15059 14116 15115 14172
rect 15115 14116 15119 14172
rect 15055 14112 15119 14116
rect 15135 14172 15199 14176
rect 15135 14116 15139 14172
rect 15139 14116 15195 14172
rect 15195 14116 15199 14172
rect 15135 14112 15199 14116
rect 15215 14172 15279 14176
rect 15215 14116 15219 14172
rect 15219 14116 15275 14172
rect 15275 14116 15279 14172
rect 15215 14112 15279 14116
rect 2861 13628 2925 13632
rect 2861 13572 2865 13628
rect 2865 13572 2921 13628
rect 2921 13572 2925 13628
rect 2861 13568 2925 13572
rect 2941 13628 3005 13632
rect 2941 13572 2945 13628
rect 2945 13572 3001 13628
rect 3001 13572 3005 13628
rect 2941 13568 3005 13572
rect 3021 13628 3085 13632
rect 3021 13572 3025 13628
rect 3025 13572 3081 13628
rect 3081 13572 3085 13628
rect 3021 13568 3085 13572
rect 3101 13628 3165 13632
rect 3101 13572 3105 13628
rect 3105 13572 3161 13628
rect 3161 13572 3165 13628
rect 3101 13568 3165 13572
rect 6679 13628 6743 13632
rect 6679 13572 6683 13628
rect 6683 13572 6739 13628
rect 6739 13572 6743 13628
rect 6679 13568 6743 13572
rect 6759 13628 6823 13632
rect 6759 13572 6763 13628
rect 6763 13572 6819 13628
rect 6819 13572 6823 13628
rect 6759 13568 6823 13572
rect 6839 13628 6903 13632
rect 6839 13572 6843 13628
rect 6843 13572 6899 13628
rect 6899 13572 6903 13628
rect 6839 13568 6903 13572
rect 6919 13628 6983 13632
rect 6919 13572 6923 13628
rect 6923 13572 6979 13628
rect 6979 13572 6983 13628
rect 6919 13568 6983 13572
rect 10497 13628 10561 13632
rect 10497 13572 10501 13628
rect 10501 13572 10557 13628
rect 10557 13572 10561 13628
rect 10497 13568 10561 13572
rect 10577 13628 10641 13632
rect 10577 13572 10581 13628
rect 10581 13572 10637 13628
rect 10637 13572 10641 13628
rect 10577 13568 10641 13572
rect 10657 13628 10721 13632
rect 10657 13572 10661 13628
rect 10661 13572 10717 13628
rect 10717 13572 10721 13628
rect 10657 13568 10721 13572
rect 10737 13628 10801 13632
rect 10737 13572 10741 13628
rect 10741 13572 10797 13628
rect 10797 13572 10801 13628
rect 10737 13568 10801 13572
rect 14315 13628 14379 13632
rect 14315 13572 14319 13628
rect 14319 13572 14375 13628
rect 14375 13572 14379 13628
rect 14315 13568 14379 13572
rect 14395 13628 14459 13632
rect 14395 13572 14399 13628
rect 14399 13572 14455 13628
rect 14455 13572 14459 13628
rect 14395 13568 14459 13572
rect 14475 13628 14539 13632
rect 14475 13572 14479 13628
rect 14479 13572 14535 13628
rect 14535 13572 14539 13628
rect 14475 13568 14539 13572
rect 14555 13628 14619 13632
rect 14555 13572 14559 13628
rect 14559 13572 14615 13628
rect 14615 13572 14619 13628
rect 14555 13568 14619 13572
rect 3521 13084 3585 13088
rect 3521 13028 3525 13084
rect 3525 13028 3581 13084
rect 3581 13028 3585 13084
rect 3521 13024 3585 13028
rect 3601 13084 3665 13088
rect 3601 13028 3605 13084
rect 3605 13028 3661 13084
rect 3661 13028 3665 13084
rect 3601 13024 3665 13028
rect 3681 13084 3745 13088
rect 3681 13028 3685 13084
rect 3685 13028 3741 13084
rect 3741 13028 3745 13084
rect 3681 13024 3745 13028
rect 3761 13084 3825 13088
rect 3761 13028 3765 13084
rect 3765 13028 3821 13084
rect 3821 13028 3825 13084
rect 3761 13024 3825 13028
rect 7339 13084 7403 13088
rect 7339 13028 7343 13084
rect 7343 13028 7399 13084
rect 7399 13028 7403 13084
rect 7339 13024 7403 13028
rect 7419 13084 7483 13088
rect 7419 13028 7423 13084
rect 7423 13028 7479 13084
rect 7479 13028 7483 13084
rect 7419 13024 7483 13028
rect 7499 13084 7563 13088
rect 7499 13028 7503 13084
rect 7503 13028 7559 13084
rect 7559 13028 7563 13084
rect 7499 13024 7563 13028
rect 7579 13084 7643 13088
rect 7579 13028 7583 13084
rect 7583 13028 7639 13084
rect 7639 13028 7643 13084
rect 7579 13024 7643 13028
rect 11157 13084 11221 13088
rect 11157 13028 11161 13084
rect 11161 13028 11217 13084
rect 11217 13028 11221 13084
rect 11157 13024 11221 13028
rect 11237 13084 11301 13088
rect 11237 13028 11241 13084
rect 11241 13028 11297 13084
rect 11297 13028 11301 13084
rect 11237 13024 11301 13028
rect 11317 13084 11381 13088
rect 11317 13028 11321 13084
rect 11321 13028 11377 13084
rect 11377 13028 11381 13084
rect 11317 13024 11381 13028
rect 11397 13084 11461 13088
rect 11397 13028 11401 13084
rect 11401 13028 11457 13084
rect 11457 13028 11461 13084
rect 11397 13024 11461 13028
rect 14975 13084 15039 13088
rect 14975 13028 14979 13084
rect 14979 13028 15035 13084
rect 15035 13028 15039 13084
rect 14975 13024 15039 13028
rect 15055 13084 15119 13088
rect 15055 13028 15059 13084
rect 15059 13028 15115 13084
rect 15115 13028 15119 13084
rect 15055 13024 15119 13028
rect 15135 13084 15199 13088
rect 15135 13028 15139 13084
rect 15139 13028 15195 13084
rect 15195 13028 15199 13084
rect 15135 13024 15199 13028
rect 15215 13084 15279 13088
rect 15215 13028 15219 13084
rect 15219 13028 15275 13084
rect 15275 13028 15279 13084
rect 15215 13024 15279 13028
rect 2861 12540 2925 12544
rect 2861 12484 2865 12540
rect 2865 12484 2921 12540
rect 2921 12484 2925 12540
rect 2861 12480 2925 12484
rect 2941 12540 3005 12544
rect 2941 12484 2945 12540
rect 2945 12484 3001 12540
rect 3001 12484 3005 12540
rect 2941 12480 3005 12484
rect 3021 12540 3085 12544
rect 3021 12484 3025 12540
rect 3025 12484 3081 12540
rect 3081 12484 3085 12540
rect 3021 12480 3085 12484
rect 3101 12540 3165 12544
rect 3101 12484 3105 12540
rect 3105 12484 3161 12540
rect 3161 12484 3165 12540
rect 3101 12480 3165 12484
rect 6679 12540 6743 12544
rect 6679 12484 6683 12540
rect 6683 12484 6739 12540
rect 6739 12484 6743 12540
rect 6679 12480 6743 12484
rect 6759 12540 6823 12544
rect 6759 12484 6763 12540
rect 6763 12484 6819 12540
rect 6819 12484 6823 12540
rect 6759 12480 6823 12484
rect 6839 12540 6903 12544
rect 6839 12484 6843 12540
rect 6843 12484 6899 12540
rect 6899 12484 6903 12540
rect 6839 12480 6903 12484
rect 6919 12540 6983 12544
rect 6919 12484 6923 12540
rect 6923 12484 6979 12540
rect 6979 12484 6983 12540
rect 6919 12480 6983 12484
rect 10497 12540 10561 12544
rect 10497 12484 10501 12540
rect 10501 12484 10557 12540
rect 10557 12484 10561 12540
rect 10497 12480 10561 12484
rect 10577 12540 10641 12544
rect 10577 12484 10581 12540
rect 10581 12484 10637 12540
rect 10637 12484 10641 12540
rect 10577 12480 10641 12484
rect 10657 12540 10721 12544
rect 10657 12484 10661 12540
rect 10661 12484 10717 12540
rect 10717 12484 10721 12540
rect 10657 12480 10721 12484
rect 10737 12540 10801 12544
rect 10737 12484 10741 12540
rect 10741 12484 10797 12540
rect 10797 12484 10801 12540
rect 10737 12480 10801 12484
rect 14315 12540 14379 12544
rect 14315 12484 14319 12540
rect 14319 12484 14375 12540
rect 14375 12484 14379 12540
rect 14315 12480 14379 12484
rect 14395 12540 14459 12544
rect 14395 12484 14399 12540
rect 14399 12484 14455 12540
rect 14455 12484 14459 12540
rect 14395 12480 14459 12484
rect 14475 12540 14539 12544
rect 14475 12484 14479 12540
rect 14479 12484 14535 12540
rect 14535 12484 14539 12540
rect 14475 12480 14539 12484
rect 14555 12540 14619 12544
rect 14555 12484 14559 12540
rect 14559 12484 14615 12540
rect 14615 12484 14619 12540
rect 14555 12480 14619 12484
rect 3521 11996 3585 12000
rect 3521 11940 3525 11996
rect 3525 11940 3581 11996
rect 3581 11940 3585 11996
rect 3521 11936 3585 11940
rect 3601 11996 3665 12000
rect 3601 11940 3605 11996
rect 3605 11940 3661 11996
rect 3661 11940 3665 11996
rect 3601 11936 3665 11940
rect 3681 11996 3745 12000
rect 3681 11940 3685 11996
rect 3685 11940 3741 11996
rect 3741 11940 3745 11996
rect 3681 11936 3745 11940
rect 3761 11996 3825 12000
rect 3761 11940 3765 11996
rect 3765 11940 3821 11996
rect 3821 11940 3825 11996
rect 3761 11936 3825 11940
rect 7339 11996 7403 12000
rect 7339 11940 7343 11996
rect 7343 11940 7399 11996
rect 7399 11940 7403 11996
rect 7339 11936 7403 11940
rect 7419 11996 7483 12000
rect 7419 11940 7423 11996
rect 7423 11940 7479 11996
rect 7479 11940 7483 11996
rect 7419 11936 7483 11940
rect 7499 11996 7563 12000
rect 7499 11940 7503 11996
rect 7503 11940 7559 11996
rect 7559 11940 7563 11996
rect 7499 11936 7563 11940
rect 7579 11996 7643 12000
rect 7579 11940 7583 11996
rect 7583 11940 7639 11996
rect 7639 11940 7643 11996
rect 7579 11936 7643 11940
rect 11157 11996 11221 12000
rect 11157 11940 11161 11996
rect 11161 11940 11217 11996
rect 11217 11940 11221 11996
rect 11157 11936 11221 11940
rect 11237 11996 11301 12000
rect 11237 11940 11241 11996
rect 11241 11940 11297 11996
rect 11297 11940 11301 11996
rect 11237 11936 11301 11940
rect 11317 11996 11381 12000
rect 11317 11940 11321 11996
rect 11321 11940 11377 11996
rect 11377 11940 11381 11996
rect 11317 11936 11381 11940
rect 11397 11996 11461 12000
rect 11397 11940 11401 11996
rect 11401 11940 11457 11996
rect 11457 11940 11461 11996
rect 11397 11936 11461 11940
rect 14975 11996 15039 12000
rect 14975 11940 14979 11996
rect 14979 11940 15035 11996
rect 15035 11940 15039 11996
rect 14975 11936 15039 11940
rect 15055 11996 15119 12000
rect 15055 11940 15059 11996
rect 15059 11940 15115 11996
rect 15115 11940 15119 11996
rect 15055 11936 15119 11940
rect 15135 11996 15199 12000
rect 15135 11940 15139 11996
rect 15139 11940 15195 11996
rect 15195 11940 15199 11996
rect 15135 11936 15199 11940
rect 15215 11996 15279 12000
rect 15215 11940 15219 11996
rect 15219 11940 15275 11996
rect 15275 11940 15279 11996
rect 15215 11936 15279 11940
rect 2861 11452 2925 11456
rect 2861 11396 2865 11452
rect 2865 11396 2921 11452
rect 2921 11396 2925 11452
rect 2861 11392 2925 11396
rect 2941 11452 3005 11456
rect 2941 11396 2945 11452
rect 2945 11396 3001 11452
rect 3001 11396 3005 11452
rect 2941 11392 3005 11396
rect 3021 11452 3085 11456
rect 3021 11396 3025 11452
rect 3025 11396 3081 11452
rect 3081 11396 3085 11452
rect 3021 11392 3085 11396
rect 3101 11452 3165 11456
rect 3101 11396 3105 11452
rect 3105 11396 3161 11452
rect 3161 11396 3165 11452
rect 3101 11392 3165 11396
rect 6679 11452 6743 11456
rect 6679 11396 6683 11452
rect 6683 11396 6739 11452
rect 6739 11396 6743 11452
rect 6679 11392 6743 11396
rect 6759 11452 6823 11456
rect 6759 11396 6763 11452
rect 6763 11396 6819 11452
rect 6819 11396 6823 11452
rect 6759 11392 6823 11396
rect 6839 11452 6903 11456
rect 6839 11396 6843 11452
rect 6843 11396 6899 11452
rect 6899 11396 6903 11452
rect 6839 11392 6903 11396
rect 6919 11452 6983 11456
rect 6919 11396 6923 11452
rect 6923 11396 6979 11452
rect 6979 11396 6983 11452
rect 6919 11392 6983 11396
rect 10497 11452 10561 11456
rect 10497 11396 10501 11452
rect 10501 11396 10557 11452
rect 10557 11396 10561 11452
rect 10497 11392 10561 11396
rect 10577 11452 10641 11456
rect 10577 11396 10581 11452
rect 10581 11396 10637 11452
rect 10637 11396 10641 11452
rect 10577 11392 10641 11396
rect 10657 11452 10721 11456
rect 10657 11396 10661 11452
rect 10661 11396 10717 11452
rect 10717 11396 10721 11452
rect 10657 11392 10721 11396
rect 10737 11452 10801 11456
rect 10737 11396 10741 11452
rect 10741 11396 10797 11452
rect 10797 11396 10801 11452
rect 10737 11392 10801 11396
rect 14315 11452 14379 11456
rect 14315 11396 14319 11452
rect 14319 11396 14375 11452
rect 14375 11396 14379 11452
rect 14315 11392 14379 11396
rect 14395 11452 14459 11456
rect 14395 11396 14399 11452
rect 14399 11396 14455 11452
rect 14455 11396 14459 11452
rect 14395 11392 14459 11396
rect 14475 11452 14539 11456
rect 14475 11396 14479 11452
rect 14479 11396 14535 11452
rect 14535 11396 14539 11452
rect 14475 11392 14539 11396
rect 14555 11452 14619 11456
rect 14555 11396 14559 11452
rect 14559 11396 14615 11452
rect 14615 11396 14619 11452
rect 14555 11392 14619 11396
rect 3521 10908 3585 10912
rect 3521 10852 3525 10908
rect 3525 10852 3581 10908
rect 3581 10852 3585 10908
rect 3521 10848 3585 10852
rect 3601 10908 3665 10912
rect 3601 10852 3605 10908
rect 3605 10852 3661 10908
rect 3661 10852 3665 10908
rect 3601 10848 3665 10852
rect 3681 10908 3745 10912
rect 3681 10852 3685 10908
rect 3685 10852 3741 10908
rect 3741 10852 3745 10908
rect 3681 10848 3745 10852
rect 3761 10908 3825 10912
rect 3761 10852 3765 10908
rect 3765 10852 3821 10908
rect 3821 10852 3825 10908
rect 3761 10848 3825 10852
rect 7339 10908 7403 10912
rect 7339 10852 7343 10908
rect 7343 10852 7399 10908
rect 7399 10852 7403 10908
rect 7339 10848 7403 10852
rect 7419 10908 7483 10912
rect 7419 10852 7423 10908
rect 7423 10852 7479 10908
rect 7479 10852 7483 10908
rect 7419 10848 7483 10852
rect 7499 10908 7563 10912
rect 7499 10852 7503 10908
rect 7503 10852 7559 10908
rect 7559 10852 7563 10908
rect 7499 10848 7563 10852
rect 7579 10908 7643 10912
rect 7579 10852 7583 10908
rect 7583 10852 7639 10908
rect 7639 10852 7643 10908
rect 7579 10848 7643 10852
rect 11157 10908 11221 10912
rect 11157 10852 11161 10908
rect 11161 10852 11217 10908
rect 11217 10852 11221 10908
rect 11157 10848 11221 10852
rect 11237 10908 11301 10912
rect 11237 10852 11241 10908
rect 11241 10852 11297 10908
rect 11297 10852 11301 10908
rect 11237 10848 11301 10852
rect 11317 10908 11381 10912
rect 11317 10852 11321 10908
rect 11321 10852 11377 10908
rect 11377 10852 11381 10908
rect 11317 10848 11381 10852
rect 11397 10908 11461 10912
rect 11397 10852 11401 10908
rect 11401 10852 11457 10908
rect 11457 10852 11461 10908
rect 11397 10848 11461 10852
rect 14975 10908 15039 10912
rect 14975 10852 14979 10908
rect 14979 10852 15035 10908
rect 15035 10852 15039 10908
rect 14975 10848 15039 10852
rect 15055 10908 15119 10912
rect 15055 10852 15059 10908
rect 15059 10852 15115 10908
rect 15115 10852 15119 10908
rect 15055 10848 15119 10852
rect 15135 10908 15199 10912
rect 15135 10852 15139 10908
rect 15139 10852 15195 10908
rect 15195 10852 15199 10908
rect 15135 10848 15199 10852
rect 15215 10908 15279 10912
rect 15215 10852 15219 10908
rect 15219 10852 15275 10908
rect 15275 10852 15279 10908
rect 15215 10848 15279 10852
rect 2861 10364 2925 10368
rect 2861 10308 2865 10364
rect 2865 10308 2921 10364
rect 2921 10308 2925 10364
rect 2861 10304 2925 10308
rect 2941 10364 3005 10368
rect 2941 10308 2945 10364
rect 2945 10308 3001 10364
rect 3001 10308 3005 10364
rect 2941 10304 3005 10308
rect 3021 10364 3085 10368
rect 3021 10308 3025 10364
rect 3025 10308 3081 10364
rect 3081 10308 3085 10364
rect 3021 10304 3085 10308
rect 3101 10364 3165 10368
rect 3101 10308 3105 10364
rect 3105 10308 3161 10364
rect 3161 10308 3165 10364
rect 3101 10304 3165 10308
rect 6679 10364 6743 10368
rect 6679 10308 6683 10364
rect 6683 10308 6739 10364
rect 6739 10308 6743 10364
rect 6679 10304 6743 10308
rect 6759 10364 6823 10368
rect 6759 10308 6763 10364
rect 6763 10308 6819 10364
rect 6819 10308 6823 10364
rect 6759 10304 6823 10308
rect 6839 10364 6903 10368
rect 6839 10308 6843 10364
rect 6843 10308 6899 10364
rect 6899 10308 6903 10364
rect 6839 10304 6903 10308
rect 6919 10364 6983 10368
rect 6919 10308 6923 10364
rect 6923 10308 6979 10364
rect 6979 10308 6983 10364
rect 6919 10304 6983 10308
rect 10497 10364 10561 10368
rect 10497 10308 10501 10364
rect 10501 10308 10557 10364
rect 10557 10308 10561 10364
rect 10497 10304 10561 10308
rect 10577 10364 10641 10368
rect 10577 10308 10581 10364
rect 10581 10308 10637 10364
rect 10637 10308 10641 10364
rect 10577 10304 10641 10308
rect 10657 10364 10721 10368
rect 10657 10308 10661 10364
rect 10661 10308 10717 10364
rect 10717 10308 10721 10364
rect 10657 10304 10721 10308
rect 10737 10364 10801 10368
rect 10737 10308 10741 10364
rect 10741 10308 10797 10364
rect 10797 10308 10801 10364
rect 10737 10304 10801 10308
rect 14315 10364 14379 10368
rect 14315 10308 14319 10364
rect 14319 10308 14375 10364
rect 14375 10308 14379 10364
rect 14315 10304 14379 10308
rect 14395 10364 14459 10368
rect 14395 10308 14399 10364
rect 14399 10308 14455 10364
rect 14455 10308 14459 10364
rect 14395 10304 14459 10308
rect 14475 10364 14539 10368
rect 14475 10308 14479 10364
rect 14479 10308 14535 10364
rect 14535 10308 14539 10364
rect 14475 10304 14539 10308
rect 14555 10364 14619 10368
rect 14555 10308 14559 10364
rect 14559 10308 14615 10364
rect 14615 10308 14619 10364
rect 14555 10304 14619 10308
rect 3521 9820 3585 9824
rect 3521 9764 3525 9820
rect 3525 9764 3581 9820
rect 3581 9764 3585 9820
rect 3521 9760 3585 9764
rect 3601 9820 3665 9824
rect 3601 9764 3605 9820
rect 3605 9764 3661 9820
rect 3661 9764 3665 9820
rect 3601 9760 3665 9764
rect 3681 9820 3745 9824
rect 3681 9764 3685 9820
rect 3685 9764 3741 9820
rect 3741 9764 3745 9820
rect 3681 9760 3745 9764
rect 3761 9820 3825 9824
rect 3761 9764 3765 9820
rect 3765 9764 3821 9820
rect 3821 9764 3825 9820
rect 3761 9760 3825 9764
rect 7339 9820 7403 9824
rect 7339 9764 7343 9820
rect 7343 9764 7399 9820
rect 7399 9764 7403 9820
rect 7339 9760 7403 9764
rect 7419 9820 7483 9824
rect 7419 9764 7423 9820
rect 7423 9764 7479 9820
rect 7479 9764 7483 9820
rect 7419 9760 7483 9764
rect 7499 9820 7563 9824
rect 7499 9764 7503 9820
rect 7503 9764 7559 9820
rect 7559 9764 7563 9820
rect 7499 9760 7563 9764
rect 7579 9820 7643 9824
rect 7579 9764 7583 9820
rect 7583 9764 7639 9820
rect 7639 9764 7643 9820
rect 7579 9760 7643 9764
rect 11157 9820 11221 9824
rect 11157 9764 11161 9820
rect 11161 9764 11217 9820
rect 11217 9764 11221 9820
rect 11157 9760 11221 9764
rect 11237 9820 11301 9824
rect 11237 9764 11241 9820
rect 11241 9764 11297 9820
rect 11297 9764 11301 9820
rect 11237 9760 11301 9764
rect 11317 9820 11381 9824
rect 11317 9764 11321 9820
rect 11321 9764 11377 9820
rect 11377 9764 11381 9820
rect 11317 9760 11381 9764
rect 11397 9820 11461 9824
rect 11397 9764 11401 9820
rect 11401 9764 11457 9820
rect 11457 9764 11461 9820
rect 11397 9760 11461 9764
rect 14975 9820 15039 9824
rect 14975 9764 14979 9820
rect 14979 9764 15035 9820
rect 15035 9764 15039 9820
rect 14975 9760 15039 9764
rect 15055 9820 15119 9824
rect 15055 9764 15059 9820
rect 15059 9764 15115 9820
rect 15115 9764 15119 9820
rect 15055 9760 15119 9764
rect 15135 9820 15199 9824
rect 15135 9764 15139 9820
rect 15139 9764 15195 9820
rect 15195 9764 15199 9820
rect 15135 9760 15199 9764
rect 15215 9820 15279 9824
rect 15215 9764 15219 9820
rect 15219 9764 15275 9820
rect 15275 9764 15279 9820
rect 15215 9760 15279 9764
rect 2861 9276 2925 9280
rect 2861 9220 2865 9276
rect 2865 9220 2921 9276
rect 2921 9220 2925 9276
rect 2861 9216 2925 9220
rect 2941 9276 3005 9280
rect 2941 9220 2945 9276
rect 2945 9220 3001 9276
rect 3001 9220 3005 9276
rect 2941 9216 3005 9220
rect 3021 9276 3085 9280
rect 3021 9220 3025 9276
rect 3025 9220 3081 9276
rect 3081 9220 3085 9276
rect 3021 9216 3085 9220
rect 3101 9276 3165 9280
rect 3101 9220 3105 9276
rect 3105 9220 3161 9276
rect 3161 9220 3165 9276
rect 3101 9216 3165 9220
rect 6679 9276 6743 9280
rect 6679 9220 6683 9276
rect 6683 9220 6739 9276
rect 6739 9220 6743 9276
rect 6679 9216 6743 9220
rect 6759 9276 6823 9280
rect 6759 9220 6763 9276
rect 6763 9220 6819 9276
rect 6819 9220 6823 9276
rect 6759 9216 6823 9220
rect 6839 9276 6903 9280
rect 6839 9220 6843 9276
rect 6843 9220 6899 9276
rect 6899 9220 6903 9276
rect 6839 9216 6903 9220
rect 6919 9276 6983 9280
rect 6919 9220 6923 9276
rect 6923 9220 6979 9276
rect 6979 9220 6983 9276
rect 6919 9216 6983 9220
rect 10497 9276 10561 9280
rect 10497 9220 10501 9276
rect 10501 9220 10557 9276
rect 10557 9220 10561 9276
rect 10497 9216 10561 9220
rect 10577 9276 10641 9280
rect 10577 9220 10581 9276
rect 10581 9220 10637 9276
rect 10637 9220 10641 9276
rect 10577 9216 10641 9220
rect 10657 9276 10721 9280
rect 10657 9220 10661 9276
rect 10661 9220 10717 9276
rect 10717 9220 10721 9276
rect 10657 9216 10721 9220
rect 10737 9276 10801 9280
rect 10737 9220 10741 9276
rect 10741 9220 10797 9276
rect 10797 9220 10801 9276
rect 10737 9216 10801 9220
rect 14315 9276 14379 9280
rect 14315 9220 14319 9276
rect 14319 9220 14375 9276
rect 14375 9220 14379 9276
rect 14315 9216 14379 9220
rect 14395 9276 14459 9280
rect 14395 9220 14399 9276
rect 14399 9220 14455 9276
rect 14455 9220 14459 9276
rect 14395 9216 14459 9220
rect 14475 9276 14539 9280
rect 14475 9220 14479 9276
rect 14479 9220 14535 9276
rect 14535 9220 14539 9276
rect 14475 9216 14539 9220
rect 14555 9276 14619 9280
rect 14555 9220 14559 9276
rect 14559 9220 14615 9276
rect 14615 9220 14619 9276
rect 14555 9216 14619 9220
rect 3521 8732 3585 8736
rect 3521 8676 3525 8732
rect 3525 8676 3581 8732
rect 3581 8676 3585 8732
rect 3521 8672 3585 8676
rect 3601 8732 3665 8736
rect 3601 8676 3605 8732
rect 3605 8676 3661 8732
rect 3661 8676 3665 8732
rect 3601 8672 3665 8676
rect 3681 8732 3745 8736
rect 3681 8676 3685 8732
rect 3685 8676 3741 8732
rect 3741 8676 3745 8732
rect 3681 8672 3745 8676
rect 3761 8732 3825 8736
rect 3761 8676 3765 8732
rect 3765 8676 3821 8732
rect 3821 8676 3825 8732
rect 3761 8672 3825 8676
rect 7339 8732 7403 8736
rect 7339 8676 7343 8732
rect 7343 8676 7399 8732
rect 7399 8676 7403 8732
rect 7339 8672 7403 8676
rect 7419 8732 7483 8736
rect 7419 8676 7423 8732
rect 7423 8676 7479 8732
rect 7479 8676 7483 8732
rect 7419 8672 7483 8676
rect 7499 8732 7563 8736
rect 7499 8676 7503 8732
rect 7503 8676 7559 8732
rect 7559 8676 7563 8732
rect 7499 8672 7563 8676
rect 7579 8732 7643 8736
rect 7579 8676 7583 8732
rect 7583 8676 7639 8732
rect 7639 8676 7643 8732
rect 7579 8672 7643 8676
rect 11157 8732 11221 8736
rect 11157 8676 11161 8732
rect 11161 8676 11217 8732
rect 11217 8676 11221 8732
rect 11157 8672 11221 8676
rect 11237 8732 11301 8736
rect 11237 8676 11241 8732
rect 11241 8676 11297 8732
rect 11297 8676 11301 8732
rect 11237 8672 11301 8676
rect 11317 8732 11381 8736
rect 11317 8676 11321 8732
rect 11321 8676 11377 8732
rect 11377 8676 11381 8732
rect 11317 8672 11381 8676
rect 11397 8732 11461 8736
rect 11397 8676 11401 8732
rect 11401 8676 11457 8732
rect 11457 8676 11461 8732
rect 11397 8672 11461 8676
rect 14975 8732 15039 8736
rect 14975 8676 14979 8732
rect 14979 8676 15035 8732
rect 15035 8676 15039 8732
rect 14975 8672 15039 8676
rect 15055 8732 15119 8736
rect 15055 8676 15059 8732
rect 15059 8676 15115 8732
rect 15115 8676 15119 8732
rect 15055 8672 15119 8676
rect 15135 8732 15199 8736
rect 15135 8676 15139 8732
rect 15139 8676 15195 8732
rect 15195 8676 15199 8732
rect 15135 8672 15199 8676
rect 15215 8732 15279 8736
rect 15215 8676 15219 8732
rect 15219 8676 15275 8732
rect 15275 8676 15279 8732
rect 15215 8672 15279 8676
rect 2861 8188 2925 8192
rect 2861 8132 2865 8188
rect 2865 8132 2921 8188
rect 2921 8132 2925 8188
rect 2861 8128 2925 8132
rect 2941 8188 3005 8192
rect 2941 8132 2945 8188
rect 2945 8132 3001 8188
rect 3001 8132 3005 8188
rect 2941 8128 3005 8132
rect 3021 8188 3085 8192
rect 3021 8132 3025 8188
rect 3025 8132 3081 8188
rect 3081 8132 3085 8188
rect 3021 8128 3085 8132
rect 3101 8188 3165 8192
rect 3101 8132 3105 8188
rect 3105 8132 3161 8188
rect 3161 8132 3165 8188
rect 3101 8128 3165 8132
rect 6679 8188 6743 8192
rect 6679 8132 6683 8188
rect 6683 8132 6739 8188
rect 6739 8132 6743 8188
rect 6679 8128 6743 8132
rect 6759 8188 6823 8192
rect 6759 8132 6763 8188
rect 6763 8132 6819 8188
rect 6819 8132 6823 8188
rect 6759 8128 6823 8132
rect 6839 8188 6903 8192
rect 6839 8132 6843 8188
rect 6843 8132 6899 8188
rect 6899 8132 6903 8188
rect 6839 8128 6903 8132
rect 6919 8188 6983 8192
rect 6919 8132 6923 8188
rect 6923 8132 6979 8188
rect 6979 8132 6983 8188
rect 6919 8128 6983 8132
rect 10497 8188 10561 8192
rect 10497 8132 10501 8188
rect 10501 8132 10557 8188
rect 10557 8132 10561 8188
rect 10497 8128 10561 8132
rect 10577 8188 10641 8192
rect 10577 8132 10581 8188
rect 10581 8132 10637 8188
rect 10637 8132 10641 8188
rect 10577 8128 10641 8132
rect 10657 8188 10721 8192
rect 10657 8132 10661 8188
rect 10661 8132 10717 8188
rect 10717 8132 10721 8188
rect 10657 8128 10721 8132
rect 10737 8188 10801 8192
rect 10737 8132 10741 8188
rect 10741 8132 10797 8188
rect 10797 8132 10801 8188
rect 10737 8128 10801 8132
rect 14315 8188 14379 8192
rect 14315 8132 14319 8188
rect 14319 8132 14375 8188
rect 14375 8132 14379 8188
rect 14315 8128 14379 8132
rect 14395 8188 14459 8192
rect 14395 8132 14399 8188
rect 14399 8132 14455 8188
rect 14455 8132 14459 8188
rect 14395 8128 14459 8132
rect 14475 8188 14539 8192
rect 14475 8132 14479 8188
rect 14479 8132 14535 8188
rect 14535 8132 14539 8188
rect 14475 8128 14539 8132
rect 14555 8188 14619 8192
rect 14555 8132 14559 8188
rect 14559 8132 14615 8188
rect 14615 8132 14619 8188
rect 14555 8128 14619 8132
rect 3521 7644 3585 7648
rect 3521 7588 3525 7644
rect 3525 7588 3581 7644
rect 3581 7588 3585 7644
rect 3521 7584 3585 7588
rect 3601 7644 3665 7648
rect 3601 7588 3605 7644
rect 3605 7588 3661 7644
rect 3661 7588 3665 7644
rect 3601 7584 3665 7588
rect 3681 7644 3745 7648
rect 3681 7588 3685 7644
rect 3685 7588 3741 7644
rect 3741 7588 3745 7644
rect 3681 7584 3745 7588
rect 3761 7644 3825 7648
rect 3761 7588 3765 7644
rect 3765 7588 3821 7644
rect 3821 7588 3825 7644
rect 3761 7584 3825 7588
rect 7339 7644 7403 7648
rect 7339 7588 7343 7644
rect 7343 7588 7399 7644
rect 7399 7588 7403 7644
rect 7339 7584 7403 7588
rect 7419 7644 7483 7648
rect 7419 7588 7423 7644
rect 7423 7588 7479 7644
rect 7479 7588 7483 7644
rect 7419 7584 7483 7588
rect 7499 7644 7563 7648
rect 7499 7588 7503 7644
rect 7503 7588 7559 7644
rect 7559 7588 7563 7644
rect 7499 7584 7563 7588
rect 7579 7644 7643 7648
rect 7579 7588 7583 7644
rect 7583 7588 7639 7644
rect 7639 7588 7643 7644
rect 7579 7584 7643 7588
rect 11157 7644 11221 7648
rect 11157 7588 11161 7644
rect 11161 7588 11217 7644
rect 11217 7588 11221 7644
rect 11157 7584 11221 7588
rect 11237 7644 11301 7648
rect 11237 7588 11241 7644
rect 11241 7588 11297 7644
rect 11297 7588 11301 7644
rect 11237 7584 11301 7588
rect 11317 7644 11381 7648
rect 11317 7588 11321 7644
rect 11321 7588 11377 7644
rect 11377 7588 11381 7644
rect 11317 7584 11381 7588
rect 11397 7644 11461 7648
rect 11397 7588 11401 7644
rect 11401 7588 11457 7644
rect 11457 7588 11461 7644
rect 11397 7584 11461 7588
rect 14975 7644 15039 7648
rect 14975 7588 14979 7644
rect 14979 7588 15035 7644
rect 15035 7588 15039 7644
rect 14975 7584 15039 7588
rect 15055 7644 15119 7648
rect 15055 7588 15059 7644
rect 15059 7588 15115 7644
rect 15115 7588 15119 7644
rect 15055 7584 15119 7588
rect 15135 7644 15199 7648
rect 15135 7588 15139 7644
rect 15139 7588 15195 7644
rect 15195 7588 15199 7644
rect 15135 7584 15199 7588
rect 15215 7644 15279 7648
rect 15215 7588 15219 7644
rect 15219 7588 15275 7644
rect 15275 7588 15279 7644
rect 15215 7584 15279 7588
rect 2861 7100 2925 7104
rect 2861 7044 2865 7100
rect 2865 7044 2921 7100
rect 2921 7044 2925 7100
rect 2861 7040 2925 7044
rect 2941 7100 3005 7104
rect 2941 7044 2945 7100
rect 2945 7044 3001 7100
rect 3001 7044 3005 7100
rect 2941 7040 3005 7044
rect 3021 7100 3085 7104
rect 3021 7044 3025 7100
rect 3025 7044 3081 7100
rect 3081 7044 3085 7100
rect 3021 7040 3085 7044
rect 3101 7100 3165 7104
rect 3101 7044 3105 7100
rect 3105 7044 3161 7100
rect 3161 7044 3165 7100
rect 3101 7040 3165 7044
rect 6679 7100 6743 7104
rect 6679 7044 6683 7100
rect 6683 7044 6739 7100
rect 6739 7044 6743 7100
rect 6679 7040 6743 7044
rect 6759 7100 6823 7104
rect 6759 7044 6763 7100
rect 6763 7044 6819 7100
rect 6819 7044 6823 7100
rect 6759 7040 6823 7044
rect 6839 7100 6903 7104
rect 6839 7044 6843 7100
rect 6843 7044 6899 7100
rect 6899 7044 6903 7100
rect 6839 7040 6903 7044
rect 6919 7100 6983 7104
rect 6919 7044 6923 7100
rect 6923 7044 6979 7100
rect 6979 7044 6983 7100
rect 6919 7040 6983 7044
rect 10497 7100 10561 7104
rect 10497 7044 10501 7100
rect 10501 7044 10557 7100
rect 10557 7044 10561 7100
rect 10497 7040 10561 7044
rect 10577 7100 10641 7104
rect 10577 7044 10581 7100
rect 10581 7044 10637 7100
rect 10637 7044 10641 7100
rect 10577 7040 10641 7044
rect 10657 7100 10721 7104
rect 10657 7044 10661 7100
rect 10661 7044 10717 7100
rect 10717 7044 10721 7100
rect 10657 7040 10721 7044
rect 10737 7100 10801 7104
rect 10737 7044 10741 7100
rect 10741 7044 10797 7100
rect 10797 7044 10801 7100
rect 10737 7040 10801 7044
rect 14315 7100 14379 7104
rect 14315 7044 14319 7100
rect 14319 7044 14375 7100
rect 14375 7044 14379 7100
rect 14315 7040 14379 7044
rect 14395 7100 14459 7104
rect 14395 7044 14399 7100
rect 14399 7044 14455 7100
rect 14455 7044 14459 7100
rect 14395 7040 14459 7044
rect 14475 7100 14539 7104
rect 14475 7044 14479 7100
rect 14479 7044 14535 7100
rect 14535 7044 14539 7100
rect 14475 7040 14539 7044
rect 14555 7100 14619 7104
rect 14555 7044 14559 7100
rect 14559 7044 14615 7100
rect 14615 7044 14619 7100
rect 14555 7040 14619 7044
rect 3521 6556 3585 6560
rect 3521 6500 3525 6556
rect 3525 6500 3581 6556
rect 3581 6500 3585 6556
rect 3521 6496 3585 6500
rect 3601 6556 3665 6560
rect 3601 6500 3605 6556
rect 3605 6500 3661 6556
rect 3661 6500 3665 6556
rect 3601 6496 3665 6500
rect 3681 6556 3745 6560
rect 3681 6500 3685 6556
rect 3685 6500 3741 6556
rect 3741 6500 3745 6556
rect 3681 6496 3745 6500
rect 3761 6556 3825 6560
rect 3761 6500 3765 6556
rect 3765 6500 3821 6556
rect 3821 6500 3825 6556
rect 3761 6496 3825 6500
rect 7339 6556 7403 6560
rect 7339 6500 7343 6556
rect 7343 6500 7399 6556
rect 7399 6500 7403 6556
rect 7339 6496 7403 6500
rect 7419 6556 7483 6560
rect 7419 6500 7423 6556
rect 7423 6500 7479 6556
rect 7479 6500 7483 6556
rect 7419 6496 7483 6500
rect 7499 6556 7563 6560
rect 7499 6500 7503 6556
rect 7503 6500 7559 6556
rect 7559 6500 7563 6556
rect 7499 6496 7563 6500
rect 7579 6556 7643 6560
rect 7579 6500 7583 6556
rect 7583 6500 7639 6556
rect 7639 6500 7643 6556
rect 7579 6496 7643 6500
rect 11157 6556 11221 6560
rect 11157 6500 11161 6556
rect 11161 6500 11217 6556
rect 11217 6500 11221 6556
rect 11157 6496 11221 6500
rect 11237 6556 11301 6560
rect 11237 6500 11241 6556
rect 11241 6500 11297 6556
rect 11297 6500 11301 6556
rect 11237 6496 11301 6500
rect 11317 6556 11381 6560
rect 11317 6500 11321 6556
rect 11321 6500 11377 6556
rect 11377 6500 11381 6556
rect 11317 6496 11381 6500
rect 11397 6556 11461 6560
rect 11397 6500 11401 6556
rect 11401 6500 11457 6556
rect 11457 6500 11461 6556
rect 11397 6496 11461 6500
rect 14975 6556 15039 6560
rect 14975 6500 14979 6556
rect 14979 6500 15035 6556
rect 15035 6500 15039 6556
rect 14975 6496 15039 6500
rect 15055 6556 15119 6560
rect 15055 6500 15059 6556
rect 15059 6500 15115 6556
rect 15115 6500 15119 6556
rect 15055 6496 15119 6500
rect 15135 6556 15199 6560
rect 15135 6500 15139 6556
rect 15139 6500 15195 6556
rect 15195 6500 15199 6556
rect 15135 6496 15199 6500
rect 15215 6556 15279 6560
rect 15215 6500 15219 6556
rect 15219 6500 15275 6556
rect 15275 6500 15279 6556
rect 15215 6496 15279 6500
rect 2861 6012 2925 6016
rect 2861 5956 2865 6012
rect 2865 5956 2921 6012
rect 2921 5956 2925 6012
rect 2861 5952 2925 5956
rect 2941 6012 3005 6016
rect 2941 5956 2945 6012
rect 2945 5956 3001 6012
rect 3001 5956 3005 6012
rect 2941 5952 3005 5956
rect 3021 6012 3085 6016
rect 3021 5956 3025 6012
rect 3025 5956 3081 6012
rect 3081 5956 3085 6012
rect 3021 5952 3085 5956
rect 3101 6012 3165 6016
rect 3101 5956 3105 6012
rect 3105 5956 3161 6012
rect 3161 5956 3165 6012
rect 3101 5952 3165 5956
rect 6679 6012 6743 6016
rect 6679 5956 6683 6012
rect 6683 5956 6739 6012
rect 6739 5956 6743 6012
rect 6679 5952 6743 5956
rect 6759 6012 6823 6016
rect 6759 5956 6763 6012
rect 6763 5956 6819 6012
rect 6819 5956 6823 6012
rect 6759 5952 6823 5956
rect 6839 6012 6903 6016
rect 6839 5956 6843 6012
rect 6843 5956 6899 6012
rect 6899 5956 6903 6012
rect 6839 5952 6903 5956
rect 6919 6012 6983 6016
rect 6919 5956 6923 6012
rect 6923 5956 6979 6012
rect 6979 5956 6983 6012
rect 6919 5952 6983 5956
rect 10497 6012 10561 6016
rect 10497 5956 10501 6012
rect 10501 5956 10557 6012
rect 10557 5956 10561 6012
rect 10497 5952 10561 5956
rect 10577 6012 10641 6016
rect 10577 5956 10581 6012
rect 10581 5956 10637 6012
rect 10637 5956 10641 6012
rect 10577 5952 10641 5956
rect 10657 6012 10721 6016
rect 10657 5956 10661 6012
rect 10661 5956 10717 6012
rect 10717 5956 10721 6012
rect 10657 5952 10721 5956
rect 10737 6012 10801 6016
rect 10737 5956 10741 6012
rect 10741 5956 10797 6012
rect 10797 5956 10801 6012
rect 10737 5952 10801 5956
rect 14315 6012 14379 6016
rect 14315 5956 14319 6012
rect 14319 5956 14375 6012
rect 14375 5956 14379 6012
rect 14315 5952 14379 5956
rect 14395 6012 14459 6016
rect 14395 5956 14399 6012
rect 14399 5956 14455 6012
rect 14455 5956 14459 6012
rect 14395 5952 14459 5956
rect 14475 6012 14539 6016
rect 14475 5956 14479 6012
rect 14479 5956 14535 6012
rect 14535 5956 14539 6012
rect 14475 5952 14539 5956
rect 14555 6012 14619 6016
rect 14555 5956 14559 6012
rect 14559 5956 14615 6012
rect 14615 5956 14619 6012
rect 14555 5952 14619 5956
rect 3521 5468 3585 5472
rect 3521 5412 3525 5468
rect 3525 5412 3581 5468
rect 3581 5412 3585 5468
rect 3521 5408 3585 5412
rect 3601 5468 3665 5472
rect 3601 5412 3605 5468
rect 3605 5412 3661 5468
rect 3661 5412 3665 5468
rect 3601 5408 3665 5412
rect 3681 5468 3745 5472
rect 3681 5412 3685 5468
rect 3685 5412 3741 5468
rect 3741 5412 3745 5468
rect 3681 5408 3745 5412
rect 3761 5468 3825 5472
rect 3761 5412 3765 5468
rect 3765 5412 3821 5468
rect 3821 5412 3825 5468
rect 3761 5408 3825 5412
rect 7339 5468 7403 5472
rect 7339 5412 7343 5468
rect 7343 5412 7399 5468
rect 7399 5412 7403 5468
rect 7339 5408 7403 5412
rect 7419 5468 7483 5472
rect 7419 5412 7423 5468
rect 7423 5412 7479 5468
rect 7479 5412 7483 5468
rect 7419 5408 7483 5412
rect 7499 5468 7563 5472
rect 7499 5412 7503 5468
rect 7503 5412 7559 5468
rect 7559 5412 7563 5468
rect 7499 5408 7563 5412
rect 7579 5468 7643 5472
rect 7579 5412 7583 5468
rect 7583 5412 7639 5468
rect 7639 5412 7643 5468
rect 7579 5408 7643 5412
rect 11157 5468 11221 5472
rect 11157 5412 11161 5468
rect 11161 5412 11217 5468
rect 11217 5412 11221 5468
rect 11157 5408 11221 5412
rect 11237 5468 11301 5472
rect 11237 5412 11241 5468
rect 11241 5412 11297 5468
rect 11297 5412 11301 5468
rect 11237 5408 11301 5412
rect 11317 5468 11381 5472
rect 11317 5412 11321 5468
rect 11321 5412 11377 5468
rect 11377 5412 11381 5468
rect 11317 5408 11381 5412
rect 11397 5468 11461 5472
rect 11397 5412 11401 5468
rect 11401 5412 11457 5468
rect 11457 5412 11461 5468
rect 11397 5408 11461 5412
rect 14975 5468 15039 5472
rect 14975 5412 14979 5468
rect 14979 5412 15035 5468
rect 15035 5412 15039 5468
rect 14975 5408 15039 5412
rect 15055 5468 15119 5472
rect 15055 5412 15059 5468
rect 15059 5412 15115 5468
rect 15115 5412 15119 5468
rect 15055 5408 15119 5412
rect 15135 5468 15199 5472
rect 15135 5412 15139 5468
rect 15139 5412 15195 5468
rect 15195 5412 15199 5468
rect 15135 5408 15199 5412
rect 15215 5468 15279 5472
rect 15215 5412 15219 5468
rect 15219 5412 15275 5468
rect 15275 5412 15279 5468
rect 15215 5408 15279 5412
rect 2861 4924 2925 4928
rect 2861 4868 2865 4924
rect 2865 4868 2921 4924
rect 2921 4868 2925 4924
rect 2861 4864 2925 4868
rect 2941 4924 3005 4928
rect 2941 4868 2945 4924
rect 2945 4868 3001 4924
rect 3001 4868 3005 4924
rect 2941 4864 3005 4868
rect 3021 4924 3085 4928
rect 3021 4868 3025 4924
rect 3025 4868 3081 4924
rect 3081 4868 3085 4924
rect 3021 4864 3085 4868
rect 3101 4924 3165 4928
rect 3101 4868 3105 4924
rect 3105 4868 3161 4924
rect 3161 4868 3165 4924
rect 3101 4864 3165 4868
rect 6679 4924 6743 4928
rect 6679 4868 6683 4924
rect 6683 4868 6739 4924
rect 6739 4868 6743 4924
rect 6679 4864 6743 4868
rect 6759 4924 6823 4928
rect 6759 4868 6763 4924
rect 6763 4868 6819 4924
rect 6819 4868 6823 4924
rect 6759 4864 6823 4868
rect 6839 4924 6903 4928
rect 6839 4868 6843 4924
rect 6843 4868 6899 4924
rect 6899 4868 6903 4924
rect 6839 4864 6903 4868
rect 6919 4924 6983 4928
rect 6919 4868 6923 4924
rect 6923 4868 6979 4924
rect 6979 4868 6983 4924
rect 6919 4864 6983 4868
rect 10497 4924 10561 4928
rect 10497 4868 10501 4924
rect 10501 4868 10557 4924
rect 10557 4868 10561 4924
rect 10497 4864 10561 4868
rect 10577 4924 10641 4928
rect 10577 4868 10581 4924
rect 10581 4868 10637 4924
rect 10637 4868 10641 4924
rect 10577 4864 10641 4868
rect 10657 4924 10721 4928
rect 10657 4868 10661 4924
rect 10661 4868 10717 4924
rect 10717 4868 10721 4924
rect 10657 4864 10721 4868
rect 10737 4924 10801 4928
rect 10737 4868 10741 4924
rect 10741 4868 10797 4924
rect 10797 4868 10801 4924
rect 10737 4864 10801 4868
rect 14315 4924 14379 4928
rect 14315 4868 14319 4924
rect 14319 4868 14375 4924
rect 14375 4868 14379 4924
rect 14315 4864 14379 4868
rect 14395 4924 14459 4928
rect 14395 4868 14399 4924
rect 14399 4868 14455 4924
rect 14455 4868 14459 4924
rect 14395 4864 14459 4868
rect 14475 4924 14539 4928
rect 14475 4868 14479 4924
rect 14479 4868 14535 4924
rect 14535 4868 14539 4924
rect 14475 4864 14539 4868
rect 14555 4924 14619 4928
rect 14555 4868 14559 4924
rect 14559 4868 14615 4924
rect 14615 4868 14619 4924
rect 14555 4864 14619 4868
rect 3521 4380 3585 4384
rect 3521 4324 3525 4380
rect 3525 4324 3581 4380
rect 3581 4324 3585 4380
rect 3521 4320 3585 4324
rect 3601 4380 3665 4384
rect 3601 4324 3605 4380
rect 3605 4324 3661 4380
rect 3661 4324 3665 4380
rect 3601 4320 3665 4324
rect 3681 4380 3745 4384
rect 3681 4324 3685 4380
rect 3685 4324 3741 4380
rect 3741 4324 3745 4380
rect 3681 4320 3745 4324
rect 3761 4380 3825 4384
rect 3761 4324 3765 4380
rect 3765 4324 3821 4380
rect 3821 4324 3825 4380
rect 3761 4320 3825 4324
rect 7339 4380 7403 4384
rect 7339 4324 7343 4380
rect 7343 4324 7399 4380
rect 7399 4324 7403 4380
rect 7339 4320 7403 4324
rect 7419 4380 7483 4384
rect 7419 4324 7423 4380
rect 7423 4324 7479 4380
rect 7479 4324 7483 4380
rect 7419 4320 7483 4324
rect 7499 4380 7563 4384
rect 7499 4324 7503 4380
rect 7503 4324 7559 4380
rect 7559 4324 7563 4380
rect 7499 4320 7563 4324
rect 7579 4380 7643 4384
rect 7579 4324 7583 4380
rect 7583 4324 7639 4380
rect 7639 4324 7643 4380
rect 7579 4320 7643 4324
rect 11157 4380 11221 4384
rect 11157 4324 11161 4380
rect 11161 4324 11217 4380
rect 11217 4324 11221 4380
rect 11157 4320 11221 4324
rect 11237 4380 11301 4384
rect 11237 4324 11241 4380
rect 11241 4324 11297 4380
rect 11297 4324 11301 4380
rect 11237 4320 11301 4324
rect 11317 4380 11381 4384
rect 11317 4324 11321 4380
rect 11321 4324 11377 4380
rect 11377 4324 11381 4380
rect 11317 4320 11381 4324
rect 11397 4380 11461 4384
rect 11397 4324 11401 4380
rect 11401 4324 11457 4380
rect 11457 4324 11461 4380
rect 11397 4320 11461 4324
rect 14975 4380 15039 4384
rect 14975 4324 14979 4380
rect 14979 4324 15035 4380
rect 15035 4324 15039 4380
rect 14975 4320 15039 4324
rect 15055 4380 15119 4384
rect 15055 4324 15059 4380
rect 15059 4324 15115 4380
rect 15115 4324 15119 4380
rect 15055 4320 15119 4324
rect 15135 4380 15199 4384
rect 15135 4324 15139 4380
rect 15139 4324 15195 4380
rect 15195 4324 15199 4380
rect 15135 4320 15199 4324
rect 15215 4380 15279 4384
rect 15215 4324 15219 4380
rect 15219 4324 15275 4380
rect 15275 4324 15279 4380
rect 15215 4320 15279 4324
rect 2861 3836 2925 3840
rect 2861 3780 2865 3836
rect 2865 3780 2921 3836
rect 2921 3780 2925 3836
rect 2861 3776 2925 3780
rect 2941 3836 3005 3840
rect 2941 3780 2945 3836
rect 2945 3780 3001 3836
rect 3001 3780 3005 3836
rect 2941 3776 3005 3780
rect 3021 3836 3085 3840
rect 3021 3780 3025 3836
rect 3025 3780 3081 3836
rect 3081 3780 3085 3836
rect 3021 3776 3085 3780
rect 3101 3836 3165 3840
rect 3101 3780 3105 3836
rect 3105 3780 3161 3836
rect 3161 3780 3165 3836
rect 3101 3776 3165 3780
rect 6679 3836 6743 3840
rect 6679 3780 6683 3836
rect 6683 3780 6739 3836
rect 6739 3780 6743 3836
rect 6679 3776 6743 3780
rect 6759 3836 6823 3840
rect 6759 3780 6763 3836
rect 6763 3780 6819 3836
rect 6819 3780 6823 3836
rect 6759 3776 6823 3780
rect 6839 3836 6903 3840
rect 6839 3780 6843 3836
rect 6843 3780 6899 3836
rect 6899 3780 6903 3836
rect 6839 3776 6903 3780
rect 6919 3836 6983 3840
rect 6919 3780 6923 3836
rect 6923 3780 6979 3836
rect 6979 3780 6983 3836
rect 6919 3776 6983 3780
rect 10497 3836 10561 3840
rect 10497 3780 10501 3836
rect 10501 3780 10557 3836
rect 10557 3780 10561 3836
rect 10497 3776 10561 3780
rect 10577 3836 10641 3840
rect 10577 3780 10581 3836
rect 10581 3780 10637 3836
rect 10637 3780 10641 3836
rect 10577 3776 10641 3780
rect 10657 3836 10721 3840
rect 10657 3780 10661 3836
rect 10661 3780 10717 3836
rect 10717 3780 10721 3836
rect 10657 3776 10721 3780
rect 10737 3836 10801 3840
rect 10737 3780 10741 3836
rect 10741 3780 10797 3836
rect 10797 3780 10801 3836
rect 10737 3776 10801 3780
rect 14315 3836 14379 3840
rect 14315 3780 14319 3836
rect 14319 3780 14375 3836
rect 14375 3780 14379 3836
rect 14315 3776 14379 3780
rect 14395 3836 14459 3840
rect 14395 3780 14399 3836
rect 14399 3780 14455 3836
rect 14455 3780 14459 3836
rect 14395 3776 14459 3780
rect 14475 3836 14539 3840
rect 14475 3780 14479 3836
rect 14479 3780 14535 3836
rect 14535 3780 14539 3836
rect 14475 3776 14539 3780
rect 14555 3836 14619 3840
rect 14555 3780 14559 3836
rect 14559 3780 14615 3836
rect 14615 3780 14619 3836
rect 14555 3776 14619 3780
rect 3521 3292 3585 3296
rect 3521 3236 3525 3292
rect 3525 3236 3581 3292
rect 3581 3236 3585 3292
rect 3521 3232 3585 3236
rect 3601 3292 3665 3296
rect 3601 3236 3605 3292
rect 3605 3236 3661 3292
rect 3661 3236 3665 3292
rect 3601 3232 3665 3236
rect 3681 3292 3745 3296
rect 3681 3236 3685 3292
rect 3685 3236 3741 3292
rect 3741 3236 3745 3292
rect 3681 3232 3745 3236
rect 3761 3292 3825 3296
rect 3761 3236 3765 3292
rect 3765 3236 3821 3292
rect 3821 3236 3825 3292
rect 3761 3232 3825 3236
rect 7339 3292 7403 3296
rect 7339 3236 7343 3292
rect 7343 3236 7399 3292
rect 7399 3236 7403 3292
rect 7339 3232 7403 3236
rect 7419 3292 7483 3296
rect 7419 3236 7423 3292
rect 7423 3236 7479 3292
rect 7479 3236 7483 3292
rect 7419 3232 7483 3236
rect 7499 3292 7563 3296
rect 7499 3236 7503 3292
rect 7503 3236 7559 3292
rect 7559 3236 7563 3292
rect 7499 3232 7563 3236
rect 7579 3292 7643 3296
rect 7579 3236 7583 3292
rect 7583 3236 7639 3292
rect 7639 3236 7643 3292
rect 7579 3232 7643 3236
rect 11157 3292 11221 3296
rect 11157 3236 11161 3292
rect 11161 3236 11217 3292
rect 11217 3236 11221 3292
rect 11157 3232 11221 3236
rect 11237 3292 11301 3296
rect 11237 3236 11241 3292
rect 11241 3236 11297 3292
rect 11297 3236 11301 3292
rect 11237 3232 11301 3236
rect 11317 3292 11381 3296
rect 11317 3236 11321 3292
rect 11321 3236 11377 3292
rect 11377 3236 11381 3292
rect 11317 3232 11381 3236
rect 11397 3292 11461 3296
rect 11397 3236 11401 3292
rect 11401 3236 11457 3292
rect 11457 3236 11461 3292
rect 11397 3232 11461 3236
rect 14975 3292 15039 3296
rect 14975 3236 14979 3292
rect 14979 3236 15035 3292
rect 15035 3236 15039 3292
rect 14975 3232 15039 3236
rect 15055 3292 15119 3296
rect 15055 3236 15059 3292
rect 15059 3236 15115 3292
rect 15115 3236 15119 3292
rect 15055 3232 15119 3236
rect 15135 3292 15199 3296
rect 15135 3236 15139 3292
rect 15139 3236 15195 3292
rect 15195 3236 15199 3292
rect 15135 3232 15199 3236
rect 15215 3292 15279 3296
rect 15215 3236 15219 3292
rect 15219 3236 15275 3292
rect 15275 3236 15279 3292
rect 15215 3232 15279 3236
rect 2861 2748 2925 2752
rect 2861 2692 2865 2748
rect 2865 2692 2921 2748
rect 2921 2692 2925 2748
rect 2861 2688 2925 2692
rect 2941 2748 3005 2752
rect 2941 2692 2945 2748
rect 2945 2692 3001 2748
rect 3001 2692 3005 2748
rect 2941 2688 3005 2692
rect 3021 2748 3085 2752
rect 3021 2692 3025 2748
rect 3025 2692 3081 2748
rect 3081 2692 3085 2748
rect 3021 2688 3085 2692
rect 3101 2748 3165 2752
rect 3101 2692 3105 2748
rect 3105 2692 3161 2748
rect 3161 2692 3165 2748
rect 3101 2688 3165 2692
rect 6679 2748 6743 2752
rect 6679 2692 6683 2748
rect 6683 2692 6739 2748
rect 6739 2692 6743 2748
rect 6679 2688 6743 2692
rect 6759 2748 6823 2752
rect 6759 2692 6763 2748
rect 6763 2692 6819 2748
rect 6819 2692 6823 2748
rect 6759 2688 6823 2692
rect 6839 2748 6903 2752
rect 6839 2692 6843 2748
rect 6843 2692 6899 2748
rect 6899 2692 6903 2748
rect 6839 2688 6903 2692
rect 6919 2748 6983 2752
rect 6919 2692 6923 2748
rect 6923 2692 6979 2748
rect 6979 2692 6983 2748
rect 6919 2688 6983 2692
rect 10497 2748 10561 2752
rect 10497 2692 10501 2748
rect 10501 2692 10557 2748
rect 10557 2692 10561 2748
rect 10497 2688 10561 2692
rect 10577 2748 10641 2752
rect 10577 2692 10581 2748
rect 10581 2692 10637 2748
rect 10637 2692 10641 2748
rect 10577 2688 10641 2692
rect 10657 2748 10721 2752
rect 10657 2692 10661 2748
rect 10661 2692 10717 2748
rect 10717 2692 10721 2748
rect 10657 2688 10721 2692
rect 10737 2748 10801 2752
rect 10737 2692 10741 2748
rect 10741 2692 10797 2748
rect 10797 2692 10801 2748
rect 10737 2688 10801 2692
rect 14315 2748 14379 2752
rect 14315 2692 14319 2748
rect 14319 2692 14375 2748
rect 14375 2692 14379 2748
rect 14315 2688 14379 2692
rect 14395 2748 14459 2752
rect 14395 2692 14399 2748
rect 14399 2692 14455 2748
rect 14455 2692 14459 2748
rect 14395 2688 14459 2692
rect 14475 2748 14539 2752
rect 14475 2692 14479 2748
rect 14479 2692 14535 2748
rect 14535 2692 14539 2748
rect 14475 2688 14539 2692
rect 14555 2748 14619 2752
rect 14555 2692 14559 2748
rect 14559 2692 14615 2748
rect 14615 2692 14619 2748
rect 14555 2688 14619 2692
rect 3521 2204 3585 2208
rect 3521 2148 3525 2204
rect 3525 2148 3581 2204
rect 3581 2148 3585 2204
rect 3521 2144 3585 2148
rect 3601 2204 3665 2208
rect 3601 2148 3605 2204
rect 3605 2148 3661 2204
rect 3661 2148 3665 2204
rect 3601 2144 3665 2148
rect 3681 2204 3745 2208
rect 3681 2148 3685 2204
rect 3685 2148 3741 2204
rect 3741 2148 3745 2204
rect 3681 2144 3745 2148
rect 3761 2204 3825 2208
rect 3761 2148 3765 2204
rect 3765 2148 3821 2204
rect 3821 2148 3825 2204
rect 3761 2144 3825 2148
rect 7339 2204 7403 2208
rect 7339 2148 7343 2204
rect 7343 2148 7399 2204
rect 7399 2148 7403 2204
rect 7339 2144 7403 2148
rect 7419 2204 7483 2208
rect 7419 2148 7423 2204
rect 7423 2148 7479 2204
rect 7479 2148 7483 2204
rect 7419 2144 7483 2148
rect 7499 2204 7563 2208
rect 7499 2148 7503 2204
rect 7503 2148 7559 2204
rect 7559 2148 7563 2204
rect 7499 2144 7563 2148
rect 7579 2204 7643 2208
rect 7579 2148 7583 2204
rect 7583 2148 7639 2204
rect 7639 2148 7643 2204
rect 7579 2144 7643 2148
rect 11157 2204 11221 2208
rect 11157 2148 11161 2204
rect 11161 2148 11217 2204
rect 11217 2148 11221 2204
rect 11157 2144 11221 2148
rect 11237 2204 11301 2208
rect 11237 2148 11241 2204
rect 11241 2148 11297 2204
rect 11297 2148 11301 2204
rect 11237 2144 11301 2148
rect 11317 2204 11381 2208
rect 11317 2148 11321 2204
rect 11321 2148 11377 2204
rect 11377 2148 11381 2204
rect 11317 2144 11381 2148
rect 11397 2204 11461 2208
rect 11397 2148 11401 2204
rect 11401 2148 11457 2204
rect 11457 2148 11461 2204
rect 11397 2144 11461 2148
rect 14975 2204 15039 2208
rect 14975 2148 14979 2204
rect 14979 2148 15035 2204
rect 15035 2148 15039 2204
rect 14975 2144 15039 2148
rect 15055 2204 15119 2208
rect 15055 2148 15059 2204
rect 15059 2148 15115 2204
rect 15115 2148 15119 2204
rect 15055 2144 15119 2148
rect 15135 2204 15199 2208
rect 15135 2148 15139 2204
rect 15139 2148 15195 2204
rect 15195 2148 15199 2204
rect 15135 2144 15199 2148
rect 15215 2204 15279 2208
rect 15215 2148 15219 2204
rect 15219 2148 15275 2204
rect 15275 2148 15279 2204
rect 15215 2144 15279 2148
<< metal4 >>
rect 2853 16896 3173 17456
rect 2853 16832 2861 16896
rect 2925 16832 2941 16896
rect 3005 16832 3021 16896
rect 3085 16832 3101 16896
rect 3165 16832 3173 16896
rect 2853 15808 3173 16832
rect 2853 15744 2861 15808
rect 2925 15744 2941 15808
rect 3005 15744 3021 15808
rect 3085 15744 3101 15808
rect 3165 15744 3173 15808
rect 2853 15622 3173 15744
rect 2853 15386 2895 15622
rect 3131 15386 3173 15622
rect 2853 14720 3173 15386
rect 2853 14656 2861 14720
rect 2925 14656 2941 14720
rect 3005 14656 3021 14720
rect 3085 14656 3101 14720
rect 3165 14656 3173 14720
rect 2853 13632 3173 14656
rect 2853 13568 2861 13632
rect 2925 13568 2941 13632
rect 3005 13568 3021 13632
rect 3085 13568 3101 13632
rect 3165 13568 3173 13632
rect 2853 12544 3173 13568
rect 2853 12480 2861 12544
rect 2925 12480 2941 12544
rect 3005 12480 3021 12544
rect 3085 12480 3101 12544
rect 3165 12480 3173 12544
rect 2853 11814 3173 12480
rect 2853 11578 2895 11814
rect 3131 11578 3173 11814
rect 2853 11456 3173 11578
rect 2853 11392 2861 11456
rect 2925 11392 2941 11456
rect 3005 11392 3021 11456
rect 3085 11392 3101 11456
rect 3165 11392 3173 11456
rect 2853 10368 3173 11392
rect 2853 10304 2861 10368
rect 2925 10304 2941 10368
rect 3005 10304 3021 10368
rect 3085 10304 3101 10368
rect 3165 10304 3173 10368
rect 2853 9280 3173 10304
rect 2853 9216 2861 9280
rect 2925 9216 2941 9280
rect 3005 9216 3021 9280
rect 3085 9216 3101 9280
rect 3165 9216 3173 9280
rect 2853 8192 3173 9216
rect 2853 8128 2861 8192
rect 2925 8128 2941 8192
rect 3005 8128 3021 8192
rect 3085 8128 3101 8192
rect 3165 8128 3173 8192
rect 2853 8006 3173 8128
rect 2853 7770 2895 8006
rect 3131 7770 3173 8006
rect 2853 7104 3173 7770
rect 2853 7040 2861 7104
rect 2925 7040 2941 7104
rect 3005 7040 3021 7104
rect 3085 7040 3101 7104
rect 3165 7040 3173 7104
rect 2853 6016 3173 7040
rect 2853 5952 2861 6016
rect 2925 5952 2941 6016
rect 3005 5952 3021 6016
rect 3085 5952 3101 6016
rect 3165 5952 3173 6016
rect 2853 4928 3173 5952
rect 2853 4864 2861 4928
rect 2925 4864 2941 4928
rect 3005 4864 3021 4928
rect 3085 4864 3101 4928
rect 3165 4864 3173 4928
rect 2853 4198 3173 4864
rect 2853 3962 2895 4198
rect 3131 3962 3173 4198
rect 2853 3840 3173 3962
rect 2853 3776 2861 3840
rect 2925 3776 2941 3840
rect 3005 3776 3021 3840
rect 3085 3776 3101 3840
rect 3165 3776 3173 3840
rect 2853 2752 3173 3776
rect 2853 2688 2861 2752
rect 2925 2688 2941 2752
rect 3005 2688 3021 2752
rect 3085 2688 3101 2752
rect 3165 2688 3173 2752
rect 2853 2128 3173 2688
rect 3513 17440 3833 17456
rect 3513 17376 3521 17440
rect 3585 17376 3601 17440
rect 3665 17376 3681 17440
rect 3745 17376 3761 17440
rect 3825 17376 3833 17440
rect 3513 16352 3833 17376
rect 3513 16288 3521 16352
rect 3585 16288 3601 16352
rect 3665 16288 3681 16352
rect 3745 16288 3761 16352
rect 3825 16288 3833 16352
rect 3513 16282 3833 16288
rect 3513 16046 3555 16282
rect 3791 16046 3833 16282
rect 3513 15264 3833 16046
rect 3513 15200 3521 15264
rect 3585 15200 3601 15264
rect 3665 15200 3681 15264
rect 3745 15200 3761 15264
rect 3825 15200 3833 15264
rect 3513 14176 3833 15200
rect 3513 14112 3521 14176
rect 3585 14112 3601 14176
rect 3665 14112 3681 14176
rect 3745 14112 3761 14176
rect 3825 14112 3833 14176
rect 3513 13088 3833 14112
rect 3513 13024 3521 13088
rect 3585 13024 3601 13088
rect 3665 13024 3681 13088
rect 3745 13024 3761 13088
rect 3825 13024 3833 13088
rect 3513 12474 3833 13024
rect 3513 12238 3555 12474
rect 3791 12238 3833 12474
rect 3513 12000 3833 12238
rect 3513 11936 3521 12000
rect 3585 11936 3601 12000
rect 3665 11936 3681 12000
rect 3745 11936 3761 12000
rect 3825 11936 3833 12000
rect 3513 10912 3833 11936
rect 3513 10848 3521 10912
rect 3585 10848 3601 10912
rect 3665 10848 3681 10912
rect 3745 10848 3761 10912
rect 3825 10848 3833 10912
rect 3513 9824 3833 10848
rect 3513 9760 3521 9824
rect 3585 9760 3601 9824
rect 3665 9760 3681 9824
rect 3745 9760 3761 9824
rect 3825 9760 3833 9824
rect 3513 8736 3833 9760
rect 3513 8672 3521 8736
rect 3585 8672 3601 8736
rect 3665 8672 3681 8736
rect 3745 8672 3761 8736
rect 3825 8672 3833 8736
rect 3513 8666 3833 8672
rect 3513 8430 3555 8666
rect 3791 8430 3833 8666
rect 3513 7648 3833 8430
rect 3513 7584 3521 7648
rect 3585 7584 3601 7648
rect 3665 7584 3681 7648
rect 3745 7584 3761 7648
rect 3825 7584 3833 7648
rect 3513 6560 3833 7584
rect 3513 6496 3521 6560
rect 3585 6496 3601 6560
rect 3665 6496 3681 6560
rect 3745 6496 3761 6560
rect 3825 6496 3833 6560
rect 3513 5472 3833 6496
rect 3513 5408 3521 5472
rect 3585 5408 3601 5472
rect 3665 5408 3681 5472
rect 3745 5408 3761 5472
rect 3825 5408 3833 5472
rect 3513 4858 3833 5408
rect 3513 4622 3555 4858
rect 3791 4622 3833 4858
rect 3513 4384 3833 4622
rect 3513 4320 3521 4384
rect 3585 4320 3601 4384
rect 3665 4320 3681 4384
rect 3745 4320 3761 4384
rect 3825 4320 3833 4384
rect 3513 3296 3833 4320
rect 3513 3232 3521 3296
rect 3585 3232 3601 3296
rect 3665 3232 3681 3296
rect 3745 3232 3761 3296
rect 3825 3232 3833 3296
rect 3513 2208 3833 3232
rect 3513 2144 3521 2208
rect 3585 2144 3601 2208
rect 3665 2144 3681 2208
rect 3745 2144 3761 2208
rect 3825 2144 3833 2208
rect 3513 2128 3833 2144
rect 6671 16896 6991 17456
rect 6671 16832 6679 16896
rect 6743 16832 6759 16896
rect 6823 16832 6839 16896
rect 6903 16832 6919 16896
rect 6983 16832 6991 16896
rect 6671 15808 6991 16832
rect 6671 15744 6679 15808
rect 6743 15744 6759 15808
rect 6823 15744 6839 15808
rect 6903 15744 6919 15808
rect 6983 15744 6991 15808
rect 6671 15622 6991 15744
rect 6671 15386 6713 15622
rect 6949 15386 6991 15622
rect 6671 14720 6991 15386
rect 6671 14656 6679 14720
rect 6743 14656 6759 14720
rect 6823 14656 6839 14720
rect 6903 14656 6919 14720
rect 6983 14656 6991 14720
rect 6671 13632 6991 14656
rect 6671 13568 6679 13632
rect 6743 13568 6759 13632
rect 6823 13568 6839 13632
rect 6903 13568 6919 13632
rect 6983 13568 6991 13632
rect 6671 12544 6991 13568
rect 6671 12480 6679 12544
rect 6743 12480 6759 12544
rect 6823 12480 6839 12544
rect 6903 12480 6919 12544
rect 6983 12480 6991 12544
rect 6671 11814 6991 12480
rect 6671 11578 6713 11814
rect 6949 11578 6991 11814
rect 6671 11456 6991 11578
rect 6671 11392 6679 11456
rect 6743 11392 6759 11456
rect 6823 11392 6839 11456
rect 6903 11392 6919 11456
rect 6983 11392 6991 11456
rect 6671 10368 6991 11392
rect 6671 10304 6679 10368
rect 6743 10304 6759 10368
rect 6823 10304 6839 10368
rect 6903 10304 6919 10368
rect 6983 10304 6991 10368
rect 6671 9280 6991 10304
rect 6671 9216 6679 9280
rect 6743 9216 6759 9280
rect 6823 9216 6839 9280
rect 6903 9216 6919 9280
rect 6983 9216 6991 9280
rect 6671 8192 6991 9216
rect 6671 8128 6679 8192
rect 6743 8128 6759 8192
rect 6823 8128 6839 8192
rect 6903 8128 6919 8192
rect 6983 8128 6991 8192
rect 6671 8006 6991 8128
rect 6671 7770 6713 8006
rect 6949 7770 6991 8006
rect 6671 7104 6991 7770
rect 6671 7040 6679 7104
rect 6743 7040 6759 7104
rect 6823 7040 6839 7104
rect 6903 7040 6919 7104
rect 6983 7040 6991 7104
rect 6671 6016 6991 7040
rect 6671 5952 6679 6016
rect 6743 5952 6759 6016
rect 6823 5952 6839 6016
rect 6903 5952 6919 6016
rect 6983 5952 6991 6016
rect 6671 4928 6991 5952
rect 6671 4864 6679 4928
rect 6743 4864 6759 4928
rect 6823 4864 6839 4928
rect 6903 4864 6919 4928
rect 6983 4864 6991 4928
rect 6671 4198 6991 4864
rect 6671 3962 6713 4198
rect 6949 3962 6991 4198
rect 6671 3840 6991 3962
rect 6671 3776 6679 3840
rect 6743 3776 6759 3840
rect 6823 3776 6839 3840
rect 6903 3776 6919 3840
rect 6983 3776 6991 3840
rect 6671 2752 6991 3776
rect 6671 2688 6679 2752
rect 6743 2688 6759 2752
rect 6823 2688 6839 2752
rect 6903 2688 6919 2752
rect 6983 2688 6991 2752
rect 6671 2128 6991 2688
rect 7331 17440 7651 17456
rect 7331 17376 7339 17440
rect 7403 17376 7419 17440
rect 7483 17376 7499 17440
rect 7563 17376 7579 17440
rect 7643 17376 7651 17440
rect 7331 16352 7651 17376
rect 7331 16288 7339 16352
rect 7403 16288 7419 16352
rect 7483 16288 7499 16352
rect 7563 16288 7579 16352
rect 7643 16288 7651 16352
rect 7331 16282 7651 16288
rect 7331 16046 7373 16282
rect 7609 16046 7651 16282
rect 7331 15264 7651 16046
rect 7331 15200 7339 15264
rect 7403 15200 7419 15264
rect 7483 15200 7499 15264
rect 7563 15200 7579 15264
rect 7643 15200 7651 15264
rect 7331 14176 7651 15200
rect 7331 14112 7339 14176
rect 7403 14112 7419 14176
rect 7483 14112 7499 14176
rect 7563 14112 7579 14176
rect 7643 14112 7651 14176
rect 7331 13088 7651 14112
rect 7331 13024 7339 13088
rect 7403 13024 7419 13088
rect 7483 13024 7499 13088
rect 7563 13024 7579 13088
rect 7643 13024 7651 13088
rect 7331 12474 7651 13024
rect 7331 12238 7373 12474
rect 7609 12238 7651 12474
rect 7331 12000 7651 12238
rect 7331 11936 7339 12000
rect 7403 11936 7419 12000
rect 7483 11936 7499 12000
rect 7563 11936 7579 12000
rect 7643 11936 7651 12000
rect 7331 10912 7651 11936
rect 7331 10848 7339 10912
rect 7403 10848 7419 10912
rect 7483 10848 7499 10912
rect 7563 10848 7579 10912
rect 7643 10848 7651 10912
rect 7331 9824 7651 10848
rect 7331 9760 7339 9824
rect 7403 9760 7419 9824
rect 7483 9760 7499 9824
rect 7563 9760 7579 9824
rect 7643 9760 7651 9824
rect 7331 8736 7651 9760
rect 7331 8672 7339 8736
rect 7403 8672 7419 8736
rect 7483 8672 7499 8736
rect 7563 8672 7579 8736
rect 7643 8672 7651 8736
rect 7331 8666 7651 8672
rect 7331 8430 7373 8666
rect 7609 8430 7651 8666
rect 7331 7648 7651 8430
rect 7331 7584 7339 7648
rect 7403 7584 7419 7648
rect 7483 7584 7499 7648
rect 7563 7584 7579 7648
rect 7643 7584 7651 7648
rect 7331 6560 7651 7584
rect 7331 6496 7339 6560
rect 7403 6496 7419 6560
rect 7483 6496 7499 6560
rect 7563 6496 7579 6560
rect 7643 6496 7651 6560
rect 7331 5472 7651 6496
rect 7331 5408 7339 5472
rect 7403 5408 7419 5472
rect 7483 5408 7499 5472
rect 7563 5408 7579 5472
rect 7643 5408 7651 5472
rect 7331 4858 7651 5408
rect 7331 4622 7373 4858
rect 7609 4622 7651 4858
rect 7331 4384 7651 4622
rect 7331 4320 7339 4384
rect 7403 4320 7419 4384
rect 7483 4320 7499 4384
rect 7563 4320 7579 4384
rect 7643 4320 7651 4384
rect 7331 3296 7651 4320
rect 7331 3232 7339 3296
rect 7403 3232 7419 3296
rect 7483 3232 7499 3296
rect 7563 3232 7579 3296
rect 7643 3232 7651 3296
rect 7331 2208 7651 3232
rect 7331 2144 7339 2208
rect 7403 2144 7419 2208
rect 7483 2144 7499 2208
rect 7563 2144 7579 2208
rect 7643 2144 7651 2208
rect 7331 2128 7651 2144
rect 10489 16896 10809 17456
rect 10489 16832 10497 16896
rect 10561 16832 10577 16896
rect 10641 16832 10657 16896
rect 10721 16832 10737 16896
rect 10801 16832 10809 16896
rect 10489 15808 10809 16832
rect 10489 15744 10497 15808
rect 10561 15744 10577 15808
rect 10641 15744 10657 15808
rect 10721 15744 10737 15808
rect 10801 15744 10809 15808
rect 10489 15622 10809 15744
rect 10489 15386 10531 15622
rect 10767 15386 10809 15622
rect 10489 14720 10809 15386
rect 10489 14656 10497 14720
rect 10561 14656 10577 14720
rect 10641 14656 10657 14720
rect 10721 14656 10737 14720
rect 10801 14656 10809 14720
rect 10489 13632 10809 14656
rect 10489 13568 10497 13632
rect 10561 13568 10577 13632
rect 10641 13568 10657 13632
rect 10721 13568 10737 13632
rect 10801 13568 10809 13632
rect 10489 12544 10809 13568
rect 10489 12480 10497 12544
rect 10561 12480 10577 12544
rect 10641 12480 10657 12544
rect 10721 12480 10737 12544
rect 10801 12480 10809 12544
rect 10489 11814 10809 12480
rect 10489 11578 10531 11814
rect 10767 11578 10809 11814
rect 10489 11456 10809 11578
rect 10489 11392 10497 11456
rect 10561 11392 10577 11456
rect 10641 11392 10657 11456
rect 10721 11392 10737 11456
rect 10801 11392 10809 11456
rect 10489 10368 10809 11392
rect 10489 10304 10497 10368
rect 10561 10304 10577 10368
rect 10641 10304 10657 10368
rect 10721 10304 10737 10368
rect 10801 10304 10809 10368
rect 10489 9280 10809 10304
rect 10489 9216 10497 9280
rect 10561 9216 10577 9280
rect 10641 9216 10657 9280
rect 10721 9216 10737 9280
rect 10801 9216 10809 9280
rect 10489 8192 10809 9216
rect 10489 8128 10497 8192
rect 10561 8128 10577 8192
rect 10641 8128 10657 8192
rect 10721 8128 10737 8192
rect 10801 8128 10809 8192
rect 10489 8006 10809 8128
rect 10489 7770 10531 8006
rect 10767 7770 10809 8006
rect 10489 7104 10809 7770
rect 10489 7040 10497 7104
rect 10561 7040 10577 7104
rect 10641 7040 10657 7104
rect 10721 7040 10737 7104
rect 10801 7040 10809 7104
rect 10489 6016 10809 7040
rect 10489 5952 10497 6016
rect 10561 5952 10577 6016
rect 10641 5952 10657 6016
rect 10721 5952 10737 6016
rect 10801 5952 10809 6016
rect 10489 4928 10809 5952
rect 10489 4864 10497 4928
rect 10561 4864 10577 4928
rect 10641 4864 10657 4928
rect 10721 4864 10737 4928
rect 10801 4864 10809 4928
rect 10489 4198 10809 4864
rect 10489 3962 10531 4198
rect 10767 3962 10809 4198
rect 10489 3840 10809 3962
rect 10489 3776 10497 3840
rect 10561 3776 10577 3840
rect 10641 3776 10657 3840
rect 10721 3776 10737 3840
rect 10801 3776 10809 3840
rect 10489 2752 10809 3776
rect 10489 2688 10497 2752
rect 10561 2688 10577 2752
rect 10641 2688 10657 2752
rect 10721 2688 10737 2752
rect 10801 2688 10809 2752
rect 10489 2128 10809 2688
rect 11149 17440 11469 17456
rect 11149 17376 11157 17440
rect 11221 17376 11237 17440
rect 11301 17376 11317 17440
rect 11381 17376 11397 17440
rect 11461 17376 11469 17440
rect 11149 16352 11469 17376
rect 11149 16288 11157 16352
rect 11221 16288 11237 16352
rect 11301 16288 11317 16352
rect 11381 16288 11397 16352
rect 11461 16288 11469 16352
rect 11149 16282 11469 16288
rect 11149 16046 11191 16282
rect 11427 16046 11469 16282
rect 11149 15264 11469 16046
rect 11149 15200 11157 15264
rect 11221 15200 11237 15264
rect 11301 15200 11317 15264
rect 11381 15200 11397 15264
rect 11461 15200 11469 15264
rect 11149 14176 11469 15200
rect 11149 14112 11157 14176
rect 11221 14112 11237 14176
rect 11301 14112 11317 14176
rect 11381 14112 11397 14176
rect 11461 14112 11469 14176
rect 11149 13088 11469 14112
rect 11149 13024 11157 13088
rect 11221 13024 11237 13088
rect 11301 13024 11317 13088
rect 11381 13024 11397 13088
rect 11461 13024 11469 13088
rect 11149 12474 11469 13024
rect 11149 12238 11191 12474
rect 11427 12238 11469 12474
rect 11149 12000 11469 12238
rect 11149 11936 11157 12000
rect 11221 11936 11237 12000
rect 11301 11936 11317 12000
rect 11381 11936 11397 12000
rect 11461 11936 11469 12000
rect 11149 10912 11469 11936
rect 11149 10848 11157 10912
rect 11221 10848 11237 10912
rect 11301 10848 11317 10912
rect 11381 10848 11397 10912
rect 11461 10848 11469 10912
rect 11149 9824 11469 10848
rect 11149 9760 11157 9824
rect 11221 9760 11237 9824
rect 11301 9760 11317 9824
rect 11381 9760 11397 9824
rect 11461 9760 11469 9824
rect 11149 8736 11469 9760
rect 11149 8672 11157 8736
rect 11221 8672 11237 8736
rect 11301 8672 11317 8736
rect 11381 8672 11397 8736
rect 11461 8672 11469 8736
rect 11149 8666 11469 8672
rect 11149 8430 11191 8666
rect 11427 8430 11469 8666
rect 11149 7648 11469 8430
rect 11149 7584 11157 7648
rect 11221 7584 11237 7648
rect 11301 7584 11317 7648
rect 11381 7584 11397 7648
rect 11461 7584 11469 7648
rect 11149 6560 11469 7584
rect 11149 6496 11157 6560
rect 11221 6496 11237 6560
rect 11301 6496 11317 6560
rect 11381 6496 11397 6560
rect 11461 6496 11469 6560
rect 11149 5472 11469 6496
rect 11149 5408 11157 5472
rect 11221 5408 11237 5472
rect 11301 5408 11317 5472
rect 11381 5408 11397 5472
rect 11461 5408 11469 5472
rect 11149 4858 11469 5408
rect 11149 4622 11191 4858
rect 11427 4622 11469 4858
rect 11149 4384 11469 4622
rect 11149 4320 11157 4384
rect 11221 4320 11237 4384
rect 11301 4320 11317 4384
rect 11381 4320 11397 4384
rect 11461 4320 11469 4384
rect 11149 3296 11469 4320
rect 11149 3232 11157 3296
rect 11221 3232 11237 3296
rect 11301 3232 11317 3296
rect 11381 3232 11397 3296
rect 11461 3232 11469 3296
rect 11149 2208 11469 3232
rect 11149 2144 11157 2208
rect 11221 2144 11237 2208
rect 11301 2144 11317 2208
rect 11381 2144 11397 2208
rect 11461 2144 11469 2208
rect 11149 2128 11469 2144
rect 14307 16896 14627 17456
rect 14307 16832 14315 16896
rect 14379 16832 14395 16896
rect 14459 16832 14475 16896
rect 14539 16832 14555 16896
rect 14619 16832 14627 16896
rect 14307 15808 14627 16832
rect 14307 15744 14315 15808
rect 14379 15744 14395 15808
rect 14459 15744 14475 15808
rect 14539 15744 14555 15808
rect 14619 15744 14627 15808
rect 14307 15622 14627 15744
rect 14307 15386 14349 15622
rect 14585 15386 14627 15622
rect 14307 14720 14627 15386
rect 14307 14656 14315 14720
rect 14379 14656 14395 14720
rect 14459 14656 14475 14720
rect 14539 14656 14555 14720
rect 14619 14656 14627 14720
rect 14307 13632 14627 14656
rect 14307 13568 14315 13632
rect 14379 13568 14395 13632
rect 14459 13568 14475 13632
rect 14539 13568 14555 13632
rect 14619 13568 14627 13632
rect 14307 12544 14627 13568
rect 14307 12480 14315 12544
rect 14379 12480 14395 12544
rect 14459 12480 14475 12544
rect 14539 12480 14555 12544
rect 14619 12480 14627 12544
rect 14307 11814 14627 12480
rect 14307 11578 14349 11814
rect 14585 11578 14627 11814
rect 14307 11456 14627 11578
rect 14307 11392 14315 11456
rect 14379 11392 14395 11456
rect 14459 11392 14475 11456
rect 14539 11392 14555 11456
rect 14619 11392 14627 11456
rect 14307 10368 14627 11392
rect 14307 10304 14315 10368
rect 14379 10304 14395 10368
rect 14459 10304 14475 10368
rect 14539 10304 14555 10368
rect 14619 10304 14627 10368
rect 14307 9280 14627 10304
rect 14307 9216 14315 9280
rect 14379 9216 14395 9280
rect 14459 9216 14475 9280
rect 14539 9216 14555 9280
rect 14619 9216 14627 9280
rect 14307 8192 14627 9216
rect 14307 8128 14315 8192
rect 14379 8128 14395 8192
rect 14459 8128 14475 8192
rect 14539 8128 14555 8192
rect 14619 8128 14627 8192
rect 14307 8006 14627 8128
rect 14307 7770 14349 8006
rect 14585 7770 14627 8006
rect 14307 7104 14627 7770
rect 14307 7040 14315 7104
rect 14379 7040 14395 7104
rect 14459 7040 14475 7104
rect 14539 7040 14555 7104
rect 14619 7040 14627 7104
rect 14307 6016 14627 7040
rect 14307 5952 14315 6016
rect 14379 5952 14395 6016
rect 14459 5952 14475 6016
rect 14539 5952 14555 6016
rect 14619 5952 14627 6016
rect 14307 4928 14627 5952
rect 14307 4864 14315 4928
rect 14379 4864 14395 4928
rect 14459 4864 14475 4928
rect 14539 4864 14555 4928
rect 14619 4864 14627 4928
rect 14307 4198 14627 4864
rect 14307 3962 14349 4198
rect 14585 3962 14627 4198
rect 14307 3840 14627 3962
rect 14307 3776 14315 3840
rect 14379 3776 14395 3840
rect 14459 3776 14475 3840
rect 14539 3776 14555 3840
rect 14619 3776 14627 3840
rect 14307 2752 14627 3776
rect 14307 2688 14315 2752
rect 14379 2688 14395 2752
rect 14459 2688 14475 2752
rect 14539 2688 14555 2752
rect 14619 2688 14627 2752
rect 14307 2128 14627 2688
rect 14967 17440 15287 17456
rect 14967 17376 14975 17440
rect 15039 17376 15055 17440
rect 15119 17376 15135 17440
rect 15199 17376 15215 17440
rect 15279 17376 15287 17440
rect 14967 16352 15287 17376
rect 14967 16288 14975 16352
rect 15039 16288 15055 16352
rect 15119 16288 15135 16352
rect 15199 16288 15215 16352
rect 15279 16288 15287 16352
rect 14967 16282 15287 16288
rect 14967 16046 15009 16282
rect 15245 16046 15287 16282
rect 14967 15264 15287 16046
rect 14967 15200 14975 15264
rect 15039 15200 15055 15264
rect 15119 15200 15135 15264
rect 15199 15200 15215 15264
rect 15279 15200 15287 15264
rect 14967 14176 15287 15200
rect 14967 14112 14975 14176
rect 15039 14112 15055 14176
rect 15119 14112 15135 14176
rect 15199 14112 15215 14176
rect 15279 14112 15287 14176
rect 14967 13088 15287 14112
rect 14967 13024 14975 13088
rect 15039 13024 15055 13088
rect 15119 13024 15135 13088
rect 15199 13024 15215 13088
rect 15279 13024 15287 13088
rect 14967 12474 15287 13024
rect 14967 12238 15009 12474
rect 15245 12238 15287 12474
rect 14967 12000 15287 12238
rect 14967 11936 14975 12000
rect 15039 11936 15055 12000
rect 15119 11936 15135 12000
rect 15199 11936 15215 12000
rect 15279 11936 15287 12000
rect 14967 10912 15287 11936
rect 14967 10848 14975 10912
rect 15039 10848 15055 10912
rect 15119 10848 15135 10912
rect 15199 10848 15215 10912
rect 15279 10848 15287 10912
rect 14967 9824 15287 10848
rect 14967 9760 14975 9824
rect 15039 9760 15055 9824
rect 15119 9760 15135 9824
rect 15199 9760 15215 9824
rect 15279 9760 15287 9824
rect 14967 8736 15287 9760
rect 14967 8672 14975 8736
rect 15039 8672 15055 8736
rect 15119 8672 15135 8736
rect 15199 8672 15215 8736
rect 15279 8672 15287 8736
rect 14967 8666 15287 8672
rect 14967 8430 15009 8666
rect 15245 8430 15287 8666
rect 14967 7648 15287 8430
rect 14967 7584 14975 7648
rect 15039 7584 15055 7648
rect 15119 7584 15135 7648
rect 15199 7584 15215 7648
rect 15279 7584 15287 7648
rect 14967 6560 15287 7584
rect 14967 6496 14975 6560
rect 15039 6496 15055 6560
rect 15119 6496 15135 6560
rect 15199 6496 15215 6560
rect 15279 6496 15287 6560
rect 14967 5472 15287 6496
rect 14967 5408 14975 5472
rect 15039 5408 15055 5472
rect 15119 5408 15135 5472
rect 15199 5408 15215 5472
rect 15279 5408 15287 5472
rect 14967 4858 15287 5408
rect 14967 4622 15009 4858
rect 15245 4622 15287 4858
rect 14967 4384 15287 4622
rect 14967 4320 14975 4384
rect 15039 4320 15055 4384
rect 15119 4320 15135 4384
rect 15199 4320 15215 4384
rect 15279 4320 15287 4384
rect 14967 3296 15287 4320
rect 14967 3232 14975 3296
rect 15039 3232 15055 3296
rect 15119 3232 15135 3296
rect 15199 3232 15215 3296
rect 15279 3232 15287 3296
rect 14967 2208 15287 3232
rect 14967 2144 14975 2208
rect 15039 2144 15055 2208
rect 15119 2144 15135 2208
rect 15199 2144 15215 2208
rect 15279 2144 15287 2208
rect 14967 2128 15287 2144
<< via4 >>
rect 2895 15386 3131 15622
rect 2895 11578 3131 11814
rect 2895 7770 3131 8006
rect 2895 3962 3131 4198
rect 3555 16046 3791 16282
rect 3555 12238 3791 12474
rect 3555 8430 3791 8666
rect 3555 4622 3791 4858
rect 6713 15386 6949 15622
rect 6713 11578 6949 11814
rect 6713 7770 6949 8006
rect 6713 3962 6949 4198
rect 7373 16046 7609 16282
rect 7373 12238 7609 12474
rect 7373 8430 7609 8666
rect 7373 4622 7609 4858
rect 10531 15386 10767 15622
rect 10531 11578 10767 11814
rect 10531 7770 10767 8006
rect 10531 3962 10767 4198
rect 11191 16046 11427 16282
rect 11191 12238 11427 12474
rect 11191 8430 11427 8666
rect 11191 4622 11427 4858
rect 14349 15386 14585 15622
rect 14349 11578 14585 11814
rect 14349 7770 14585 8006
rect 14349 3962 14585 4198
rect 15009 16046 15245 16282
rect 15009 12238 15245 12474
rect 15009 8430 15245 8666
rect 15009 4622 15245 4858
<< metal5 >>
rect 1056 16282 16424 16324
rect 1056 16046 3555 16282
rect 3791 16046 7373 16282
rect 7609 16046 11191 16282
rect 11427 16046 15009 16282
rect 15245 16046 16424 16282
rect 1056 16004 16424 16046
rect 1056 15622 16424 15664
rect 1056 15386 2895 15622
rect 3131 15386 6713 15622
rect 6949 15386 10531 15622
rect 10767 15386 14349 15622
rect 14585 15386 16424 15622
rect 1056 15344 16424 15386
rect 1056 12474 16424 12516
rect 1056 12238 3555 12474
rect 3791 12238 7373 12474
rect 7609 12238 11191 12474
rect 11427 12238 15009 12474
rect 15245 12238 16424 12474
rect 1056 12196 16424 12238
rect 1056 11814 16424 11856
rect 1056 11578 2895 11814
rect 3131 11578 6713 11814
rect 6949 11578 10531 11814
rect 10767 11578 14349 11814
rect 14585 11578 16424 11814
rect 1056 11536 16424 11578
rect 1056 8666 16424 8708
rect 1056 8430 3555 8666
rect 3791 8430 7373 8666
rect 7609 8430 11191 8666
rect 11427 8430 15009 8666
rect 15245 8430 16424 8666
rect 1056 8388 16424 8430
rect 1056 8006 16424 8048
rect 1056 7770 2895 8006
rect 3131 7770 6713 8006
rect 6949 7770 10531 8006
rect 10767 7770 14349 8006
rect 14585 7770 16424 8006
rect 1056 7728 16424 7770
rect 1056 4858 16424 4900
rect 1056 4622 3555 4858
rect 3791 4622 7373 4858
rect 7609 4622 11191 4858
rect 11427 4622 15009 4858
rect 15245 4622 16424 4858
rect 1056 4580 16424 4622
rect 1056 4198 16424 4240
rect 1056 3962 2895 4198
rect 3131 3962 6713 4198
rect 6949 3962 10531 4198
rect 10767 3962 14349 4198
rect 14585 3962 16424 4198
rect 1056 3920 16424 3962
use sky130_fd_sc_hd__mux2_1  _14_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 4784 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _15_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 5060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _16_
timestamp 1694700623
transform -1 0 6164 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _17_
timestamp 1694700623
transform -1 0 5336 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _18_
timestamp 1694700623
transform -1 0 7268 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _19_
timestamp 1694700623
transform 1 0 6808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _20_
timestamp 1694700623
transform 1 0 7820 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _21_
timestamp 1694700623
transform 1 0 7268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _22_
timestamp 1694700623
transform 1 0 9108 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 1694700623
transform -1 0 8832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _24_
timestamp 1694700623
transform -1 0 10856 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _25_
timestamp 1694700623
transform 1 0 11408 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _26_
timestamp 1694700623
transform 1 0 9844 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _27_
timestamp 1694700623
transform -1 0 9384 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _28_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 6256 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _29_
timestamp 1694700623
transform 1 0 4968 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _30_
timestamp 1694700623
transform 1 0 4416 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _31_
timestamp 1694700623
transform 1 0 6624 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _32_
timestamp 1694700623
transform -1 0 9108 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _33_
timestamp 1694700623
transform 1 0 9108 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _34_
timestamp 1694700623
transform 1 0 9384 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_sclk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 7268 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_sclk
timestamp 1694700623
transform -1 0 6624 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_sclk
timestamp 1694700623
transform 1 0 9568 0 1 3264
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_35
timestamp 1694700623
transform 1 0 4324 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_82
timestamp 1694700623
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 1694700623
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_96
timestamp 1694700623
transform 1 0 9936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_117
timestamp 1694700623
transform 1 0 11868 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_124
timestamp 1694700623
transform 1 0 12512 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_136
timestamp 1694700623
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_147
timestamp 1694700623
transform 1 0 14628 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_159
timestamp 1694700623
transform 1 0 15732 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1694700623
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1694700623
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_27
timestamp 1694700623
transform 1 0 3588 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_57
timestamp 1694700623
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_107
timestamp 1694700623
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1694700623
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_121
timestamp 1694700623
transform 1 0 12236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_133
timestamp 1694700623
transform 1 0 13340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_145
timestamp 1694700623
transform 1 0 14444 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_157
timestamp 1694700623
transform 1 0 15548 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1694700623
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1694700623
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1694700623
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_29
timestamp 1694700623
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_80
timestamp 1694700623
transform 1 0 8464 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_85
timestamp 1694700623
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_91
timestamp 1694700623
transform 1 0 9476 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_115
timestamp 1694700623
transform 1 0 11684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_127
timestamp 1694700623
transform 1 0 12788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1694700623
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1694700623
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_153 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 15180 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_161
timestamp 1694700623
transform 1 0 15916 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1694700623
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1694700623
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1694700623
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_39
timestamp 1694700623
transform 1 0 4692 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1694700623
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_65
timestamp 1694700623
transform 1 0 7084 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_110
timestamp 1694700623
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1694700623
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1694700623
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1694700623
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1694700623
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_161
timestamp 1694700623
transform 1 0 15916 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1694700623
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1694700623
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1694700623
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1694700623
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_41
timestamp 1694700623
transform 1 0 4876 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_65
timestamp 1694700623
transform 1 0 7084 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_82
timestamp 1694700623
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_85
timestamp 1694700623
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_93
timestamp 1694700623
transform 1 0 9660 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_104
timestamp 1694700623
transform 1 0 10672 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_116
timestamp 1694700623
transform 1 0 11776 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_128
timestamp 1694700623
transform 1 0 12880 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1694700623
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_153
timestamp 1694700623
transform 1 0 15180 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_161
timestamp 1694700623
transform 1 0 15916 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1694700623
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1694700623
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1694700623
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_39
timestamp 1694700623
transform 1 0 4692 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1694700623
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_69
timestamp 1694700623
transform 1 0 7452 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1694700623
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1694700623
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1694700623
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1694700623
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1694700623
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1694700623
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1694700623
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1694700623
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_161
timestamp 1694700623
transform 1 0 15916 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1694700623
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1694700623
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1694700623
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1694700623
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1694700623
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1694700623
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1694700623
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1694700623
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1694700623
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1694700623
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1694700623
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1694700623
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1694700623
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1694700623
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1694700623
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1694700623
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_153
timestamp 1694700623
transform 1 0 15180 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_161
timestamp 1694700623
transform 1 0 15916 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1694700623
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1694700623
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1694700623
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1694700623
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1694700623
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1694700623
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1694700623
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1694700623
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1694700623
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1694700623
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1694700623
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1694700623
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1694700623
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1694700623
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1694700623
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1694700623
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_161
timestamp 1694700623
transform 1 0 15916 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1694700623
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1694700623
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1694700623
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1694700623
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1694700623
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1694700623
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1694700623
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1694700623
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1694700623
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1694700623
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1694700623
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1694700623
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1694700623
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1694700623
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1694700623
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1694700623
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_153
timestamp 1694700623
transform 1 0 15180 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_161
timestamp 1694700623
transform 1 0 15916 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1694700623
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1694700623
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1694700623
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1694700623
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1694700623
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1694700623
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1694700623
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1694700623
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1694700623
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1694700623
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1694700623
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1694700623
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1694700623
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1694700623
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1694700623
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1694700623
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_161
timestamp 1694700623
transform 1 0 15916 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1694700623
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1694700623
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1694700623
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1694700623
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1694700623
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1694700623
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1694700623
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1694700623
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1694700623
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1694700623
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1694700623
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1694700623
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1694700623
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1694700623
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1694700623
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1694700623
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_153
timestamp 1694700623
transform 1 0 15180 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_161
timestamp 1694700623
transform 1 0 15916 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1694700623
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1694700623
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1694700623
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1694700623
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1694700623
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1694700623
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1694700623
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1694700623
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1694700623
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1694700623
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1694700623
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1694700623
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1694700623
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1694700623
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1694700623
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1694700623
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_161
timestamp 1694700623
transform 1 0 15916 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1694700623
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1694700623
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1694700623
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1694700623
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1694700623
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1694700623
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1694700623
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1694700623
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1694700623
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1694700623
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1694700623
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1694700623
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1694700623
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1694700623
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1694700623
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1694700623
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_153
timestamp 1694700623
transform 1 0 15180 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_161
timestamp 1694700623
transform 1 0 15916 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1694700623
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1694700623
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1694700623
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1694700623
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1694700623
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1694700623
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1694700623
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1694700623
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1694700623
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1694700623
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1694700623
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1694700623
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1694700623
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1694700623
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1694700623
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1694700623
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_161
timestamp 1694700623
transform 1 0 15916 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1694700623
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1694700623
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1694700623
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1694700623
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1694700623
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1694700623
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1694700623
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1694700623
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1694700623
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1694700623
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1694700623
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1694700623
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1694700623
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1694700623
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1694700623
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1694700623
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_153
timestamp 1694700623
transform 1 0 15180 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_161
timestamp 1694700623
transform 1 0 15916 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1694700623
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1694700623
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1694700623
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1694700623
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1694700623
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1694700623
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1694700623
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1694700623
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1694700623
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1694700623
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1694700623
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1694700623
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1694700623
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1694700623
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1694700623
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1694700623
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_161
timestamp 1694700623
transform 1 0 15916 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1694700623
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1694700623
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1694700623
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1694700623
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1694700623
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1694700623
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1694700623
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1694700623
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1694700623
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1694700623
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1694700623
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1694700623
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1694700623
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1694700623
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1694700623
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1694700623
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_153
timestamp 1694700623
transform 1 0 15180 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_161
timestamp 1694700623
transform 1 0 15916 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1694700623
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1694700623
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1694700623
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1694700623
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1694700623
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1694700623
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1694700623
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1694700623
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1694700623
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1694700623
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1694700623
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1694700623
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1694700623
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1694700623
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1694700623
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 1694700623
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_161
timestamp 1694700623
transform 1 0 15916 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1694700623
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1694700623
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1694700623
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1694700623
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1694700623
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1694700623
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1694700623
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1694700623
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1694700623
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1694700623
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1694700623
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1694700623
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1694700623
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1694700623
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1694700623
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1694700623
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_153
timestamp 1694700623
transform 1 0 15180 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_161
timestamp 1694700623
transform 1 0 15916 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1694700623
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1694700623
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1694700623
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1694700623
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1694700623
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1694700623
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1694700623
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1694700623
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1694700623
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1694700623
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1694700623
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1694700623
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1694700623
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1694700623
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1694700623
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 1694700623
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_161
timestamp 1694700623
transform 1 0 15916 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1694700623
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1694700623
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1694700623
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1694700623
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1694700623
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1694700623
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1694700623
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1694700623
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1694700623
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1694700623
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1694700623
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 1694700623
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 1694700623
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 1694700623
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1694700623
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1694700623
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_153
timestamp 1694700623
transform 1 0 15180 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_161
timestamp 1694700623
transform 1 0 15916 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1694700623
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1694700623
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1694700623
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1694700623
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1694700623
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1694700623
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1694700623
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1694700623
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1694700623
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1694700623
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1694700623
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1694700623
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1694700623
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1694700623
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 1694700623
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 1694700623
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_161
timestamp 1694700623
transform 1 0 15916 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1694700623
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1694700623
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1694700623
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1694700623
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1694700623
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1694700623
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1694700623
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1694700623
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1694700623
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1694700623
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1694700623
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1694700623
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 1694700623
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1694700623
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1694700623
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1694700623
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_153
timestamp 1694700623
transform 1 0 15180 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_161
timestamp 1694700623
transform 1 0 15916 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1694700623
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1694700623
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1694700623
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1694700623
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1694700623
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1694700623
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1694700623
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1694700623
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1694700623
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1694700623
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1694700623
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1694700623
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1694700623
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1694700623
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 1694700623
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 1694700623
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_161
timestamp 1694700623
transform 1 0 15916 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1694700623
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1694700623
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1694700623
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1694700623
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1694700623
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1694700623
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1694700623
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1694700623
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1694700623
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1694700623
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1694700623
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1694700623
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1694700623
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1694700623
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1694700623
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1694700623
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_153
timestamp 1694700623
transform 1 0 15180 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_161
timestamp 1694700623
transform 1 0 15916 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1694700623
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1694700623
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1694700623
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1694700623
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1694700623
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1694700623
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1694700623
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1694700623
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1694700623
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1694700623
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1694700623
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1694700623
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1694700623
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1694700623
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 1694700623
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1694700623
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_161
timestamp 1694700623
transform 1 0 15916 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1694700623
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1694700623
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1694700623
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1694700623
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1694700623
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1694700623
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1694700623
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1694700623
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1694700623
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1694700623
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1694700623
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1694700623
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1694700623
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1694700623
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1694700623
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1694700623
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_153
timestamp 1694700623
transform 1 0 15180 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_161
timestamp 1694700623
transform 1 0 15916 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_3
timestamp 1694700623
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_11
timestamp 1694700623
transform 1 0 2116 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_19
timestamp 1694700623
transform 1 0 2852 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_27
timestamp 1694700623
transform 1 0 3588 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_29
timestamp 1694700623
transform 1 0 3772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_41
timestamp 1694700623
transform 1 0 4876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_53
timestamp 1694700623
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1694700623
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1694700623
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_81
timestamp 1694700623
transform 1 0 8556 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_85
timestamp 1694700623
transform 1 0 8924 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_97
timestamp 1694700623
transform 1 0 10028 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_105
timestamp 1694700623
transform 1 0 10764 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_110
timestamp 1694700623
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1694700623
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1694700623
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_137
timestamp 1694700623
transform 1 0 13708 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_141
timestamp 1694700623
transform 1 0 14076 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_153
timestamp 1694700623
transform 1 0 15180 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_160
timestamp 1694700623
transform 1 0 15824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3680 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1694700623
transform -1 0 7084 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1694700623
transform -1 0 5980 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1694700623
transform -1 0 8556 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1694700623
transform -1 0 12236 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1694700623
transform -1 0 7268 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 15272 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 11224 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input3
timestamp 1694700623
transform 1 0 2300 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output4
timestamp 1694700623
transform -1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output5
timestamp 1694700623
transform -1 0 4324 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output6
timestamp 1694700623
transform 1 0 8096 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output7
timestamp 1694700623
transform -1 0 8096 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output8
timestamp 1694700623
transform 1 0 10856 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output9
timestamp 1694700623
transform 1 0 11960 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output10
timestamp 1694700623
transform 1 0 14076 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_28
timestamp 1694700623
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1694700623
transform -1 0 16376 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_29
timestamp 1694700623
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1694700623
transform -1 0 16376 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_30
timestamp 1694700623
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1694700623
transform -1 0 16376 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_31
timestamp 1694700623
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1694700623
transform -1 0 16376 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_32
timestamp 1694700623
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1694700623
transform -1 0 16376 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_33
timestamp 1694700623
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1694700623
transform -1 0 16376 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_34
timestamp 1694700623
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1694700623
transform -1 0 16376 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_35
timestamp 1694700623
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1694700623
transform -1 0 16376 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_36
timestamp 1694700623
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1694700623
transform -1 0 16376 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_37
timestamp 1694700623
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1694700623
transform -1 0 16376 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_38
timestamp 1694700623
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1694700623
transform -1 0 16376 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_39
timestamp 1694700623
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1694700623
transform -1 0 16376 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_40
timestamp 1694700623
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1694700623
transform -1 0 16376 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_41
timestamp 1694700623
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1694700623
transform -1 0 16376 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_42
timestamp 1694700623
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1694700623
transform -1 0 16376 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_43
timestamp 1694700623
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1694700623
transform -1 0 16376 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_44
timestamp 1694700623
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1694700623
transform -1 0 16376 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_45
timestamp 1694700623
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1694700623
transform -1 0 16376 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_46
timestamp 1694700623
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1694700623
transform -1 0 16376 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_47
timestamp 1694700623
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1694700623
transform -1 0 16376 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_48
timestamp 1694700623
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1694700623
transform -1 0 16376 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_49
timestamp 1694700623
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1694700623
transform -1 0 16376 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_50
timestamp 1694700623
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1694700623
transform -1 0 16376 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_51
timestamp 1694700623
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1694700623
transform -1 0 16376 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_52
timestamp 1694700623
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1694700623
transform -1 0 16376 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_53
timestamp 1694700623
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1694700623
transform -1 0 16376 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_54
timestamp 1694700623
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1694700623
transform -1 0 16376 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_55
timestamp 1694700623
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1694700623
transform -1 0 16376 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sr_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 15824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_57
timestamp 1694700623
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_58
timestamp 1694700623
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_59
timestamp 1694700623
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_60
timestamp 1694700623
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_61
timestamp 1694700623
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_62
timestamp 1694700623
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_63
timestamp 1694700623
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_64
timestamp 1694700623
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_65
timestamp 1694700623
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_66
timestamp 1694700623
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_67
timestamp 1694700623
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_68
timestamp 1694700623
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_69
timestamp 1694700623
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_70
timestamp 1694700623
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_71
timestamp 1694700623
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_72
timestamp 1694700623
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_73
timestamp 1694700623
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_74
timestamp 1694700623
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_75
timestamp 1694700623
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_76
timestamp 1694700623
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_77
timestamp 1694700623
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_78
timestamp 1694700623
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_79
timestamp 1694700623
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_80
timestamp 1694700623
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_81
timestamp 1694700623
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_82
timestamp 1694700623
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_83
timestamp 1694700623
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_84
timestamp 1694700623
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_85
timestamp 1694700623
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_86
timestamp 1694700623
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_87
timestamp 1694700623
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_88
timestamp 1694700623
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_89
timestamp 1694700623
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_90
timestamp 1694700623
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_91
timestamp 1694700623
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_92
timestamp 1694700623
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_93
timestamp 1694700623
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_94
timestamp 1694700623
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_95
timestamp 1694700623
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_96
timestamp 1694700623
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_97
timestamp 1694700623
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_98
timestamp 1694700623
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_99
timestamp 1694700623
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_100
timestamp 1694700623
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_101
timestamp 1694700623
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_102
timestamp 1694700623
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_103
timestamp 1694700623
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_104
timestamp 1694700623
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_105
timestamp 1694700623
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_106
timestamp 1694700623
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_107
timestamp 1694700623
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_108
timestamp 1694700623
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_109
timestamp 1694700623
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_110
timestamp 1694700623
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_111
timestamp 1694700623
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_112
timestamp 1694700623
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_113
timestamp 1694700623
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_114
timestamp 1694700623
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_115
timestamp 1694700623
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_116
timestamp 1694700623
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_117
timestamp 1694700623
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_118
timestamp 1694700623
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_119
timestamp 1694700623
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_120
timestamp 1694700623
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_121
timestamp 1694700623
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_122
timestamp 1694700623
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_123
timestamp 1694700623
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_124
timestamp 1694700623
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_125
timestamp 1694700623
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_126
timestamp 1694700623
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_127
timestamp 1694700623
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_128
timestamp 1694700623
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_129
timestamp 1694700623
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_130
timestamp 1694700623
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
<< labels >>
flabel metal4 s 3513 2128 3833 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7331 2128 7651 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 11149 2128 11469 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 14967 2128 15287 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 4580 16424 4900 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 8388 16424 8708 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 12196 16424 12516 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 16004 16424 16324 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2853 2128 3173 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6671 2128 6991 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 10489 2128 10809 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 14307 2128 14627 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 3920 16424 4240 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 7728 16424 8048 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 11536 16424 11856 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 15344 16424 15664 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 data[0]
port 2 nsew signal tristate
flabel metal2 s 3422 0 3478 800 0 FreeSans 224 90 0 0 data[1]
port 3 nsew signal tristate
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 data[2]
port 4 nsew signal tristate
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 data[3]
port 5 nsew signal tristate
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 data[4]
port 6 nsew signal tristate
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 data[5]
port 7 nsew signal tristate
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 data[6]
port 8 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 data[7]
port 9 nsew signal tristate
flabel metal2 s 15198 18856 15254 19656 0 FreeSans 224 90 0 0 reset
port 10 nsew signal input
flabel metal2 s 6550 18856 6606 19656 0 FreeSans 224 90 0 0 sclk
port 11 nsew signal input
flabel metal2 s 10874 18856 10930 19656 0 FreeSans 224 90 0 0 sdi
port 12 nsew signal input
flabel metal2 s 2226 18856 2282 19656 0 FreeSans 224 90 0 0 ss
port 13 nsew signal input
rlabel metal1 8740 17408 8740 17408 0 VGND
rlabel metal1 8740 16864 8740 16864 0 VPWR
rlabel metal1 5520 2958 5520 2958 0 _00_
rlabel metal1 7268 2618 7268 2618 0 _01_
rlabel metal2 8786 3162 8786 3162 0 _02_
rlabel metal1 10074 2958 10074 2958 0 _03_
rlabel metal1 9614 4046 9614 4046 0 _04_
rlabel metal1 5750 2482 5750 2482 0 _05_
rlabel metal2 5290 4386 5290 4386 0 _06_
rlabel metal1 4784 3706 4784 3706 0 _07_
rlabel metal1 6026 4250 6026 4250 0 _08_
rlabel metal1 7130 2890 7130 2890 0 _09_
rlabel metal1 7682 2414 7682 2414 0 _10_
rlabel metal1 8878 2618 8878 2618 0 _11_
rlabel metal1 11224 2550 11224 2550 0 _12_
rlabel metal1 9292 4114 9292 4114 0 _13_
rlabel metal2 6578 3706 6578 3706 0 clknet_0_sclk
rlabel metal1 5060 3706 5060 3706 0 clknet_1_0__leaf_sclk
rlabel metal2 9430 3876 9430 3876 0 clknet_1_1__leaf_sclk
rlabel metal2 1334 1554 1334 1554 0 data[0]
rlabel metal2 3450 1554 3450 1554 0 data[1]
rlabel metal2 5566 959 5566 959 0 data[2]
rlabel metal2 7682 959 7682 959 0 data[3]
rlabel metal2 9798 1792 9798 1792 0 data[4]
rlabel metal2 11914 1520 11914 1520 0 data[5]
rlabel metal2 14030 1520 14030 1520 0 data[6]
rlabel metal1 5789 3026 5789 3026 0 net1
rlabel metal1 10994 2414 10994 2414 0 net10
rlabel metal2 16146 1027 16146 1027 0 net11
rlabel metal1 4324 3162 4324 3162 0 net12
rlabel metal1 6072 4114 6072 4114 0 net13
rlabel metal1 5152 4114 5152 4114 0 net14
rlabel metal1 8234 4692 8234 4692 0 net15
rlabel metal1 10948 2482 10948 2482 0 net16
rlabel metal2 6578 2856 6578 2856 0 net17
rlabel metal1 10626 16966 10626 16966 0 net2
rlabel metal1 3358 3570 3358 3570 0 net3
rlabel metal2 3726 2686 3726 2686 0 net4
rlabel metal2 5658 4352 5658 4352 0 net5
rlabel metal2 7130 3434 7130 3434 0 net6
rlabel metal1 6854 2992 6854 2992 0 net7
rlabel metal1 7866 2822 7866 2822 0 net8
rlabel metal1 11500 2958 11500 2958 0 net9
rlabel metal2 15410 18105 15410 18105 0 reset
rlabel metal2 6578 17146 6578 17146 0 sclk
rlabel metal1 11132 17170 11132 17170 0 sdi
rlabel metal1 2346 17238 2346 17238 0 ss
<< properties >>
string FIXED_BBOX 0 0 17512 19656
<< end >>
