magic
tech sky130A
magscale 1 2
timestamp 1698518340
<< error_p >>
rect -29 581 29 587
rect -29 547 -17 581
rect -29 541 29 547
rect -29 -547 29 -541
rect -29 -581 -17 -547
rect -29 -587 29 -581
<< nwell >>
rect -109 -600 109 600
<< pmos >>
rect -15 -500 15 500
<< pdiff >>
rect -73 488 -15 500
rect -73 -488 -61 488
rect -27 -488 -15 488
rect -73 -500 -15 -488
rect 15 488 73 500
rect 15 -488 27 488
rect 61 -488 73 488
rect 15 -500 73 -488
<< pdiffc >>
rect -61 -488 -27 488
rect 27 -488 61 488
<< poly >>
rect -33 581 33 597
rect -33 547 -17 581
rect 17 547 33 581
rect -33 531 33 547
rect -15 500 15 531
rect -15 -531 15 -500
rect -33 -547 33 -531
rect -33 -581 -17 -547
rect 17 -581 33 -547
rect -33 -597 33 -581
<< polycont >>
rect -17 547 17 581
rect -17 -581 17 -547
<< locali >>
rect -33 547 -17 581
rect 17 547 33 581
rect -61 488 -27 504
rect -61 -504 -27 -488
rect 27 488 61 504
rect 27 -504 61 -488
rect -33 -581 -17 -547
rect 17 -581 33 -547
<< viali >>
rect -17 547 17 581
rect -61 -17 -27 471
rect 27 -17 61 471
rect -17 -581 17 -547
<< metal1 >>
rect -29 581 29 587
rect -29 547 -17 581
rect 17 547 29 581
rect -29 541 29 547
rect -67 471 -21 483
rect -67 -17 -61 471
rect -27 -17 -21 471
rect -67 -29 -21 -17
rect 21 471 67 483
rect 21 -17 27 471
rect 61 -17 67 471
rect 21 -29 67 -17
rect -29 -547 29 -541
rect -29 -581 -17 -547
rect 17 -581 29 -547
rect -29 -587 29 -581
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc -50 viadrn -50 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
