magic
tech sky130A
magscale 1 2
timestamp 1698604040
<< nwell >>
rect 4910 26581 20258 27147
rect 4910 25493 20258 26059
rect 4910 24405 20258 24971
rect 4910 23317 20258 23883
rect 4910 22229 20258 22795
rect 4910 21141 20258 21707
rect 4910 20053 20258 20619
rect 4910 18965 20258 19531
rect 4910 17877 20258 18443
rect 4910 16789 20258 17355
rect 4910 15701 20258 16267
rect 4910 14613 20258 15179
rect 4910 13525 20258 14091
rect 4910 12437 20258 13003
rect 29520 4870 34880 7110
rect 1250 2960 3450 4520
rect 4550 2960 6750 4520
rect 7850 2960 10050 4520
rect 11150 2960 13350 4520
rect 14750 2960 16950 4520
rect 18250 2960 20450 4520
rect 21950 2960 24150 4520
rect 25750 2960 27950 4520
<< pwell >>
rect 4977 27387 5011 27425
rect 5437 27387 5471 27425
rect 5989 27387 6023 27425
rect 6092 27397 6116 27419
rect 7185 27387 7219 27425
rect 7553 27387 7587 27425
rect 8657 27387 8691 27425
rect 9761 27387 9795 27425
rect 10037 27396 10069 27418
rect 10131 27387 10165 27425
rect 10497 27396 10529 27418
rect 11233 27387 11267 27425
rect 12337 27387 12371 27425
rect 12705 27387 12739 27425
rect 13809 27387 13843 27425
rect 14913 27387 14947 27425
rect 15281 27387 15315 27425
rect 16385 27387 16419 27425
rect 17489 27387 17523 27425
rect 17684 27397 17708 27419
rect 18409 27387 18443 27425
rect 18961 27387 18995 27425
rect 19145 27396 19177 27418
rect 19881 27387 19915 27425
rect 20157 27387 20191 27425
rect 4949 27225 5223 27387
rect 5225 27225 5499 27387
rect 5503 27251 6051 27387
rect 6145 27225 7247 27387
rect 7251 27213 7337 27370
rect 7341 27225 7615 27387
rect 7617 27225 8719 27387
rect 8721 27225 9823 27387
rect 9827 27213 9913 27370
rect 10101 27231 10375 27387
rect 10561 27225 11295 27387
rect 11297 27225 12399 27387
rect 12403 27213 12489 27370
rect 12493 27225 12767 27387
rect 12769 27225 13871 27387
rect 13873 27225 14975 27387
rect 14979 27213 15065 27370
rect 15069 27225 15343 27387
rect 15345 27225 16447 27387
rect 16449 27225 17551 27387
rect 17555 27213 17641 27370
rect 17737 27225 18471 27387
rect 18475 27251 19023 27387
rect 19209 27225 19943 27387
rect 19945 27225 20219 27387
rect 4949 26341 5223 26503
rect 5409 26341 6143 26503
rect 6145 26341 7247 26503
rect 7251 26358 7337 26515
rect 7433 26341 7983 26503
rect 7985 26341 9087 26503
rect 9089 26341 10191 26503
rect 10193 26341 11295 26503
rect 11297 26341 12399 26503
rect 12403 26358 12489 26515
rect 12585 26341 13135 26503
rect 13137 26341 14239 26503
rect 14241 26341 15343 26503
rect 15345 26341 16447 26503
rect 16449 26341 17551 26503
rect 17555 26358 17641 26515
rect 17737 26341 18839 26503
rect 18841 26341 19943 26503
rect 19945 26341 20219 26503
rect 4977 26299 5011 26341
rect 5345 26308 5377 26332
rect 6081 26303 6115 26341
rect 6449 26299 6483 26337
rect 7185 26303 7219 26341
rect 7380 26309 7404 26331
rect 7553 26299 7587 26337
rect 7921 26303 7955 26341
rect 8657 26299 8691 26337
rect 9025 26303 9059 26341
rect 9761 26299 9795 26337
rect 9956 26309 9980 26331
rect 10129 26303 10163 26341
rect 10497 26299 10531 26337
rect 11233 26303 11267 26341
rect 11601 26299 11635 26337
rect 12337 26303 12371 26341
rect 12532 26309 12556 26331
rect 12705 26299 12739 26337
rect 13073 26303 13107 26341
rect 13809 26299 13843 26337
rect 14177 26303 14211 26341
rect 14913 26299 14947 26337
rect 15108 26309 15132 26331
rect 15281 26303 15315 26341
rect 15465 26299 15499 26337
rect 16385 26303 16419 26341
rect 16569 26299 16603 26337
rect 17489 26303 17523 26341
rect 17673 26331 17707 26337
rect 17673 26309 17708 26331
rect 17673 26299 17707 26309
rect 18777 26299 18811 26341
rect 19881 26299 19915 26341
rect 20157 26299 20191 26341
rect 4949 26137 5223 26299
rect 5409 26137 6511 26299
rect 6513 26137 7615 26299
rect 7617 26137 8719 26299
rect 8721 26137 9823 26299
rect 9827 26125 9913 26282
rect 10009 26137 10559 26299
rect 10561 26137 11663 26299
rect 11665 26137 12767 26299
rect 12769 26137 13871 26299
rect 13873 26137 14975 26299
rect 14979 26125 15065 26282
rect 15161 26137 15527 26299
rect 15529 26137 16631 26299
rect 16633 26137 17735 26299
rect 17737 26137 18839 26299
rect 18841 26137 19943 26299
rect 19945 26137 20219 26299
rect 4949 25253 5223 25415
rect 5409 25253 6143 25415
rect 6145 25253 7247 25415
rect 7251 25270 7337 25427
rect 7433 25253 7983 25415
rect 7985 25253 9087 25415
rect 9089 25253 10191 25415
rect 10193 25253 11295 25415
rect 11297 25253 12399 25415
rect 12403 25270 12489 25427
rect 12585 25253 13135 25415
rect 13137 25253 14239 25415
rect 14241 25253 15343 25415
rect 15345 25253 16447 25415
rect 16449 25253 17551 25415
rect 17555 25270 17641 25427
rect 17737 25253 18839 25415
rect 18841 25253 19943 25415
rect 19945 25253 20219 25415
rect 4977 25211 5011 25253
rect 5345 25220 5377 25244
rect 6081 25215 6115 25253
rect 6449 25211 6483 25249
rect 7185 25215 7219 25253
rect 7380 25221 7404 25243
rect 7553 25211 7587 25249
rect 7921 25215 7955 25253
rect 8657 25211 8691 25249
rect 9025 25215 9059 25253
rect 9761 25211 9795 25249
rect 9956 25221 9980 25243
rect 10129 25215 10163 25253
rect 10497 25211 10531 25249
rect 11233 25215 11267 25253
rect 11601 25211 11635 25249
rect 12337 25215 12371 25253
rect 12532 25221 12556 25243
rect 12705 25211 12739 25249
rect 13073 25215 13107 25253
rect 13809 25211 13843 25249
rect 14177 25215 14211 25253
rect 14913 25211 14947 25249
rect 15108 25221 15132 25243
rect 15281 25215 15315 25253
rect 15465 25211 15499 25249
rect 16385 25215 16419 25253
rect 16569 25211 16603 25249
rect 17489 25215 17523 25253
rect 17673 25243 17707 25249
rect 17673 25221 17708 25243
rect 17673 25211 17707 25221
rect 18777 25211 18811 25253
rect 19881 25211 19915 25253
rect 20157 25211 20191 25253
rect 4949 25049 5223 25211
rect 5409 25049 6511 25211
rect 6513 25049 7615 25211
rect 7617 25049 8719 25211
rect 8721 25049 9823 25211
rect 9827 25037 9913 25194
rect 10009 25049 10559 25211
rect 10561 25049 11663 25211
rect 11665 25049 12767 25211
rect 12769 25049 13871 25211
rect 13873 25049 14975 25211
rect 14979 25037 15065 25194
rect 15161 25049 15527 25211
rect 15529 25049 16631 25211
rect 16633 25049 17735 25211
rect 17737 25049 18839 25211
rect 18841 25049 19943 25211
rect 19945 25049 20219 25211
rect 4949 24165 5223 24327
rect 5409 24165 6143 24327
rect 6145 24165 7247 24327
rect 7251 24182 7337 24339
rect 7433 24165 7983 24327
rect 7985 24165 9087 24327
rect 9089 24165 10191 24327
rect 10193 24165 11295 24327
rect 11297 24165 12399 24327
rect 12403 24182 12489 24339
rect 12585 24165 13135 24327
rect 13137 24165 14239 24327
rect 14241 24165 15343 24327
rect 15345 24165 16447 24327
rect 16449 24165 17551 24327
rect 17555 24182 17641 24339
rect 17737 24165 18839 24327
rect 18841 24165 19943 24327
rect 19945 24165 20219 24327
rect 4977 24123 5011 24165
rect 5345 24132 5377 24156
rect 6081 24127 6115 24165
rect 6449 24123 6483 24161
rect 7185 24127 7219 24165
rect 7380 24133 7404 24155
rect 7553 24123 7587 24161
rect 7921 24127 7955 24165
rect 8657 24123 8691 24161
rect 9025 24127 9059 24165
rect 9761 24123 9795 24161
rect 9956 24133 9980 24155
rect 10129 24127 10163 24165
rect 10497 24123 10531 24161
rect 11233 24127 11267 24165
rect 11601 24123 11635 24161
rect 12337 24127 12371 24165
rect 12532 24133 12556 24155
rect 12705 24123 12739 24161
rect 13073 24127 13107 24165
rect 13809 24123 13843 24161
rect 14177 24127 14211 24165
rect 14913 24123 14947 24161
rect 15108 24133 15132 24155
rect 15281 24127 15315 24165
rect 15465 24123 15499 24161
rect 16385 24127 16419 24165
rect 16569 24123 16603 24161
rect 17489 24127 17523 24165
rect 17673 24155 17707 24161
rect 17673 24133 17708 24155
rect 17673 24123 17707 24133
rect 18777 24123 18811 24165
rect 19881 24123 19915 24165
rect 20157 24123 20191 24165
rect 4949 23961 5223 24123
rect 5409 23961 6511 24123
rect 6513 23961 7615 24123
rect 7617 23961 8719 24123
rect 8721 23961 9823 24123
rect 9827 23949 9913 24106
rect 10009 23961 10559 24123
rect 10561 23961 11663 24123
rect 11665 23961 12767 24123
rect 12769 23961 13871 24123
rect 13873 23961 14975 24123
rect 14979 23949 15065 24106
rect 15161 23961 15527 24123
rect 15529 23961 16631 24123
rect 16633 23961 17735 24123
rect 17737 23961 18839 24123
rect 18841 23961 19943 24123
rect 19945 23961 20219 24123
rect 4949 23077 5223 23239
rect 5409 23077 6143 23239
rect 6145 23077 7247 23239
rect 7251 23094 7337 23251
rect 7433 23077 7983 23239
rect 7985 23077 9087 23239
rect 9089 23077 10191 23239
rect 10193 23077 11295 23239
rect 11297 23077 12399 23239
rect 12403 23094 12489 23251
rect 12585 23077 13135 23239
rect 13137 23077 14239 23239
rect 14241 23077 15343 23239
rect 15345 23077 16447 23239
rect 16449 23077 17551 23239
rect 17555 23094 17641 23251
rect 17737 23077 18839 23239
rect 18841 23077 19943 23239
rect 19945 23077 20219 23239
rect 4977 23035 5011 23077
rect 5345 23044 5377 23068
rect 6081 23039 6115 23077
rect 6449 23035 6483 23073
rect 7185 23039 7219 23077
rect 7380 23045 7404 23067
rect 7553 23035 7587 23073
rect 7921 23039 7955 23077
rect 8657 23035 8691 23073
rect 9025 23039 9059 23077
rect 9761 23035 9795 23073
rect 9956 23045 9980 23067
rect 10129 23039 10163 23077
rect 10497 23035 10531 23073
rect 11233 23039 11267 23077
rect 11601 23035 11635 23073
rect 12337 23039 12371 23077
rect 12532 23045 12556 23067
rect 12705 23035 12739 23073
rect 13073 23039 13107 23077
rect 13809 23035 13843 23073
rect 14177 23039 14211 23077
rect 14913 23035 14947 23073
rect 15108 23045 15132 23067
rect 15281 23039 15315 23077
rect 15465 23035 15499 23073
rect 16385 23039 16419 23077
rect 16569 23035 16603 23073
rect 17489 23039 17523 23077
rect 17673 23067 17707 23073
rect 17673 23045 17708 23067
rect 17673 23035 17707 23045
rect 18777 23035 18811 23077
rect 19881 23035 19915 23077
rect 20157 23035 20191 23077
rect 4949 22873 5223 23035
rect 5409 22873 6511 23035
rect 6513 22873 7615 23035
rect 7617 22873 8719 23035
rect 8721 22873 9823 23035
rect 9827 22861 9913 23018
rect 10009 22873 10559 23035
rect 10561 22873 11663 23035
rect 11665 22873 12767 23035
rect 12769 22873 13871 23035
rect 13873 22873 14975 23035
rect 14979 22861 15065 23018
rect 15161 22873 15527 23035
rect 15529 22873 16631 23035
rect 16633 22873 17735 23035
rect 17737 22873 18839 23035
rect 18841 22873 19943 23035
rect 19945 22873 20219 23035
rect 4949 21989 5223 22151
rect 5409 21989 6143 22151
rect 6145 21989 7247 22151
rect 7251 22006 7337 22163
rect 7433 21989 7983 22151
rect 7985 21989 9087 22151
rect 9089 21989 10191 22151
rect 10193 21989 11295 22151
rect 11297 21989 12399 22151
rect 12403 22006 12489 22163
rect 12585 21989 13135 22151
rect 13137 21989 14239 22151
rect 14241 21989 15343 22151
rect 15345 21989 16447 22151
rect 16449 21989 17551 22151
rect 17555 22006 17641 22163
rect 17737 21989 18839 22151
rect 18841 21989 19943 22151
rect 19945 21989 20219 22151
rect 4977 21947 5011 21989
rect 5345 21956 5377 21980
rect 6081 21951 6115 21989
rect 6449 21947 6483 21985
rect 7185 21951 7219 21989
rect 7380 21957 7404 21979
rect 7553 21947 7587 21985
rect 7921 21951 7955 21989
rect 8657 21947 8691 21985
rect 9025 21951 9059 21989
rect 9761 21947 9795 21985
rect 9956 21957 9980 21979
rect 10129 21951 10163 21989
rect 10497 21947 10531 21985
rect 11233 21951 11267 21989
rect 11601 21947 11635 21985
rect 12337 21951 12371 21989
rect 12532 21957 12556 21979
rect 12705 21947 12739 21985
rect 13073 21951 13107 21989
rect 13809 21947 13843 21985
rect 14177 21951 14211 21989
rect 14913 21947 14947 21985
rect 15108 21957 15132 21979
rect 15281 21951 15315 21989
rect 15465 21947 15499 21985
rect 16385 21951 16419 21989
rect 16569 21947 16603 21985
rect 17489 21951 17523 21989
rect 17673 21979 17707 21985
rect 17673 21957 17708 21979
rect 17673 21947 17707 21957
rect 18777 21947 18811 21989
rect 19881 21947 19915 21989
rect 20157 21947 20191 21989
rect 4949 21785 5223 21947
rect 5409 21785 6511 21947
rect 6513 21785 7615 21947
rect 7617 21785 8719 21947
rect 8721 21785 9823 21947
rect 9827 21773 9913 21930
rect 10009 21785 10559 21947
rect 10561 21785 11663 21947
rect 11665 21785 12767 21947
rect 12769 21785 13871 21947
rect 13873 21785 14975 21947
rect 14979 21773 15065 21930
rect 15161 21785 15527 21947
rect 15529 21785 16631 21947
rect 16633 21785 17735 21947
rect 17737 21785 18839 21947
rect 18841 21785 19943 21947
rect 19945 21785 20219 21947
rect 4949 20901 5223 21063
rect 5409 20901 6143 21063
rect 6145 20901 7247 21063
rect 7251 20918 7337 21075
rect 7433 20901 7983 21063
rect 7985 20901 9087 21063
rect 9089 20901 10191 21063
rect 10193 20901 11295 21063
rect 11297 20901 12399 21063
rect 12403 20918 12489 21075
rect 12585 20901 13135 21063
rect 13137 20901 14239 21063
rect 14241 20901 15343 21063
rect 15345 20901 16447 21063
rect 16449 20901 17551 21063
rect 17555 20918 17641 21075
rect 17737 20901 18839 21063
rect 18841 20901 19943 21063
rect 19945 20901 20219 21063
rect 4977 20859 5011 20901
rect 5345 20868 5377 20892
rect 6081 20863 6115 20901
rect 6449 20859 6483 20897
rect 7185 20863 7219 20901
rect 7380 20869 7404 20891
rect 7553 20859 7587 20897
rect 7921 20863 7955 20901
rect 8657 20859 8691 20897
rect 9025 20863 9059 20901
rect 9761 20859 9795 20897
rect 9956 20869 9980 20891
rect 10129 20863 10163 20901
rect 10497 20859 10531 20897
rect 11233 20863 11267 20901
rect 11601 20859 11635 20897
rect 12337 20863 12371 20901
rect 12532 20869 12556 20891
rect 12705 20859 12739 20897
rect 13073 20863 13107 20901
rect 13809 20859 13843 20897
rect 14177 20863 14211 20901
rect 14913 20859 14947 20897
rect 15108 20869 15132 20891
rect 15281 20863 15315 20901
rect 15465 20859 15499 20897
rect 16385 20863 16419 20901
rect 16569 20859 16603 20897
rect 17489 20863 17523 20901
rect 17673 20891 17707 20897
rect 17673 20869 17708 20891
rect 17673 20859 17707 20869
rect 18777 20859 18811 20901
rect 19881 20859 19915 20901
rect 20157 20859 20191 20901
rect 4949 20697 5223 20859
rect 5409 20697 6511 20859
rect 6513 20697 7615 20859
rect 7617 20697 8719 20859
rect 8721 20697 9823 20859
rect 9827 20685 9913 20842
rect 10009 20697 10559 20859
rect 10561 20697 11663 20859
rect 11665 20697 12767 20859
rect 12769 20697 13871 20859
rect 13873 20697 14975 20859
rect 14979 20685 15065 20842
rect 15161 20697 15527 20859
rect 15529 20697 16631 20859
rect 16633 20697 17735 20859
rect 17737 20697 18839 20859
rect 18841 20697 19943 20859
rect 19945 20697 20219 20859
rect 4949 19813 5223 19975
rect 5409 19813 6143 19975
rect 6145 19813 7247 19975
rect 7251 19830 7337 19987
rect 7433 19813 7983 19975
rect 7985 19813 9087 19975
rect 9089 19813 10191 19975
rect 10193 19813 11295 19975
rect 11297 19813 12399 19975
rect 12403 19830 12489 19987
rect 12585 19813 13135 19975
rect 13137 19813 14239 19975
rect 14241 19813 15343 19975
rect 15345 19813 16447 19975
rect 16449 19813 17551 19975
rect 17555 19830 17641 19987
rect 17737 19813 18839 19975
rect 18841 19813 19943 19975
rect 19945 19813 20219 19975
rect 4977 19771 5011 19813
rect 5345 19780 5377 19804
rect 6081 19775 6115 19813
rect 6449 19771 6483 19809
rect 7185 19775 7219 19813
rect 7380 19781 7404 19803
rect 7553 19771 7587 19809
rect 7921 19775 7955 19813
rect 8657 19771 8691 19809
rect 9025 19775 9059 19813
rect 9761 19771 9795 19809
rect 9956 19781 9980 19803
rect 10129 19775 10163 19813
rect 10497 19771 10531 19809
rect 11233 19775 11267 19813
rect 11601 19771 11635 19809
rect 12337 19775 12371 19813
rect 12532 19781 12556 19803
rect 12705 19771 12739 19809
rect 13073 19775 13107 19813
rect 13809 19771 13843 19809
rect 14177 19775 14211 19813
rect 14913 19771 14947 19809
rect 15108 19781 15132 19803
rect 15281 19775 15315 19813
rect 15465 19771 15499 19809
rect 16385 19775 16419 19813
rect 16569 19771 16603 19809
rect 17489 19775 17523 19813
rect 17673 19803 17707 19809
rect 17673 19781 17708 19803
rect 17673 19771 17707 19781
rect 18777 19771 18811 19813
rect 19881 19771 19915 19813
rect 20157 19771 20191 19813
rect 4949 19609 5223 19771
rect 5409 19609 6511 19771
rect 6513 19609 7615 19771
rect 7617 19609 8719 19771
rect 8721 19609 9823 19771
rect 9827 19597 9913 19754
rect 10009 19609 10559 19771
rect 10561 19609 11663 19771
rect 11665 19609 12767 19771
rect 12769 19609 13871 19771
rect 13873 19609 14975 19771
rect 14979 19597 15065 19754
rect 15161 19609 15527 19771
rect 15529 19609 16631 19771
rect 16633 19609 17735 19771
rect 17737 19609 18839 19771
rect 18841 19609 19943 19771
rect 19945 19609 20219 19771
rect 4949 18725 5223 18887
rect 5409 18725 6143 18887
rect 6145 18725 7247 18887
rect 7251 18742 7337 18899
rect 7433 18725 7983 18887
rect 7985 18725 9087 18887
rect 9089 18725 10191 18887
rect 10193 18725 11295 18887
rect 11297 18725 12399 18887
rect 12403 18742 12489 18899
rect 12585 18725 13135 18887
rect 13137 18725 14239 18887
rect 14241 18725 15343 18887
rect 15345 18725 16447 18887
rect 16449 18725 17551 18887
rect 17555 18742 17641 18899
rect 17737 18725 18839 18887
rect 18841 18725 19943 18887
rect 19945 18725 20219 18887
rect 4977 18683 5011 18725
rect 5345 18692 5377 18716
rect 6081 18687 6115 18725
rect 6449 18683 6483 18721
rect 7185 18687 7219 18725
rect 7380 18693 7404 18715
rect 7553 18683 7587 18721
rect 7921 18687 7955 18725
rect 8657 18683 8691 18721
rect 9025 18687 9059 18725
rect 9761 18683 9795 18721
rect 9956 18693 9980 18715
rect 10129 18687 10163 18725
rect 10497 18683 10531 18721
rect 11233 18687 11267 18725
rect 11601 18683 11635 18721
rect 12337 18687 12371 18725
rect 12532 18693 12556 18715
rect 12705 18683 12739 18721
rect 13073 18687 13107 18725
rect 13809 18683 13843 18721
rect 14177 18687 14211 18725
rect 14913 18683 14947 18721
rect 15108 18693 15132 18715
rect 15281 18687 15315 18725
rect 15465 18683 15499 18721
rect 16385 18687 16419 18725
rect 16569 18683 16603 18721
rect 17489 18687 17523 18725
rect 17673 18715 17707 18721
rect 17673 18693 17708 18715
rect 17673 18683 17707 18693
rect 18777 18683 18811 18725
rect 19881 18683 19915 18725
rect 20157 18683 20191 18725
rect 4949 18521 5223 18683
rect 5409 18521 6511 18683
rect 6513 18521 7615 18683
rect 7617 18521 8719 18683
rect 8721 18521 9823 18683
rect 9827 18509 9913 18666
rect 10009 18521 10559 18683
rect 10561 18521 11663 18683
rect 11665 18521 12767 18683
rect 12769 18521 13871 18683
rect 13873 18521 14975 18683
rect 14979 18509 15065 18666
rect 15161 18521 15527 18683
rect 15529 18521 16631 18683
rect 16633 18521 17735 18683
rect 17737 18521 18839 18683
rect 18841 18521 19943 18683
rect 19945 18521 20219 18683
rect 4949 17637 5223 17799
rect 5409 17637 6143 17799
rect 6145 17637 7247 17799
rect 7251 17654 7337 17811
rect 7433 17637 7983 17799
rect 7985 17637 9087 17799
rect 9089 17637 10191 17799
rect 10193 17637 11295 17799
rect 11297 17637 12399 17799
rect 12403 17654 12489 17811
rect 12585 17637 13135 17799
rect 13137 17637 14239 17799
rect 14241 17637 15343 17799
rect 15345 17637 16447 17799
rect 16449 17637 17551 17799
rect 17555 17654 17641 17811
rect 17737 17637 18839 17799
rect 18841 17637 19943 17799
rect 19945 17637 20219 17799
rect 4977 17595 5011 17637
rect 5345 17604 5377 17628
rect 6081 17599 6115 17637
rect 6449 17595 6483 17633
rect 7185 17599 7219 17637
rect 7380 17605 7404 17627
rect 7553 17595 7587 17633
rect 7921 17599 7955 17637
rect 8657 17595 8691 17633
rect 9025 17599 9059 17637
rect 9761 17595 9795 17633
rect 9956 17605 9980 17627
rect 10129 17599 10163 17637
rect 10497 17595 10531 17633
rect 11233 17599 11267 17637
rect 11601 17595 11635 17633
rect 12337 17599 12371 17637
rect 12532 17605 12556 17627
rect 12705 17595 12739 17633
rect 13073 17599 13107 17637
rect 13809 17595 13843 17633
rect 14177 17599 14211 17637
rect 14913 17595 14947 17633
rect 15108 17605 15132 17627
rect 15281 17599 15315 17637
rect 15465 17595 15499 17633
rect 16385 17599 16419 17637
rect 16569 17595 16603 17633
rect 17489 17599 17523 17637
rect 17673 17627 17707 17633
rect 17673 17605 17708 17627
rect 17673 17595 17707 17605
rect 18777 17595 18811 17637
rect 19881 17595 19915 17637
rect 20157 17595 20191 17637
rect 4949 17433 5223 17595
rect 5409 17433 6511 17595
rect 6513 17433 7615 17595
rect 7617 17433 8719 17595
rect 8721 17433 9823 17595
rect 9827 17421 9913 17578
rect 10009 17433 10559 17595
rect 10561 17433 11663 17595
rect 11665 17433 12767 17595
rect 12769 17433 13871 17595
rect 13873 17433 14975 17595
rect 14979 17421 15065 17578
rect 15161 17433 15527 17595
rect 15529 17433 16631 17595
rect 16633 17433 17735 17595
rect 17737 17433 18839 17595
rect 18841 17433 19943 17595
rect 19945 17433 20219 17595
rect 4949 16549 5223 16711
rect 5409 16549 6143 16711
rect 6145 16549 7247 16711
rect 7251 16566 7337 16723
rect 7433 16549 7983 16711
rect 7985 16549 9087 16711
rect 9089 16549 10191 16711
rect 10193 16549 11295 16711
rect 11297 16549 12399 16711
rect 12403 16566 12489 16723
rect 12585 16549 13135 16711
rect 13137 16549 14239 16711
rect 14241 16549 15343 16711
rect 15345 16549 16447 16711
rect 16449 16549 17551 16711
rect 17555 16566 17641 16723
rect 17737 16549 18839 16711
rect 18841 16549 19943 16711
rect 19945 16549 20219 16711
rect 4977 16507 5011 16549
rect 5345 16516 5377 16540
rect 6081 16511 6115 16549
rect 6449 16507 6483 16545
rect 7185 16511 7219 16549
rect 7380 16517 7404 16539
rect 7553 16507 7587 16545
rect 7921 16511 7955 16549
rect 8657 16507 8691 16545
rect 9025 16511 9059 16549
rect 9761 16507 9795 16545
rect 9956 16517 9980 16539
rect 10129 16511 10163 16549
rect 10497 16507 10531 16545
rect 11233 16511 11267 16549
rect 11601 16507 11635 16545
rect 12337 16511 12371 16549
rect 12532 16517 12556 16539
rect 12705 16507 12739 16545
rect 13073 16511 13107 16549
rect 13809 16507 13843 16545
rect 14177 16511 14211 16549
rect 14913 16507 14947 16545
rect 15108 16517 15132 16539
rect 15281 16511 15315 16549
rect 15465 16507 15499 16545
rect 16385 16511 16419 16549
rect 16569 16507 16603 16545
rect 17489 16511 17523 16549
rect 17673 16539 17707 16545
rect 17673 16517 17708 16539
rect 17673 16507 17707 16517
rect 18777 16507 18811 16549
rect 19881 16507 19915 16549
rect 20157 16507 20191 16549
rect 4949 16345 5223 16507
rect 5409 16345 6511 16507
rect 6513 16345 7615 16507
rect 7617 16345 8719 16507
rect 8721 16345 9823 16507
rect 9827 16333 9913 16490
rect 10009 16345 10559 16507
rect 10561 16345 11663 16507
rect 11665 16345 12767 16507
rect 12769 16345 13871 16507
rect 13873 16345 14975 16507
rect 14979 16333 15065 16490
rect 15161 16345 15527 16507
rect 15529 16345 16631 16507
rect 16633 16345 17735 16507
rect 17737 16345 18839 16507
rect 18841 16345 19943 16507
rect 19945 16345 20219 16507
rect 4949 15461 5223 15623
rect 5409 15461 6143 15623
rect 6145 15461 7247 15623
rect 7251 15478 7337 15635
rect 7433 15461 7983 15623
rect 7985 15461 9087 15623
rect 9089 15461 10191 15623
rect 10193 15461 11295 15623
rect 11297 15461 12399 15623
rect 12403 15478 12489 15635
rect 12585 15461 13135 15623
rect 13137 15461 14239 15623
rect 14241 15461 15343 15623
rect 15345 15461 16447 15623
rect 16449 15461 17551 15623
rect 17555 15478 17641 15635
rect 17737 15461 18839 15623
rect 18841 15461 19943 15623
rect 19945 15461 20219 15623
rect 4977 15419 5011 15461
rect 5345 15428 5377 15452
rect 6081 15423 6115 15461
rect 6449 15419 6483 15457
rect 7185 15423 7219 15461
rect 7380 15429 7404 15451
rect 7553 15419 7587 15457
rect 7921 15423 7955 15461
rect 8657 15419 8691 15457
rect 9025 15423 9059 15461
rect 9761 15419 9795 15457
rect 9956 15429 9980 15451
rect 10129 15423 10163 15461
rect 10497 15419 10531 15457
rect 11233 15423 11267 15461
rect 11601 15419 11635 15457
rect 12337 15423 12371 15461
rect 12532 15429 12556 15451
rect 12705 15419 12739 15457
rect 12797 15419 12831 15457
rect 13073 15423 13107 15461
rect 13809 15419 13843 15457
rect 14177 15423 14211 15461
rect 14913 15419 14947 15457
rect 15281 15419 15315 15461
rect 15373 15419 15407 15457
rect 16385 15423 16419 15461
rect 16569 15419 16603 15457
rect 17489 15423 17523 15461
rect 17673 15451 17707 15457
rect 17673 15429 17708 15451
rect 17673 15419 17707 15429
rect 18777 15419 18811 15461
rect 19881 15419 19915 15461
rect 20157 15419 20191 15461
rect 4949 15257 5223 15419
rect 5409 15257 6511 15419
rect 6513 15257 7615 15419
rect 7617 15257 8719 15419
rect 8721 15257 9823 15419
rect 9827 15245 9913 15402
rect 10009 15257 10559 15419
rect 10561 15257 11663 15419
rect 11665 15257 12767 15419
rect 12791 15283 13484 15419
rect 13300 15237 13484 15283
rect 13505 15257 13871 15419
rect 13873 15257 14975 15419
rect 14979 15245 15065 15402
rect 15069 15257 15343 15419
rect 15367 15283 16060 15419
rect 15876 15237 16060 15283
rect 16081 15257 16631 15419
rect 16633 15257 17735 15419
rect 17737 15257 18839 15419
rect 18841 15257 19943 15419
rect 19945 15257 20219 15419
rect 4949 14373 5223 14535
rect 5409 14373 6143 14535
rect 6145 14373 7247 14535
rect 7251 14390 7337 14547
rect 7341 14373 8443 14535
rect 8445 14373 9547 14535
rect 9549 14373 10651 14535
rect 11293 14509 11479 14555
rect 10699 14373 11479 14509
rect 11665 14373 12399 14535
rect 12403 14390 12489 14547
rect 13317 14509 13503 14555
rect 12723 14373 13503 14509
rect 13505 14373 14239 14535
rect 14241 14373 14515 14529
rect 14517 14509 14701 14555
rect 15267 14509 15453 14553
rect 14517 14373 16355 14509
rect 16449 14373 17551 14535
rect 17555 14390 17641 14547
rect 17737 14373 18839 14535
rect 18841 14373 19943 14535
rect 19945 14373 20219 14535
rect 4977 14331 5011 14373
rect 5345 14340 5377 14364
rect 6081 14335 6115 14373
rect 6449 14331 6483 14369
rect 7185 14335 7219 14373
rect 7553 14331 7587 14369
rect 8381 14335 8415 14373
rect 8657 14331 8691 14369
rect 9485 14335 9519 14373
rect 9761 14331 9795 14369
rect 10037 14340 10069 14362
rect 10589 14335 10623 14373
rect 11362 14335 11396 14373
rect 11601 14342 11633 14364
rect 11877 14331 11911 14369
rect 12153 14331 12187 14369
rect 12337 14335 12371 14373
rect 12613 14342 12645 14364
rect 13386 14335 13420 14373
rect 13993 14331 14027 14369
rect 14177 14335 14211 14373
rect 14269 14331 14303 14373
rect 15108 14341 15132 14363
rect 15244 14331 15278 14369
rect 16201 14331 16235 14369
rect 16293 14335 16327 14373
rect 16396 14341 16420 14363
rect 16477 14331 16511 14369
rect 16580 14341 16604 14363
rect 17489 14335 17523 14373
rect 17673 14363 17707 14369
rect 17673 14341 17708 14363
rect 17673 14331 17707 14341
rect 18777 14331 18811 14373
rect 19881 14331 19915 14373
rect 20157 14331 20191 14373
rect 4949 14169 5223 14331
rect 5409 14169 6511 14331
rect 6513 14169 7615 14331
rect 7617 14169 8719 14331
rect 8721 14169 9823 14331
rect 9827 14157 9913 14314
rect 10101 14195 11939 14331
rect 10101 14149 10285 14195
rect 10851 14151 11037 14195
rect 11941 14175 12215 14331
rect 12234 14195 14055 14331
rect 14263 14195 14956 14331
rect 14772 14149 14956 14195
rect 14979 14157 15065 14314
rect 15161 14195 15941 14331
rect 15161 14149 15347 14195
rect 15989 14175 16263 14331
rect 16265 14175 16539 14331
rect 16633 14169 17735 14331
rect 17737 14169 18839 14331
rect 18841 14169 19943 14331
rect 19945 14169 20219 14331
rect 4949 13285 5223 13447
rect 5409 13285 6143 13447
rect 6145 13285 7247 13447
rect 7251 13302 7337 13459
rect 7433 13285 8535 13447
rect 8537 13285 9639 13447
rect 9641 13285 9915 13441
rect 9934 13285 11755 13421
rect 11849 13285 12399 13447
rect 12403 13302 12489 13459
rect 12493 13285 12767 13441
rect 12861 13421 13045 13467
rect 13611 13421 13797 13465
rect 16541 13421 16727 13467
rect 12861 13285 14699 13421
rect 14701 13285 16522 13421
rect 16541 13285 17321 13421
rect 17555 13302 17641 13459
rect 17737 13285 18839 13447
rect 18841 13285 19943 13447
rect 19945 13285 20219 13447
rect 4977 13243 5011 13285
rect 5345 13254 5377 13276
rect 5713 13243 5747 13281
rect 6081 13247 6115 13285
rect 6817 13243 6851 13281
rect 7185 13247 7219 13285
rect 7380 13253 7404 13275
rect 7921 13243 7955 13281
rect 8473 13247 8507 13285
rect 9025 13243 9059 13281
rect 9117 13243 9151 13281
rect 9577 13247 9611 13285
rect 9669 13247 9703 13285
rect 9956 13253 9980 13275
rect 10313 13243 10347 13281
rect 11693 13247 11727 13285
rect 11796 13253 11820 13275
rect 12153 13243 12187 13281
rect 12245 13243 12279 13281
rect 12337 13247 12371 13285
rect 12705 13247 12739 13285
rect 12808 13253 12832 13275
rect 14140 13243 14174 13281
rect 14637 13247 14671 13285
rect 14729 13247 14763 13285
rect 14924 13253 14948 13275
rect 16624 13247 16658 13285
rect 16845 13243 16879 13281
rect 17489 13254 17521 13276
rect 17581 13243 17615 13281
rect 17684 13253 17708 13275
rect 18777 13243 18811 13285
rect 19881 13243 19915 13285
rect 20157 13243 20191 13285
rect 4949 13081 5223 13243
rect 5225 13081 5775 13243
rect 5777 13081 6879 13243
rect 6881 13081 7983 13243
rect 7985 13081 9087 13243
rect 9111 13107 9804 13243
rect 9620 13061 9804 13107
rect 9827 13069 9913 13226
rect 10009 13081 10375 13243
rect 10377 13107 12215 13243
rect 12217 13107 14055 13243
rect 10377 13061 10561 13107
rect 11127 13063 11313 13107
rect 13119 13063 13305 13107
rect 13871 13061 14055 13107
rect 14057 13107 14837 13243
rect 14057 13061 14243 13107
rect 14979 13069 15065 13226
rect 15069 13107 16907 13243
rect 16928 13107 17621 13243
rect 15069 13061 15253 13107
rect 15819 13063 16005 13107
rect 16928 13061 17112 13107
rect 17737 13081 18839 13243
rect 18841 13081 19943 13243
rect 19945 13081 20219 13243
rect 4949 12197 5223 12359
rect 5593 12197 6695 12359
rect 6699 12197 7247 12333
rect 7251 12214 7337 12371
rect 7341 12197 7707 12359
rect 7709 12197 8811 12359
rect 8815 12197 9363 12333
rect 9457 12197 9823 12359
rect 9827 12214 9913 12371
rect 10469 12333 10655 12379
rect 12029 12333 12215 12379
rect 9919 12197 10467 12333
rect 10469 12197 11249 12333
rect 11435 12197 12215 12333
rect 12403 12214 12489 12371
rect 12679 12197 13227 12333
rect 13229 12197 13777 12333
rect 13781 12197 14055 12353
rect 14588 12333 14772 12379
rect 14079 12197 14772 12333
rect 14979 12214 15065 12371
rect 15971 12333 16157 12377
rect 16723 12333 16907 12379
rect 15069 12197 16907 12333
rect 17001 12197 17549 12333
rect 17555 12214 17641 12371
rect 17737 12197 18287 12359
rect 18289 12197 19391 12359
rect 19393 12197 19941 12333
rect 19945 12197 20219 12359
rect 4977 12159 5011 12197
rect 5437 12159 5471 12193
rect 5540 12165 5564 12187
rect 6633 12159 6667 12197
rect 7185 12159 7219 12197
rect 7645 12159 7679 12197
rect 8749 12159 8783 12197
rect 9301 12159 9335 12197
rect 9404 12165 9428 12187
rect 9761 12159 9795 12197
rect 10405 12159 10439 12197
rect 10552 12159 10586 12197
rect 11336 12165 11360 12187
rect 12098 12159 12132 12197
rect 12337 12166 12369 12188
rect 12613 12166 12645 12188
rect 13165 12159 13199 12197
rect 13257 12159 13291 12197
rect 13809 12159 13843 12197
rect 14085 12159 14119 12197
rect 14913 12166 14945 12188
rect 15097 12159 15131 12197
rect 16948 12165 16972 12187
rect 17029 12159 17063 12197
rect 17684 12165 17708 12187
rect 18225 12159 18259 12197
rect 19329 12159 19363 12197
rect 19421 12159 19455 12197
rect 20157 12159 20191 12197
rect 25680 6980 28308 9260
rect 3350 4640 3752 6036
rect 6650 4640 7052 5940
rect 9950 4640 10352 6080
rect 13250 4640 13652 6360
rect 16850 4640 17252 6920
rect 20050 4640 20770 6920
rect 23150 4640 24506 6920
rect 25650 4640 28278 6920
rect 29520 3930 34880 4860
rect 1250 1440 3430 2960
rect 4550 1440 6730 2960
rect 7850 1440 10030 2960
rect 11150 1440 13330 2960
rect 14750 1440 16930 2960
rect 18250 1440 20430 2960
rect 21950 1440 24130 2960
rect 25750 1440 27930 2960
<< nmos >>
rect 29918 4358 30118 4558
rect 30298 4358 30498 4558
rect 30698 4358 30898 4558
rect 31078 4358 31278 4558
rect 31336 4358 31536 4558
rect 31594 4358 31794 4558
rect 31852 4358 32052 4558
rect 32110 4358 32310 4558
rect 32368 4358 32568 4558
rect 32626 4358 32826 4558
rect 32884 4358 33084 4558
rect 33142 4358 33342 4558
rect 33518 4358 33718 4558
rect 1488 1708 1518 2708
rect 1688 2508 1718 2708
rect 1905 1701 1935 2701
rect 2001 1701 2031 2701
rect 2097 1701 2127 2701
rect 2193 1701 2223 2701
rect 2289 1701 2319 2701
rect 2385 1701 2415 2701
rect 2481 1701 2511 2701
rect 2577 1701 2607 2701
rect 2673 1701 2703 2701
rect 2769 1701 2799 2701
rect 2865 1701 2895 2701
rect 2961 1701 2991 2701
rect 3168 1708 3198 2708
rect 4788 1708 4818 2708
rect 4988 2508 5018 2708
rect 5205 1701 5235 2701
rect 5301 1701 5331 2701
rect 5397 1701 5427 2701
rect 5493 1701 5523 2701
rect 5589 1701 5619 2701
rect 5685 1701 5715 2701
rect 5781 1701 5811 2701
rect 5877 1701 5907 2701
rect 5973 1701 6003 2701
rect 6069 1701 6099 2701
rect 6165 1701 6195 2701
rect 6261 1701 6291 2701
rect 6468 1708 6498 2708
rect 8088 1708 8118 2708
rect 8288 2508 8318 2708
rect 8505 1701 8535 2701
rect 8601 1701 8631 2701
rect 8697 1701 8727 2701
rect 8793 1701 8823 2701
rect 8889 1701 8919 2701
rect 8985 1701 9015 2701
rect 9081 1701 9111 2701
rect 9177 1701 9207 2701
rect 9273 1701 9303 2701
rect 9369 1701 9399 2701
rect 9465 1701 9495 2701
rect 9561 1701 9591 2701
rect 9768 1708 9798 2708
rect 11388 1708 11418 2708
rect 11588 2508 11618 2708
rect 11805 1701 11835 2701
rect 11901 1701 11931 2701
rect 11997 1701 12027 2701
rect 12093 1701 12123 2701
rect 12189 1701 12219 2701
rect 12285 1701 12315 2701
rect 12381 1701 12411 2701
rect 12477 1701 12507 2701
rect 12573 1701 12603 2701
rect 12669 1701 12699 2701
rect 12765 1701 12795 2701
rect 12861 1701 12891 2701
rect 13068 1708 13098 2708
rect 14988 1708 15018 2708
rect 15188 2508 15218 2708
rect 15405 1701 15435 2701
rect 15501 1701 15531 2701
rect 15597 1701 15627 2701
rect 15693 1701 15723 2701
rect 15789 1701 15819 2701
rect 15885 1701 15915 2701
rect 15981 1701 16011 2701
rect 16077 1701 16107 2701
rect 16173 1701 16203 2701
rect 16269 1701 16299 2701
rect 16365 1701 16395 2701
rect 16461 1701 16491 2701
rect 16668 1708 16698 2708
rect 18488 1708 18518 2708
rect 18688 2508 18718 2708
rect 18905 1701 18935 2701
rect 19001 1701 19031 2701
rect 19097 1701 19127 2701
rect 19193 1701 19223 2701
rect 19289 1701 19319 2701
rect 19385 1701 19415 2701
rect 19481 1701 19511 2701
rect 19577 1701 19607 2701
rect 19673 1701 19703 2701
rect 19769 1701 19799 2701
rect 19865 1701 19895 2701
rect 19961 1701 19991 2701
rect 20168 1708 20198 2708
rect 22188 1708 22218 2708
rect 22388 2508 22418 2708
rect 22605 1701 22635 2701
rect 22701 1701 22731 2701
rect 22797 1701 22827 2701
rect 22893 1701 22923 2701
rect 22989 1701 23019 2701
rect 23085 1701 23115 2701
rect 23181 1701 23211 2701
rect 23277 1701 23307 2701
rect 23373 1701 23403 2701
rect 23469 1701 23499 2701
rect 23565 1701 23595 2701
rect 23661 1701 23691 2701
rect 23868 1708 23898 2708
rect 25988 1708 26018 2708
rect 26188 2508 26218 2708
rect 26405 1701 26435 2701
rect 26501 1701 26531 2701
rect 26597 1701 26627 2701
rect 26693 1701 26723 2701
rect 26789 1701 26819 2701
rect 26885 1701 26915 2701
rect 26981 1701 27011 2701
rect 27077 1701 27107 2701
rect 27173 1701 27203 2701
rect 27269 1701 27299 2701
rect 27365 1701 27395 2701
rect 27461 1701 27491 2701
rect 27668 1708 27698 2708
<< scnmos >>
rect 5027 27251 5145 27361
rect 5303 27251 5421 27361
rect 5587 27277 5617 27361
rect 5673 27277 5703 27361
rect 5759 27277 5789 27361
rect 5845 27277 5875 27361
rect 5942 27277 5972 27361
rect 6223 27251 7169 27361
rect 7419 27251 7537 27361
rect 7695 27251 8641 27361
rect 8799 27251 9745 27361
rect 10179 27257 10209 27361
rect 10267 27257 10297 27361
rect 10639 27251 11217 27361
rect 11375 27251 12321 27361
rect 12571 27251 12689 27361
rect 12847 27251 13793 27361
rect 13951 27251 14897 27361
rect 15147 27251 15265 27361
rect 15423 27251 16369 27361
rect 16527 27251 17473 27361
rect 17815 27251 18393 27361
rect 18559 27277 18589 27361
rect 18645 27277 18675 27361
rect 18731 27277 18761 27361
rect 18817 27277 18847 27361
rect 18914 27277 18944 27361
rect 19287 27251 19865 27361
rect 20023 27251 20141 27361
rect 5027 26367 5145 26477
rect 5487 26367 6065 26477
rect 6223 26367 7169 26477
rect 7511 26367 7905 26477
rect 8063 26367 9009 26477
rect 9167 26367 10113 26477
rect 10271 26367 11217 26477
rect 11375 26367 12321 26477
rect 12663 26367 13057 26477
rect 13215 26367 14161 26477
rect 14319 26367 15265 26477
rect 15423 26367 16369 26477
rect 16527 26367 17473 26477
rect 17815 26367 18761 26477
rect 18919 26367 19865 26477
rect 20023 26367 20141 26477
rect 5027 26163 5145 26273
rect 5487 26163 6433 26273
rect 6591 26163 7537 26273
rect 7695 26163 8641 26273
rect 8799 26163 9745 26273
rect 10087 26163 10481 26273
rect 10639 26163 11585 26273
rect 11743 26163 12689 26273
rect 12847 26163 13793 26273
rect 13951 26163 14897 26273
rect 15239 26163 15449 26273
rect 15607 26163 16553 26273
rect 16711 26163 17657 26273
rect 17815 26163 18761 26273
rect 18919 26163 19865 26273
rect 20023 26163 20141 26273
rect 5027 25279 5145 25389
rect 5487 25279 6065 25389
rect 6223 25279 7169 25389
rect 7511 25279 7905 25389
rect 8063 25279 9009 25389
rect 9167 25279 10113 25389
rect 10271 25279 11217 25389
rect 11375 25279 12321 25389
rect 12663 25279 13057 25389
rect 13215 25279 14161 25389
rect 14319 25279 15265 25389
rect 15423 25279 16369 25389
rect 16527 25279 17473 25389
rect 17815 25279 18761 25389
rect 18919 25279 19865 25389
rect 20023 25279 20141 25389
rect 5027 25075 5145 25185
rect 5487 25075 6433 25185
rect 6591 25075 7537 25185
rect 7695 25075 8641 25185
rect 8799 25075 9745 25185
rect 10087 25075 10481 25185
rect 10639 25075 11585 25185
rect 11743 25075 12689 25185
rect 12847 25075 13793 25185
rect 13951 25075 14897 25185
rect 15239 25075 15449 25185
rect 15607 25075 16553 25185
rect 16711 25075 17657 25185
rect 17815 25075 18761 25185
rect 18919 25075 19865 25185
rect 20023 25075 20141 25185
rect 5027 24191 5145 24301
rect 5487 24191 6065 24301
rect 6223 24191 7169 24301
rect 7511 24191 7905 24301
rect 8063 24191 9009 24301
rect 9167 24191 10113 24301
rect 10271 24191 11217 24301
rect 11375 24191 12321 24301
rect 12663 24191 13057 24301
rect 13215 24191 14161 24301
rect 14319 24191 15265 24301
rect 15423 24191 16369 24301
rect 16527 24191 17473 24301
rect 17815 24191 18761 24301
rect 18919 24191 19865 24301
rect 20023 24191 20141 24301
rect 5027 23987 5145 24097
rect 5487 23987 6433 24097
rect 6591 23987 7537 24097
rect 7695 23987 8641 24097
rect 8799 23987 9745 24097
rect 10087 23987 10481 24097
rect 10639 23987 11585 24097
rect 11743 23987 12689 24097
rect 12847 23987 13793 24097
rect 13951 23987 14897 24097
rect 15239 23987 15449 24097
rect 15607 23987 16553 24097
rect 16711 23987 17657 24097
rect 17815 23987 18761 24097
rect 18919 23987 19865 24097
rect 20023 23987 20141 24097
rect 5027 23103 5145 23213
rect 5487 23103 6065 23213
rect 6223 23103 7169 23213
rect 7511 23103 7905 23213
rect 8063 23103 9009 23213
rect 9167 23103 10113 23213
rect 10271 23103 11217 23213
rect 11375 23103 12321 23213
rect 12663 23103 13057 23213
rect 13215 23103 14161 23213
rect 14319 23103 15265 23213
rect 15423 23103 16369 23213
rect 16527 23103 17473 23213
rect 17815 23103 18761 23213
rect 18919 23103 19865 23213
rect 20023 23103 20141 23213
rect 5027 22899 5145 23009
rect 5487 22899 6433 23009
rect 6591 22899 7537 23009
rect 7695 22899 8641 23009
rect 8799 22899 9745 23009
rect 10087 22899 10481 23009
rect 10639 22899 11585 23009
rect 11743 22899 12689 23009
rect 12847 22899 13793 23009
rect 13951 22899 14897 23009
rect 15239 22899 15449 23009
rect 15607 22899 16553 23009
rect 16711 22899 17657 23009
rect 17815 22899 18761 23009
rect 18919 22899 19865 23009
rect 20023 22899 20141 23009
rect 5027 22015 5145 22125
rect 5487 22015 6065 22125
rect 6223 22015 7169 22125
rect 7511 22015 7905 22125
rect 8063 22015 9009 22125
rect 9167 22015 10113 22125
rect 10271 22015 11217 22125
rect 11375 22015 12321 22125
rect 12663 22015 13057 22125
rect 13215 22015 14161 22125
rect 14319 22015 15265 22125
rect 15423 22015 16369 22125
rect 16527 22015 17473 22125
rect 17815 22015 18761 22125
rect 18919 22015 19865 22125
rect 20023 22015 20141 22125
rect 5027 21811 5145 21921
rect 5487 21811 6433 21921
rect 6591 21811 7537 21921
rect 7695 21811 8641 21921
rect 8799 21811 9745 21921
rect 10087 21811 10481 21921
rect 10639 21811 11585 21921
rect 11743 21811 12689 21921
rect 12847 21811 13793 21921
rect 13951 21811 14897 21921
rect 15239 21811 15449 21921
rect 15607 21811 16553 21921
rect 16711 21811 17657 21921
rect 17815 21811 18761 21921
rect 18919 21811 19865 21921
rect 20023 21811 20141 21921
rect 5027 20927 5145 21037
rect 5487 20927 6065 21037
rect 6223 20927 7169 21037
rect 7511 20927 7905 21037
rect 8063 20927 9009 21037
rect 9167 20927 10113 21037
rect 10271 20927 11217 21037
rect 11375 20927 12321 21037
rect 12663 20927 13057 21037
rect 13215 20927 14161 21037
rect 14319 20927 15265 21037
rect 15423 20927 16369 21037
rect 16527 20927 17473 21037
rect 17815 20927 18761 21037
rect 18919 20927 19865 21037
rect 20023 20927 20141 21037
rect 5027 20723 5145 20833
rect 5487 20723 6433 20833
rect 6591 20723 7537 20833
rect 7695 20723 8641 20833
rect 8799 20723 9745 20833
rect 10087 20723 10481 20833
rect 10639 20723 11585 20833
rect 11743 20723 12689 20833
rect 12847 20723 13793 20833
rect 13951 20723 14897 20833
rect 15239 20723 15449 20833
rect 15607 20723 16553 20833
rect 16711 20723 17657 20833
rect 17815 20723 18761 20833
rect 18919 20723 19865 20833
rect 20023 20723 20141 20833
rect 5027 19839 5145 19949
rect 5487 19839 6065 19949
rect 6223 19839 7169 19949
rect 7511 19839 7905 19949
rect 8063 19839 9009 19949
rect 9167 19839 10113 19949
rect 10271 19839 11217 19949
rect 11375 19839 12321 19949
rect 12663 19839 13057 19949
rect 13215 19839 14161 19949
rect 14319 19839 15265 19949
rect 15423 19839 16369 19949
rect 16527 19839 17473 19949
rect 17815 19839 18761 19949
rect 18919 19839 19865 19949
rect 20023 19839 20141 19949
rect 5027 19635 5145 19745
rect 5487 19635 6433 19745
rect 6591 19635 7537 19745
rect 7695 19635 8641 19745
rect 8799 19635 9745 19745
rect 10087 19635 10481 19745
rect 10639 19635 11585 19745
rect 11743 19635 12689 19745
rect 12847 19635 13793 19745
rect 13951 19635 14897 19745
rect 15239 19635 15449 19745
rect 15607 19635 16553 19745
rect 16711 19635 17657 19745
rect 17815 19635 18761 19745
rect 18919 19635 19865 19745
rect 20023 19635 20141 19745
rect 5027 18751 5145 18861
rect 5487 18751 6065 18861
rect 6223 18751 7169 18861
rect 7511 18751 7905 18861
rect 8063 18751 9009 18861
rect 9167 18751 10113 18861
rect 10271 18751 11217 18861
rect 11375 18751 12321 18861
rect 12663 18751 13057 18861
rect 13215 18751 14161 18861
rect 14319 18751 15265 18861
rect 15423 18751 16369 18861
rect 16527 18751 17473 18861
rect 17815 18751 18761 18861
rect 18919 18751 19865 18861
rect 20023 18751 20141 18861
rect 5027 18547 5145 18657
rect 5487 18547 6433 18657
rect 6591 18547 7537 18657
rect 7695 18547 8641 18657
rect 8799 18547 9745 18657
rect 10087 18547 10481 18657
rect 10639 18547 11585 18657
rect 11743 18547 12689 18657
rect 12847 18547 13793 18657
rect 13951 18547 14897 18657
rect 15239 18547 15449 18657
rect 15607 18547 16553 18657
rect 16711 18547 17657 18657
rect 17815 18547 18761 18657
rect 18919 18547 19865 18657
rect 20023 18547 20141 18657
rect 5027 17663 5145 17773
rect 5487 17663 6065 17773
rect 6223 17663 7169 17773
rect 7511 17663 7905 17773
rect 8063 17663 9009 17773
rect 9167 17663 10113 17773
rect 10271 17663 11217 17773
rect 11375 17663 12321 17773
rect 12663 17663 13057 17773
rect 13215 17663 14161 17773
rect 14319 17663 15265 17773
rect 15423 17663 16369 17773
rect 16527 17663 17473 17773
rect 17815 17663 18761 17773
rect 18919 17663 19865 17773
rect 20023 17663 20141 17773
rect 5027 17459 5145 17569
rect 5487 17459 6433 17569
rect 6591 17459 7537 17569
rect 7695 17459 8641 17569
rect 8799 17459 9745 17569
rect 10087 17459 10481 17569
rect 10639 17459 11585 17569
rect 11743 17459 12689 17569
rect 12847 17459 13793 17569
rect 13951 17459 14897 17569
rect 15239 17459 15449 17569
rect 15607 17459 16553 17569
rect 16711 17459 17657 17569
rect 17815 17459 18761 17569
rect 18919 17459 19865 17569
rect 20023 17459 20141 17569
rect 5027 16575 5145 16685
rect 5487 16575 6065 16685
rect 6223 16575 7169 16685
rect 7511 16575 7905 16685
rect 8063 16575 9009 16685
rect 9167 16575 10113 16685
rect 10271 16575 11217 16685
rect 11375 16575 12321 16685
rect 12663 16575 13057 16685
rect 13215 16575 14161 16685
rect 14319 16575 15265 16685
rect 15423 16575 16369 16685
rect 16527 16575 17473 16685
rect 17815 16575 18761 16685
rect 18919 16575 19865 16685
rect 20023 16575 20141 16685
rect 5027 16371 5145 16481
rect 5487 16371 6433 16481
rect 6591 16371 7537 16481
rect 7695 16371 8641 16481
rect 8799 16371 9745 16481
rect 10087 16371 10481 16481
rect 10639 16371 11585 16481
rect 11743 16371 12689 16481
rect 12847 16371 13793 16481
rect 13951 16371 14897 16481
rect 15239 16371 15449 16481
rect 15607 16371 16553 16481
rect 16711 16371 17657 16481
rect 17815 16371 18761 16481
rect 18919 16371 19865 16481
rect 20023 16371 20141 16481
rect 5027 15487 5145 15597
rect 5487 15487 6065 15597
rect 6223 15487 7169 15597
rect 7511 15487 7905 15597
rect 8063 15487 9009 15597
rect 9167 15487 10113 15597
rect 10271 15487 11217 15597
rect 11375 15487 12321 15597
rect 12663 15487 13057 15597
rect 13215 15487 14161 15597
rect 14319 15487 15265 15597
rect 15423 15487 16369 15597
rect 16527 15487 17473 15597
rect 17815 15487 18761 15597
rect 18919 15487 19865 15597
rect 20023 15487 20141 15597
rect 5027 15283 5145 15393
rect 5487 15283 6433 15393
rect 6591 15283 7537 15393
rect 7695 15283 8641 15393
rect 8799 15283 9745 15393
rect 10087 15283 10481 15393
rect 10639 15283 11585 15393
rect 11743 15283 12689 15393
rect 12869 15309 12899 15393
rect 12953 15309 13053 15393
rect 13211 15309 13311 15393
rect 13376 15263 13406 15393
rect 13583 15283 13793 15393
rect 13951 15283 14897 15393
rect 15147 15283 15265 15393
rect 15445 15309 15475 15393
rect 15529 15309 15629 15393
rect 15787 15309 15887 15393
rect 15952 15263 15982 15393
rect 16159 15283 16553 15393
rect 16711 15283 17657 15393
rect 17815 15283 18761 15393
rect 18919 15283 19865 15393
rect 20023 15283 20141 15393
rect 5027 14399 5145 14509
rect 5487 14399 6065 14509
rect 6223 14399 7169 14509
rect 7419 14399 8365 14509
rect 8523 14399 9469 14509
rect 9627 14399 10573 14509
rect 10777 14399 10807 14483
rect 10945 14399 10975 14483
rect 11041 14399 11071 14483
rect 11166 14399 11196 14483
rect 11262 14399 11292 14483
rect 11371 14399 11401 14529
rect 11743 14399 12321 14509
rect 12801 14399 12831 14483
rect 12969 14399 12999 14483
rect 13065 14399 13095 14483
rect 13190 14399 13220 14483
rect 13286 14399 13316 14483
rect 13395 14399 13425 14529
rect 13583 14399 14161 14509
rect 14319 14399 14349 14503
rect 14407 14399 14437 14503
rect 14595 14399 14625 14529
rect 14803 14399 14833 14483
rect 14894 14399 14924 14483
rect 15043 14399 15073 14483
rect 15139 14399 15169 14471
rect 15248 14399 15278 14471
rect 15347 14399 15377 14527
rect 15479 14399 15509 14483
rect 15551 14399 15581 14483
rect 15717 14399 15747 14471
rect 15813 14399 15843 14471
rect 15908 14399 15938 14483
rect 16163 14399 16193 14483
rect 16247 14399 16277 14483
rect 16527 14399 17473 14509
rect 17815 14399 18761 14509
rect 18919 14399 19865 14509
rect 20023 14399 20141 14509
rect 5027 14195 5145 14305
rect 5487 14195 6433 14305
rect 6591 14195 7537 14305
rect 7695 14195 8641 14305
rect 8799 14195 9745 14305
rect 10179 14175 10209 14305
rect 10387 14221 10417 14305
rect 10478 14221 10508 14305
rect 10627 14221 10657 14305
rect 10723 14233 10753 14305
rect 10832 14233 10862 14305
rect 10931 14177 10961 14305
rect 11063 14221 11093 14305
rect 11135 14221 11165 14305
rect 11301 14233 11331 14305
rect 11397 14233 11427 14305
rect 11492 14221 11522 14305
rect 11747 14221 11777 14305
rect 11831 14221 11861 14305
rect 12019 14201 12049 14305
rect 12107 14201 12137 14305
rect 12313 14221 12343 14305
rect 12399 14221 12429 14305
rect 12485 14221 12515 14305
rect 12571 14221 12601 14305
rect 12657 14221 12687 14305
rect 12743 14221 12773 14305
rect 12829 14221 12859 14305
rect 12915 14221 12945 14305
rect 13000 14221 13030 14305
rect 13086 14221 13116 14305
rect 13172 14221 13202 14305
rect 13258 14221 13288 14305
rect 13344 14221 13374 14305
rect 13430 14221 13460 14305
rect 13516 14221 13546 14305
rect 13602 14221 13632 14305
rect 13688 14221 13718 14305
rect 13774 14221 13804 14305
rect 13860 14221 13890 14305
rect 13946 14221 13976 14305
rect 14341 14221 14371 14305
rect 14425 14221 14525 14305
rect 14683 14221 14783 14305
rect 14848 14175 14878 14305
rect 15239 14175 15269 14305
rect 15348 14221 15378 14305
rect 15444 14221 15474 14305
rect 15569 14221 15599 14305
rect 15665 14221 15695 14305
rect 15833 14221 15863 14305
rect 16067 14201 16097 14305
rect 16155 14201 16185 14305
rect 16343 14201 16373 14305
rect 16431 14201 16461 14305
rect 16711 14195 17657 14305
rect 17815 14195 18761 14305
rect 18919 14195 19865 14305
rect 20023 14195 20141 14305
rect 5027 13311 5145 13421
rect 5487 13311 6065 13421
rect 6223 13311 7169 13421
rect 7511 13311 8457 13421
rect 8615 13311 9561 13421
rect 9719 13311 9749 13415
rect 9807 13311 9837 13415
rect 10013 13311 10043 13395
rect 10099 13311 10129 13395
rect 10185 13311 10215 13395
rect 10271 13311 10301 13395
rect 10357 13311 10387 13395
rect 10443 13311 10473 13395
rect 10529 13311 10559 13395
rect 10615 13311 10645 13395
rect 10700 13311 10730 13395
rect 10786 13311 10816 13395
rect 10872 13311 10902 13395
rect 10958 13311 10988 13395
rect 11044 13311 11074 13395
rect 11130 13311 11160 13395
rect 11216 13311 11246 13395
rect 11302 13311 11332 13395
rect 11388 13311 11418 13395
rect 11474 13311 11504 13395
rect 11560 13311 11590 13395
rect 11646 13311 11676 13395
rect 11927 13311 12321 13421
rect 12571 13311 12601 13415
rect 12659 13311 12689 13415
rect 12939 13311 12969 13441
rect 13147 13311 13177 13395
rect 13238 13311 13268 13395
rect 13387 13311 13417 13395
rect 13483 13311 13513 13383
rect 13592 13311 13622 13383
rect 13691 13311 13721 13439
rect 13823 13311 13853 13395
rect 13895 13311 13925 13395
rect 14061 13311 14091 13383
rect 14157 13311 14187 13383
rect 14252 13311 14282 13395
rect 14507 13311 14537 13395
rect 14591 13311 14621 13395
rect 14780 13311 14810 13395
rect 14866 13311 14896 13395
rect 14952 13311 14982 13395
rect 15038 13311 15068 13395
rect 15124 13311 15154 13395
rect 15210 13311 15240 13395
rect 15296 13311 15326 13395
rect 15382 13311 15412 13395
rect 15468 13311 15498 13395
rect 15554 13311 15584 13395
rect 15640 13311 15670 13395
rect 15726 13311 15756 13395
rect 15811 13311 15841 13395
rect 15897 13311 15927 13395
rect 15983 13311 16013 13395
rect 16069 13311 16099 13395
rect 16155 13311 16185 13395
rect 16241 13311 16271 13395
rect 16327 13311 16357 13395
rect 16413 13311 16443 13395
rect 16619 13311 16649 13441
rect 16728 13311 16758 13395
rect 16824 13311 16854 13395
rect 16949 13311 16979 13395
rect 17045 13311 17075 13395
rect 17213 13311 17243 13395
rect 17815 13311 18761 13421
rect 18919 13311 19865 13421
rect 20023 13311 20141 13421
rect 5027 13107 5145 13217
rect 5303 13107 5697 13217
rect 5855 13107 6801 13217
rect 6959 13107 7905 13217
rect 8063 13107 9009 13217
rect 9189 13133 9219 13217
rect 9273 13133 9373 13217
rect 9531 13133 9631 13217
rect 9696 13087 9726 13217
rect 10087 13107 10297 13217
rect 10455 13087 10485 13217
rect 10663 13133 10693 13217
rect 10754 13133 10784 13217
rect 10903 13133 10933 13217
rect 10999 13145 11029 13217
rect 11108 13145 11138 13217
rect 11207 13089 11237 13217
rect 11339 13133 11369 13217
rect 11411 13133 11441 13217
rect 11577 13145 11607 13217
rect 11673 13145 11703 13217
rect 11768 13133 11798 13217
rect 12023 13133 12053 13217
rect 12107 13133 12137 13217
rect 12295 13133 12325 13217
rect 12379 13133 12409 13217
rect 12634 13133 12664 13217
rect 12729 13145 12759 13217
rect 12825 13145 12855 13217
rect 12991 13133 13021 13217
rect 13063 13133 13093 13217
rect 13195 13089 13225 13217
rect 13294 13145 13324 13217
rect 13403 13145 13433 13217
rect 13499 13133 13529 13217
rect 13648 13133 13678 13217
rect 13739 13133 13769 13217
rect 13947 13087 13977 13217
rect 14135 13087 14165 13217
rect 14244 13133 14274 13217
rect 14340 13133 14370 13217
rect 14465 13133 14495 13217
rect 14561 13133 14591 13217
rect 14729 13133 14759 13217
rect 15147 13087 15177 13217
rect 15355 13133 15385 13217
rect 15446 13133 15476 13217
rect 15595 13133 15625 13217
rect 15691 13145 15721 13217
rect 15800 13145 15830 13217
rect 15899 13089 15929 13217
rect 16031 13133 16061 13217
rect 16103 13133 16133 13217
rect 16269 13145 16299 13217
rect 16365 13145 16395 13217
rect 16460 13133 16490 13217
rect 16715 13133 16745 13217
rect 16799 13133 16829 13217
rect 17006 13087 17036 13217
rect 17101 13133 17201 13217
rect 17359 13133 17459 13217
rect 17513 13133 17543 13217
rect 17815 13107 18761 13217
rect 18919 13107 19865 13217
rect 20023 13107 20141 13217
rect 5027 12223 5145 12333
rect 5671 12223 6617 12333
rect 6783 12223 6813 12307
rect 6869 12223 6899 12307
rect 6955 12223 6985 12307
rect 7041 12223 7071 12307
rect 7138 12223 7168 12307
rect 7419 12223 7629 12333
rect 7787 12223 8733 12333
rect 8899 12223 8929 12307
rect 8985 12223 9015 12307
rect 9071 12223 9101 12307
rect 9157 12223 9187 12307
rect 9254 12223 9284 12307
rect 9535 12223 9745 12333
rect 10003 12223 10033 12307
rect 10089 12223 10119 12307
rect 10175 12223 10205 12307
rect 10261 12223 10291 12307
rect 10358 12223 10388 12307
rect 10547 12223 10577 12353
rect 10656 12223 10686 12307
rect 10752 12223 10782 12307
rect 10877 12223 10907 12307
rect 10973 12223 11003 12307
rect 11141 12223 11171 12307
rect 11513 12223 11543 12307
rect 11681 12223 11711 12307
rect 11777 12223 11807 12307
rect 11902 12223 11932 12307
rect 11998 12223 12028 12307
rect 12107 12223 12137 12353
rect 12763 12223 12793 12307
rect 12849 12223 12879 12307
rect 12935 12223 12965 12307
rect 13021 12223 13051 12307
rect 13118 12223 13148 12307
rect 13308 12223 13338 12307
rect 13405 12223 13435 12307
rect 13491 12223 13521 12307
rect 13577 12223 13607 12307
rect 13663 12223 13693 12307
rect 13859 12223 13889 12327
rect 13947 12223 13977 12327
rect 14157 12223 14187 12307
rect 14241 12223 14341 12307
rect 14499 12223 14599 12307
rect 14664 12223 14694 12353
rect 15147 12223 15177 12307
rect 15231 12223 15261 12307
rect 15486 12223 15516 12307
rect 15581 12223 15611 12295
rect 15677 12223 15707 12295
rect 15843 12223 15873 12307
rect 15915 12223 15945 12307
rect 16047 12223 16077 12351
rect 16146 12223 16176 12295
rect 16255 12223 16285 12295
rect 16351 12223 16381 12307
rect 16500 12223 16530 12307
rect 16591 12223 16621 12307
rect 16799 12223 16829 12353
rect 17080 12223 17110 12307
rect 17177 12223 17207 12307
rect 17263 12223 17293 12307
rect 17349 12223 17379 12307
rect 17435 12223 17465 12307
rect 17815 12223 18209 12333
rect 18367 12223 19313 12333
rect 19472 12223 19502 12307
rect 19569 12223 19599 12307
rect 19655 12223 19685 12307
rect 19741 12223 19771 12307
rect 19827 12223 19857 12307
rect 20023 12223 20141 12333
<< pmos >>
rect 29814 6150 30014 6750
rect 30194 6150 30394 6750
rect 30452 6150 30652 6750
rect 30834 6150 31034 6750
rect 31092 6150 31292 6750
rect 31350 6150 31550 6750
rect 31734 6150 31934 6750
rect 31992 6150 32192 6750
rect 32250 6150 32450 6750
rect 32508 6150 32708 6750
rect 32766 6150 32966 6750
rect 33024 6150 33224 6750
rect 33282 6150 33482 6750
rect 33540 6150 33740 6750
rect 33798 6150 33998 6750
rect 34056 6150 34256 6750
rect 34434 6150 34634 6750
rect 30074 5130 30104 5730
rect 30298 5130 30328 5730
rect 30394 5130 30424 5730
rect 30490 5130 30520 5730
rect 30698 5130 30728 5730
rect 30794 5130 30824 5730
rect 30890 5130 30920 5730
rect 31094 5130 31124 5730
rect 1484 3230 1514 4230
rect 1684 3230 1714 3830
rect 1901 3223 1931 4223
rect 1997 3223 2027 4223
rect 2093 3223 2123 4223
rect 2189 3223 2219 4223
rect 2285 3223 2315 4223
rect 2381 3223 2411 4223
rect 2477 3223 2507 4223
rect 2573 3223 2603 4223
rect 2669 3223 2699 4223
rect 2765 3223 2795 4223
rect 2861 3223 2891 4223
rect 2957 3223 2987 4223
rect 3184 3230 3214 4230
rect 4784 3230 4814 4230
rect 4984 3230 5014 3830
rect 5201 3223 5231 4223
rect 5297 3223 5327 4223
rect 5393 3223 5423 4223
rect 5489 3223 5519 4223
rect 5585 3223 5615 4223
rect 5681 3223 5711 4223
rect 5777 3223 5807 4223
rect 5873 3223 5903 4223
rect 5969 3223 5999 4223
rect 6065 3223 6095 4223
rect 6161 3223 6191 4223
rect 6257 3223 6287 4223
rect 6484 3230 6514 4230
rect 8084 3230 8114 4230
rect 8284 3230 8314 3830
rect 8501 3223 8531 4223
rect 8597 3223 8627 4223
rect 8693 3223 8723 4223
rect 8789 3223 8819 4223
rect 8885 3223 8915 4223
rect 8981 3223 9011 4223
rect 9077 3223 9107 4223
rect 9173 3223 9203 4223
rect 9269 3223 9299 4223
rect 9365 3223 9395 4223
rect 9461 3223 9491 4223
rect 9557 3223 9587 4223
rect 9784 3230 9814 4230
rect 11384 3230 11414 4230
rect 11584 3230 11614 3830
rect 11801 3223 11831 4223
rect 11897 3223 11927 4223
rect 11993 3223 12023 4223
rect 12089 3223 12119 4223
rect 12185 3223 12215 4223
rect 12281 3223 12311 4223
rect 12377 3223 12407 4223
rect 12473 3223 12503 4223
rect 12569 3223 12599 4223
rect 12665 3223 12695 4223
rect 12761 3223 12791 4223
rect 12857 3223 12887 4223
rect 13084 3230 13114 4230
rect 14984 3230 15014 4230
rect 15184 3230 15214 3830
rect 15401 3223 15431 4223
rect 15497 3223 15527 4223
rect 15593 3223 15623 4223
rect 15689 3223 15719 4223
rect 15785 3223 15815 4223
rect 15881 3223 15911 4223
rect 15977 3223 16007 4223
rect 16073 3223 16103 4223
rect 16169 3223 16199 4223
rect 16265 3223 16295 4223
rect 16361 3223 16391 4223
rect 16457 3223 16487 4223
rect 16684 3230 16714 4230
rect 18484 3230 18514 4230
rect 18684 3230 18714 3830
rect 18901 3223 18931 4223
rect 18997 3223 19027 4223
rect 19093 3223 19123 4223
rect 19189 3223 19219 4223
rect 19285 3223 19315 4223
rect 19381 3223 19411 4223
rect 19477 3223 19507 4223
rect 19573 3223 19603 4223
rect 19669 3223 19699 4223
rect 19765 3223 19795 4223
rect 19861 3223 19891 4223
rect 19957 3223 19987 4223
rect 20184 3230 20214 4230
rect 22184 3230 22214 4230
rect 22384 3230 22414 3830
rect 22601 3223 22631 4223
rect 22697 3223 22727 4223
rect 22793 3223 22823 4223
rect 22889 3223 22919 4223
rect 22985 3223 23015 4223
rect 23081 3223 23111 4223
rect 23177 3223 23207 4223
rect 23273 3223 23303 4223
rect 23369 3223 23399 4223
rect 23465 3223 23495 4223
rect 23561 3223 23591 4223
rect 23657 3223 23687 4223
rect 23884 3230 23914 4230
rect 25984 3230 26014 4230
rect 26184 3230 26214 3830
rect 26401 3223 26431 4223
rect 26497 3223 26527 4223
rect 26593 3223 26623 4223
rect 26689 3223 26719 4223
rect 26785 3223 26815 4223
rect 26881 3223 26911 4223
rect 26977 3223 27007 4223
rect 27073 3223 27103 4223
rect 27169 3223 27199 4223
rect 27265 3223 27295 4223
rect 27361 3223 27391 4223
rect 27457 3223 27487 4223
rect 27684 3230 27714 4230
<< scpmoshvt >>
rect 5027 26911 5145 27085
rect 5303 26911 5421 27085
rect 5588 26911 5618 27111
rect 5674 26911 5704 27111
rect 5760 26911 5790 27111
rect 5846 26911 5876 27111
rect 5942 26911 5972 27111
rect 6223 26911 7169 27085
rect 7419 26911 7537 27085
rect 7695 26911 8641 27085
rect 8799 26911 9745 27085
rect 10179 26911 10209 27069
rect 10267 26911 10297 27069
rect 10639 26911 11217 27085
rect 11375 26911 12321 27085
rect 12571 26911 12689 27085
rect 12847 26911 13793 27085
rect 13951 26911 14897 27085
rect 15147 26911 15265 27085
rect 15423 26911 16369 27085
rect 16527 26911 17473 27085
rect 17815 26911 18393 27085
rect 18560 26911 18590 27111
rect 18646 26911 18676 27111
rect 18732 26911 18762 27111
rect 18818 26911 18848 27111
rect 18914 26911 18944 27111
rect 19287 26911 19865 27085
rect 20023 26911 20141 27085
rect 5027 26643 5145 26817
rect 5487 26643 6065 26817
rect 6223 26643 7169 26817
rect 7511 26643 7905 26817
rect 8063 26643 9009 26817
rect 9167 26643 10113 26817
rect 10271 26643 11217 26817
rect 11375 26643 12321 26817
rect 12663 26643 13057 26817
rect 13215 26643 14161 26817
rect 14319 26643 15265 26817
rect 15423 26643 16369 26817
rect 16527 26643 17473 26817
rect 17815 26643 18761 26817
rect 18919 26643 19865 26817
rect 20023 26643 20141 26817
rect 5027 25823 5145 25997
rect 5487 25823 6433 25997
rect 6591 25823 7537 25997
rect 7695 25823 8641 25997
rect 8799 25823 9745 25997
rect 10087 25823 10481 25997
rect 10639 25823 11585 25997
rect 11743 25823 12689 25997
rect 12847 25823 13793 25997
rect 13951 25823 14897 25997
rect 15239 25823 15449 25997
rect 15607 25823 16553 25997
rect 16711 25823 17657 25997
rect 17815 25823 18761 25997
rect 18919 25823 19865 25997
rect 20023 25823 20141 25997
rect 5027 25555 5145 25729
rect 5487 25555 6065 25729
rect 6223 25555 7169 25729
rect 7511 25555 7905 25729
rect 8063 25555 9009 25729
rect 9167 25555 10113 25729
rect 10271 25555 11217 25729
rect 11375 25555 12321 25729
rect 12663 25555 13057 25729
rect 13215 25555 14161 25729
rect 14319 25555 15265 25729
rect 15423 25555 16369 25729
rect 16527 25555 17473 25729
rect 17815 25555 18761 25729
rect 18919 25555 19865 25729
rect 20023 25555 20141 25729
rect 5027 24735 5145 24909
rect 5487 24735 6433 24909
rect 6591 24735 7537 24909
rect 7695 24735 8641 24909
rect 8799 24735 9745 24909
rect 10087 24735 10481 24909
rect 10639 24735 11585 24909
rect 11743 24735 12689 24909
rect 12847 24735 13793 24909
rect 13951 24735 14897 24909
rect 15239 24735 15449 24909
rect 15607 24735 16553 24909
rect 16711 24735 17657 24909
rect 17815 24735 18761 24909
rect 18919 24735 19865 24909
rect 20023 24735 20141 24909
rect 5027 24467 5145 24641
rect 5487 24467 6065 24641
rect 6223 24467 7169 24641
rect 7511 24467 7905 24641
rect 8063 24467 9009 24641
rect 9167 24467 10113 24641
rect 10271 24467 11217 24641
rect 11375 24467 12321 24641
rect 12663 24467 13057 24641
rect 13215 24467 14161 24641
rect 14319 24467 15265 24641
rect 15423 24467 16369 24641
rect 16527 24467 17473 24641
rect 17815 24467 18761 24641
rect 18919 24467 19865 24641
rect 20023 24467 20141 24641
rect 5027 23647 5145 23821
rect 5487 23647 6433 23821
rect 6591 23647 7537 23821
rect 7695 23647 8641 23821
rect 8799 23647 9745 23821
rect 10087 23647 10481 23821
rect 10639 23647 11585 23821
rect 11743 23647 12689 23821
rect 12847 23647 13793 23821
rect 13951 23647 14897 23821
rect 15239 23647 15449 23821
rect 15607 23647 16553 23821
rect 16711 23647 17657 23821
rect 17815 23647 18761 23821
rect 18919 23647 19865 23821
rect 20023 23647 20141 23821
rect 5027 23379 5145 23553
rect 5487 23379 6065 23553
rect 6223 23379 7169 23553
rect 7511 23379 7905 23553
rect 8063 23379 9009 23553
rect 9167 23379 10113 23553
rect 10271 23379 11217 23553
rect 11375 23379 12321 23553
rect 12663 23379 13057 23553
rect 13215 23379 14161 23553
rect 14319 23379 15265 23553
rect 15423 23379 16369 23553
rect 16527 23379 17473 23553
rect 17815 23379 18761 23553
rect 18919 23379 19865 23553
rect 20023 23379 20141 23553
rect 5027 22559 5145 22733
rect 5487 22559 6433 22733
rect 6591 22559 7537 22733
rect 7695 22559 8641 22733
rect 8799 22559 9745 22733
rect 10087 22559 10481 22733
rect 10639 22559 11585 22733
rect 11743 22559 12689 22733
rect 12847 22559 13793 22733
rect 13951 22559 14897 22733
rect 15239 22559 15449 22733
rect 15607 22559 16553 22733
rect 16711 22559 17657 22733
rect 17815 22559 18761 22733
rect 18919 22559 19865 22733
rect 20023 22559 20141 22733
rect 5027 22291 5145 22465
rect 5487 22291 6065 22465
rect 6223 22291 7169 22465
rect 7511 22291 7905 22465
rect 8063 22291 9009 22465
rect 9167 22291 10113 22465
rect 10271 22291 11217 22465
rect 11375 22291 12321 22465
rect 12663 22291 13057 22465
rect 13215 22291 14161 22465
rect 14319 22291 15265 22465
rect 15423 22291 16369 22465
rect 16527 22291 17473 22465
rect 17815 22291 18761 22465
rect 18919 22291 19865 22465
rect 20023 22291 20141 22465
rect 5027 21471 5145 21645
rect 5487 21471 6433 21645
rect 6591 21471 7537 21645
rect 7695 21471 8641 21645
rect 8799 21471 9745 21645
rect 10087 21471 10481 21645
rect 10639 21471 11585 21645
rect 11743 21471 12689 21645
rect 12847 21471 13793 21645
rect 13951 21471 14897 21645
rect 15239 21471 15449 21645
rect 15607 21471 16553 21645
rect 16711 21471 17657 21645
rect 17815 21471 18761 21645
rect 18919 21471 19865 21645
rect 20023 21471 20141 21645
rect 5027 21203 5145 21377
rect 5487 21203 6065 21377
rect 6223 21203 7169 21377
rect 7511 21203 7905 21377
rect 8063 21203 9009 21377
rect 9167 21203 10113 21377
rect 10271 21203 11217 21377
rect 11375 21203 12321 21377
rect 12663 21203 13057 21377
rect 13215 21203 14161 21377
rect 14319 21203 15265 21377
rect 15423 21203 16369 21377
rect 16527 21203 17473 21377
rect 17815 21203 18761 21377
rect 18919 21203 19865 21377
rect 20023 21203 20141 21377
rect 5027 20383 5145 20557
rect 5487 20383 6433 20557
rect 6591 20383 7537 20557
rect 7695 20383 8641 20557
rect 8799 20383 9745 20557
rect 10087 20383 10481 20557
rect 10639 20383 11585 20557
rect 11743 20383 12689 20557
rect 12847 20383 13793 20557
rect 13951 20383 14897 20557
rect 15239 20383 15449 20557
rect 15607 20383 16553 20557
rect 16711 20383 17657 20557
rect 17815 20383 18761 20557
rect 18919 20383 19865 20557
rect 20023 20383 20141 20557
rect 5027 20115 5145 20289
rect 5487 20115 6065 20289
rect 6223 20115 7169 20289
rect 7511 20115 7905 20289
rect 8063 20115 9009 20289
rect 9167 20115 10113 20289
rect 10271 20115 11217 20289
rect 11375 20115 12321 20289
rect 12663 20115 13057 20289
rect 13215 20115 14161 20289
rect 14319 20115 15265 20289
rect 15423 20115 16369 20289
rect 16527 20115 17473 20289
rect 17815 20115 18761 20289
rect 18919 20115 19865 20289
rect 20023 20115 20141 20289
rect 5027 19295 5145 19469
rect 5487 19295 6433 19469
rect 6591 19295 7537 19469
rect 7695 19295 8641 19469
rect 8799 19295 9745 19469
rect 10087 19295 10481 19469
rect 10639 19295 11585 19469
rect 11743 19295 12689 19469
rect 12847 19295 13793 19469
rect 13951 19295 14897 19469
rect 15239 19295 15449 19469
rect 15607 19295 16553 19469
rect 16711 19295 17657 19469
rect 17815 19295 18761 19469
rect 18919 19295 19865 19469
rect 20023 19295 20141 19469
rect 5027 19027 5145 19201
rect 5487 19027 6065 19201
rect 6223 19027 7169 19201
rect 7511 19027 7905 19201
rect 8063 19027 9009 19201
rect 9167 19027 10113 19201
rect 10271 19027 11217 19201
rect 11375 19027 12321 19201
rect 12663 19027 13057 19201
rect 13215 19027 14161 19201
rect 14319 19027 15265 19201
rect 15423 19027 16369 19201
rect 16527 19027 17473 19201
rect 17815 19027 18761 19201
rect 18919 19027 19865 19201
rect 20023 19027 20141 19201
rect 5027 18207 5145 18381
rect 5487 18207 6433 18381
rect 6591 18207 7537 18381
rect 7695 18207 8641 18381
rect 8799 18207 9745 18381
rect 10087 18207 10481 18381
rect 10639 18207 11585 18381
rect 11743 18207 12689 18381
rect 12847 18207 13793 18381
rect 13951 18207 14897 18381
rect 15239 18207 15449 18381
rect 15607 18207 16553 18381
rect 16711 18207 17657 18381
rect 17815 18207 18761 18381
rect 18919 18207 19865 18381
rect 20023 18207 20141 18381
rect 5027 17939 5145 18113
rect 5487 17939 6065 18113
rect 6223 17939 7169 18113
rect 7511 17939 7905 18113
rect 8063 17939 9009 18113
rect 9167 17939 10113 18113
rect 10271 17939 11217 18113
rect 11375 17939 12321 18113
rect 12663 17939 13057 18113
rect 13215 17939 14161 18113
rect 14319 17939 15265 18113
rect 15423 17939 16369 18113
rect 16527 17939 17473 18113
rect 17815 17939 18761 18113
rect 18919 17939 19865 18113
rect 20023 17939 20141 18113
rect 5027 17119 5145 17293
rect 5487 17119 6433 17293
rect 6591 17119 7537 17293
rect 7695 17119 8641 17293
rect 8799 17119 9745 17293
rect 10087 17119 10481 17293
rect 10639 17119 11585 17293
rect 11743 17119 12689 17293
rect 12847 17119 13793 17293
rect 13951 17119 14897 17293
rect 15239 17119 15449 17293
rect 15607 17119 16553 17293
rect 16711 17119 17657 17293
rect 17815 17119 18761 17293
rect 18919 17119 19865 17293
rect 20023 17119 20141 17293
rect 5027 16851 5145 17025
rect 5487 16851 6065 17025
rect 6223 16851 7169 17025
rect 7511 16851 7905 17025
rect 8063 16851 9009 17025
rect 9167 16851 10113 17025
rect 10271 16851 11217 17025
rect 11375 16851 12321 17025
rect 12663 16851 13057 17025
rect 13215 16851 14161 17025
rect 14319 16851 15265 17025
rect 15423 16851 16369 17025
rect 16527 16851 17473 17025
rect 17815 16851 18761 17025
rect 18919 16851 19865 17025
rect 20023 16851 20141 17025
rect 5027 16031 5145 16205
rect 5487 16031 6433 16205
rect 6591 16031 7537 16205
rect 7695 16031 8641 16205
rect 8799 16031 9745 16205
rect 10087 16031 10481 16205
rect 10639 16031 11585 16205
rect 11743 16031 12689 16205
rect 12847 16031 13793 16205
rect 13951 16031 14897 16205
rect 15239 16031 15449 16205
rect 15607 16031 16553 16205
rect 16711 16031 17657 16205
rect 17815 16031 18761 16205
rect 18919 16031 19865 16205
rect 20023 16031 20141 16205
rect 5027 15763 5145 15937
rect 5487 15763 6065 15937
rect 6223 15763 7169 15937
rect 7511 15763 7905 15937
rect 8063 15763 9009 15937
rect 9167 15763 10113 15937
rect 10271 15763 11217 15937
rect 11375 15763 12321 15937
rect 12663 15763 13057 15937
rect 13215 15763 14161 15937
rect 14319 15763 15265 15937
rect 15423 15763 16369 15937
rect 16527 15763 17473 15937
rect 17815 15763 18761 15937
rect 18919 15763 19865 15937
rect 20023 15763 20141 15937
rect 5027 14943 5145 15117
rect 5487 14943 6433 15117
rect 6591 14943 7537 15117
rect 7695 14943 8641 15117
rect 8799 14943 9745 15117
rect 10087 14943 10481 15117
rect 10639 14943 11585 15117
rect 11743 14943 12689 15117
rect 12869 14943 12899 15027
rect 12953 14943 13053 15027
rect 13211 14943 13311 15027
rect 13376 14943 13406 15143
rect 13583 14943 13793 15117
rect 13951 14943 14897 15117
rect 15147 14943 15265 15117
rect 15445 14943 15475 15027
rect 15529 14943 15629 15027
rect 15787 14943 15887 15027
rect 15952 14943 15982 15143
rect 16159 14943 16553 15117
rect 16711 14943 17657 15117
rect 17815 14943 18761 15117
rect 18919 14943 19865 15117
rect 20023 14943 20141 15117
rect 5027 14675 5145 14849
rect 5487 14675 6065 14849
rect 6223 14675 7169 14849
rect 7419 14675 8365 14849
rect 8523 14675 9469 14849
rect 9627 14675 10573 14849
rect 10777 14726 10807 14810
rect 10873 14726 10903 14810
rect 10945 14726 10975 14810
rect 11159 14726 11189 14810
rect 11262 14726 11292 14810
rect 11371 14649 11401 14849
rect 11743 14675 12321 14849
rect 12801 14726 12831 14810
rect 12897 14726 12927 14810
rect 12969 14726 12999 14810
rect 13183 14726 13213 14810
rect 13286 14726 13316 14810
rect 13395 14649 13425 14849
rect 13583 14675 14161 14849
rect 14319 14691 14349 14849
rect 14407 14691 14437 14849
rect 14595 14649 14625 14849
rect 14810 14765 14840 14849
rect 14894 14765 14924 14849
rect 15002 14765 15032 14849
rect 15086 14765 15116 14849
rect 15172 14765 15202 14849
rect 15271 14681 15301 14849
rect 15468 14765 15498 14849
rect 15565 14765 15595 14849
rect 15705 14765 15735 14849
rect 15804 14765 15834 14849
rect 15896 14765 15926 14849
rect 16163 14715 16193 14843
rect 16247 14715 16277 14843
rect 16527 14675 17473 14849
rect 17815 14675 18761 14849
rect 18919 14675 19865 14849
rect 20023 14675 20141 14849
rect 5027 13855 5145 14029
rect 5487 13855 6433 14029
rect 6591 13855 7537 14029
rect 7695 13855 8641 14029
rect 8799 13855 9745 14029
rect 10179 13855 10209 14055
rect 10394 13855 10424 13939
rect 10478 13855 10508 13939
rect 10586 13855 10616 13939
rect 10670 13855 10700 13939
rect 10756 13855 10786 13939
rect 10855 13855 10885 14023
rect 11052 13855 11082 13939
rect 11149 13855 11179 13939
rect 11289 13855 11319 13939
rect 11388 13855 11418 13939
rect 11480 13855 11510 13939
rect 11747 13861 11777 13989
rect 11831 13861 11861 13989
rect 12019 13855 12049 14013
rect 12107 13855 12137 14013
rect 12313 13855 12343 14055
rect 12399 13855 12429 14055
rect 12485 13855 12515 14055
rect 12571 13855 12601 14055
rect 12657 13855 12687 14055
rect 12743 13855 12773 14055
rect 12829 13855 12859 14055
rect 12915 13855 12945 14055
rect 13000 13855 13030 14055
rect 13086 13855 13116 14055
rect 13172 13855 13202 14055
rect 13258 13855 13288 14055
rect 13344 13855 13374 14055
rect 13430 13855 13460 14055
rect 13516 13855 13546 14055
rect 13602 13855 13632 14055
rect 13688 13855 13718 14055
rect 13774 13855 13804 14055
rect 13860 13855 13890 14055
rect 13946 13855 13976 14055
rect 14341 13855 14371 13939
rect 14425 13855 14525 13939
rect 14683 13855 14783 13939
rect 14848 13855 14878 14055
rect 15239 13855 15269 14055
rect 15348 13894 15378 13978
rect 15451 13894 15481 13978
rect 15665 13894 15695 13978
rect 15737 13894 15767 13978
rect 15833 13894 15863 13978
rect 16067 13855 16097 14013
rect 16155 13855 16185 14013
rect 16343 13855 16373 14013
rect 16431 13855 16461 14013
rect 16711 13855 17657 14029
rect 17815 13855 18761 14029
rect 18919 13855 19865 14029
rect 20023 13855 20141 14029
rect 5027 13587 5145 13761
rect 5487 13587 6065 13761
rect 6223 13587 7169 13761
rect 7511 13587 8457 13761
rect 8615 13587 9561 13761
rect 9719 13603 9749 13761
rect 9807 13603 9837 13761
rect 10013 13561 10043 13761
rect 10099 13561 10129 13761
rect 10185 13561 10215 13761
rect 10271 13561 10301 13761
rect 10357 13561 10387 13761
rect 10443 13561 10473 13761
rect 10529 13561 10559 13761
rect 10615 13561 10645 13761
rect 10700 13561 10730 13761
rect 10786 13561 10816 13761
rect 10872 13561 10902 13761
rect 10958 13561 10988 13761
rect 11044 13561 11074 13761
rect 11130 13561 11160 13761
rect 11216 13561 11246 13761
rect 11302 13561 11332 13761
rect 11388 13561 11418 13761
rect 11474 13561 11504 13761
rect 11560 13561 11590 13761
rect 11646 13561 11676 13761
rect 11927 13587 12321 13761
rect 12571 13603 12601 13761
rect 12659 13603 12689 13761
rect 12939 13561 12969 13761
rect 13154 13677 13184 13761
rect 13238 13677 13268 13761
rect 13346 13677 13376 13761
rect 13430 13677 13460 13761
rect 13516 13677 13546 13761
rect 13615 13593 13645 13761
rect 13812 13677 13842 13761
rect 13909 13677 13939 13761
rect 14049 13677 14079 13761
rect 14148 13677 14178 13761
rect 14240 13677 14270 13761
rect 14507 13627 14537 13755
rect 14591 13627 14621 13755
rect 14780 13561 14810 13761
rect 14866 13561 14896 13761
rect 14952 13561 14982 13761
rect 15038 13561 15068 13761
rect 15124 13561 15154 13761
rect 15210 13561 15240 13761
rect 15296 13561 15326 13761
rect 15382 13561 15412 13761
rect 15468 13561 15498 13761
rect 15554 13561 15584 13761
rect 15640 13561 15670 13761
rect 15726 13561 15756 13761
rect 15811 13561 15841 13761
rect 15897 13561 15927 13761
rect 15983 13561 16013 13761
rect 16069 13561 16099 13761
rect 16155 13561 16185 13761
rect 16241 13561 16271 13761
rect 16327 13561 16357 13761
rect 16413 13561 16443 13761
rect 16619 13561 16649 13761
rect 16728 13638 16758 13722
rect 16831 13638 16861 13722
rect 17045 13638 17075 13722
rect 17117 13638 17147 13722
rect 17213 13638 17243 13722
rect 17815 13587 18761 13761
rect 18919 13587 19865 13761
rect 20023 13587 20141 13761
rect 5027 12767 5145 12941
rect 5303 12767 5697 12941
rect 5855 12767 6801 12941
rect 6959 12767 7905 12941
rect 8063 12767 9009 12941
rect 9189 12767 9219 12851
rect 9273 12767 9373 12851
rect 9531 12767 9631 12851
rect 9696 12767 9726 12967
rect 10087 12767 10297 12941
rect 10455 12767 10485 12967
rect 10670 12767 10700 12851
rect 10754 12767 10784 12851
rect 10862 12767 10892 12851
rect 10946 12767 10976 12851
rect 11032 12767 11062 12851
rect 11131 12767 11161 12935
rect 11328 12767 11358 12851
rect 11425 12767 11455 12851
rect 11565 12767 11595 12851
rect 11664 12767 11694 12851
rect 11756 12767 11786 12851
rect 12023 12773 12053 12901
rect 12107 12773 12137 12901
rect 12295 12773 12325 12901
rect 12379 12773 12409 12901
rect 12646 12767 12676 12851
rect 12738 12767 12768 12851
rect 12837 12767 12867 12851
rect 12977 12767 13007 12851
rect 13074 12767 13104 12851
rect 13271 12767 13301 12935
rect 13370 12767 13400 12851
rect 13456 12767 13486 12851
rect 13540 12767 13570 12851
rect 13648 12767 13678 12851
rect 13732 12767 13762 12851
rect 13947 12767 13977 12967
rect 14135 12767 14165 12967
rect 14244 12806 14274 12890
rect 14347 12806 14377 12890
rect 14561 12806 14591 12890
rect 14633 12806 14663 12890
rect 14729 12806 14759 12890
rect 15147 12767 15177 12967
rect 15362 12767 15392 12851
rect 15446 12767 15476 12851
rect 15554 12767 15584 12851
rect 15638 12767 15668 12851
rect 15724 12767 15754 12851
rect 15823 12767 15853 12935
rect 16020 12767 16050 12851
rect 16117 12767 16147 12851
rect 16257 12767 16287 12851
rect 16356 12767 16386 12851
rect 16448 12767 16478 12851
rect 16715 12773 16745 12901
rect 16799 12773 16829 12901
rect 17006 12767 17036 12967
rect 17101 12767 17201 12851
rect 17359 12767 17459 12851
rect 17513 12767 17543 12851
rect 17815 12767 18761 12941
rect 18919 12767 19865 12941
rect 20023 12767 20141 12941
rect 5027 12499 5145 12673
rect 5671 12499 6617 12673
rect 6784 12473 6814 12673
rect 6870 12473 6900 12673
rect 6956 12473 6986 12673
rect 7042 12473 7072 12673
rect 7138 12473 7168 12673
rect 7419 12499 7629 12673
rect 7787 12499 8733 12673
rect 8900 12473 8930 12673
rect 8986 12473 9016 12673
rect 9072 12473 9102 12673
rect 9158 12473 9188 12673
rect 9254 12473 9284 12673
rect 9535 12499 9745 12673
rect 10004 12473 10034 12673
rect 10090 12473 10120 12673
rect 10176 12473 10206 12673
rect 10262 12473 10292 12673
rect 10358 12473 10388 12673
rect 10547 12473 10577 12673
rect 10656 12550 10686 12634
rect 10759 12550 10789 12634
rect 10973 12550 11003 12634
rect 11045 12550 11075 12634
rect 11141 12550 11171 12634
rect 11513 12550 11543 12634
rect 11609 12550 11639 12634
rect 11681 12550 11711 12634
rect 11895 12550 11925 12634
rect 11998 12550 12028 12634
rect 12107 12473 12137 12673
rect 12764 12473 12794 12673
rect 12850 12473 12880 12673
rect 12936 12473 12966 12673
rect 13022 12473 13052 12673
rect 13118 12473 13148 12673
rect 13308 12473 13338 12673
rect 13404 12473 13434 12673
rect 13490 12473 13520 12673
rect 13576 12473 13606 12673
rect 13662 12473 13692 12673
rect 13859 12515 13889 12673
rect 13947 12515 13977 12673
rect 14157 12589 14187 12673
rect 14241 12589 14341 12673
rect 14499 12589 14599 12673
rect 14664 12473 14694 12673
rect 15147 12539 15177 12667
rect 15231 12539 15261 12667
rect 15498 12589 15528 12673
rect 15590 12589 15620 12673
rect 15689 12589 15719 12673
rect 15829 12589 15859 12673
rect 15926 12589 15956 12673
rect 16123 12505 16153 12673
rect 16222 12589 16252 12673
rect 16308 12589 16338 12673
rect 16392 12589 16422 12673
rect 16500 12589 16530 12673
rect 16584 12589 16614 12673
rect 16799 12473 16829 12673
rect 17080 12473 17110 12673
rect 17176 12473 17206 12673
rect 17262 12473 17292 12673
rect 17348 12473 17378 12673
rect 17434 12473 17464 12673
rect 17815 12499 18209 12673
rect 18367 12499 19313 12673
rect 19472 12473 19502 12673
rect 19568 12473 19598 12673
rect 19654 12473 19684 12673
rect 19740 12473 19770 12673
rect 19826 12473 19856 12673
rect 20023 12499 20141 12673
<< ndiff >>
rect 4975 27328 5027 27361
rect 4975 27294 4983 27328
rect 5017 27294 5027 27328
rect 4975 27251 5027 27294
rect 5145 27328 5197 27361
rect 5145 27294 5155 27328
rect 5189 27294 5197 27328
rect 5145 27251 5197 27294
rect 5251 27328 5303 27361
rect 5251 27294 5259 27328
rect 5293 27294 5303 27328
rect 5251 27251 5303 27294
rect 5421 27328 5473 27361
rect 5421 27294 5431 27328
rect 5465 27294 5473 27328
rect 5421 27251 5473 27294
rect 5529 27345 5587 27361
rect 5529 27311 5542 27345
rect 5576 27311 5587 27345
rect 5529 27277 5587 27311
rect 5617 27323 5673 27361
rect 5617 27289 5628 27323
rect 5662 27289 5673 27323
rect 5617 27277 5673 27289
rect 5703 27345 5759 27361
rect 5703 27311 5714 27345
rect 5748 27311 5759 27345
rect 5703 27277 5759 27311
rect 5789 27323 5845 27361
rect 5789 27289 5800 27323
rect 5834 27289 5845 27323
rect 5789 27277 5845 27289
rect 5875 27345 5942 27361
rect 5875 27311 5897 27345
rect 5931 27311 5942 27345
rect 5875 27277 5942 27311
rect 5972 27341 6025 27361
rect 5972 27307 5983 27341
rect 6017 27307 6025 27341
rect 5972 27277 6025 27307
rect 6171 27330 6223 27361
rect 6171 27296 6179 27330
rect 6213 27296 6223 27330
rect 6171 27251 6223 27296
rect 7169 27330 7221 27361
rect 7169 27296 7179 27330
rect 7213 27296 7221 27330
rect 7169 27251 7221 27296
rect 7367 27328 7419 27361
rect 7367 27294 7375 27328
rect 7409 27294 7419 27328
rect 7367 27251 7419 27294
rect 7537 27328 7589 27361
rect 7537 27294 7547 27328
rect 7581 27294 7589 27328
rect 7537 27251 7589 27294
rect 7643 27330 7695 27361
rect 7643 27296 7651 27330
rect 7685 27296 7695 27330
rect 7643 27251 7695 27296
rect 8641 27330 8693 27361
rect 8641 27296 8651 27330
rect 8685 27296 8693 27330
rect 8641 27251 8693 27296
rect 8747 27330 8799 27361
rect 8747 27296 8755 27330
rect 8789 27296 8799 27330
rect 8747 27251 8799 27296
rect 9745 27330 9797 27361
rect 9745 27296 9755 27330
rect 9789 27296 9797 27330
rect 9745 27251 9797 27296
rect 10127 27336 10179 27361
rect 10127 27302 10135 27336
rect 10169 27302 10179 27336
rect 10127 27257 10179 27302
rect 10209 27349 10267 27361
rect 10209 27315 10221 27349
rect 10255 27315 10267 27349
rect 10209 27257 10267 27315
rect 10297 27319 10349 27361
rect 10297 27285 10307 27319
rect 10341 27285 10349 27319
rect 10297 27257 10349 27285
rect 10587 27330 10639 27361
rect 10587 27296 10595 27330
rect 10629 27296 10639 27330
rect 10587 27251 10639 27296
rect 11217 27330 11269 27361
rect 11217 27296 11227 27330
rect 11261 27296 11269 27330
rect 11217 27251 11269 27296
rect 11323 27330 11375 27361
rect 11323 27296 11331 27330
rect 11365 27296 11375 27330
rect 11323 27251 11375 27296
rect 12321 27330 12373 27361
rect 12321 27296 12331 27330
rect 12365 27296 12373 27330
rect 12321 27251 12373 27296
rect 12519 27328 12571 27361
rect 12519 27294 12527 27328
rect 12561 27294 12571 27328
rect 12519 27251 12571 27294
rect 12689 27328 12741 27361
rect 12689 27294 12699 27328
rect 12733 27294 12741 27328
rect 12689 27251 12741 27294
rect 12795 27330 12847 27361
rect 12795 27296 12803 27330
rect 12837 27296 12847 27330
rect 12795 27251 12847 27296
rect 13793 27330 13845 27361
rect 13793 27296 13803 27330
rect 13837 27296 13845 27330
rect 13793 27251 13845 27296
rect 13899 27330 13951 27361
rect 13899 27296 13907 27330
rect 13941 27296 13951 27330
rect 13899 27251 13951 27296
rect 14897 27330 14949 27361
rect 14897 27296 14907 27330
rect 14941 27296 14949 27330
rect 14897 27251 14949 27296
rect 15095 27328 15147 27361
rect 15095 27294 15103 27328
rect 15137 27294 15147 27328
rect 15095 27251 15147 27294
rect 15265 27328 15317 27361
rect 15265 27294 15275 27328
rect 15309 27294 15317 27328
rect 15265 27251 15317 27294
rect 15371 27330 15423 27361
rect 15371 27296 15379 27330
rect 15413 27296 15423 27330
rect 15371 27251 15423 27296
rect 16369 27330 16421 27361
rect 16369 27296 16379 27330
rect 16413 27296 16421 27330
rect 16369 27251 16421 27296
rect 16475 27330 16527 27361
rect 16475 27296 16483 27330
rect 16517 27296 16527 27330
rect 16475 27251 16527 27296
rect 17473 27330 17525 27361
rect 17473 27296 17483 27330
rect 17517 27296 17525 27330
rect 17473 27251 17525 27296
rect 17763 27330 17815 27361
rect 17763 27296 17771 27330
rect 17805 27296 17815 27330
rect 17763 27251 17815 27296
rect 18393 27330 18445 27361
rect 18393 27296 18403 27330
rect 18437 27296 18445 27330
rect 18393 27251 18445 27296
rect 18501 27345 18559 27361
rect 18501 27311 18514 27345
rect 18548 27311 18559 27345
rect 18501 27277 18559 27311
rect 18589 27323 18645 27361
rect 18589 27289 18600 27323
rect 18634 27289 18645 27323
rect 18589 27277 18645 27289
rect 18675 27345 18731 27361
rect 18675 27311 18686 27345
rect 18720 27311 18731 27345
rect 18675 27277 18731 27311
rect 18761 27323 18817 27361
rect 18761 27289 18772 27323
rect 18806 27289 18817 27323
rect 18761 27277 18817 27289
rect 18847 27345 18914 27361
rect 18847 27311 18869 27345
rect 18903 27311 18914 27345
rect 18847 27277 18914 27311
rect 18944 27341 18997 27361
rect 18944 27307 18955 27341
rect 18989 27307 18997 27341
rect 18944 27277 18997 27307
rect 19235 27330 19287 27361
rect 19235 27296 19243 27330
rect 19277 27296 19287 27330
rect 19235 27251 19287 27296
rect 19865 27330 19917 27361
rect 19865 27296 19875 27330
rect 19909 27296 19917 27330
rect 19865 27251 19917 27296
rect 19971 27328 20023 27361
rect 19971 27294 19979 27328
rect 20013 27294 20023 27328
rect 19971 27251 20023 27294
rect 20141 27328 20193 27361
rect 20141 27294 20151 27328
rect 20185 27294 20193 27328
rect 20141 27251 20193 27294
rect 4975 26434 5027 26477
rect 4975 26400 4983 26434
rect 5017 26400 5027 26434
rect 4975 26367 5027 26400
rect 5145 26434 5197 26477
rect 5145 26400 5155 26434
rect 5189 26400 5197 26434
rect 5145 26367 5197 26400
rect 5435 26432 5487 26477
rect 5435 26398 5443 26432
rect 5477 26398 5487 26432
rect 5435 26367 5487 26398
rect 6065 26432 6117 26477
rect 6065 26398 6075 26432
rect 6109 26398 6117 26432
rect 6065 26367 6117 26398
rect 6171 26432 6223 26477
rect 6171 26398 6179 26432
rect 6213 26398 6223 26432
rect 6171 26367 6223 26398
rect 7169 26432 7221 26477
rect 7169 26398 7179 26432
rect 7213 26398 7221 26432
rect 7169 26367 7221 26398
rect 7459 26432 7511 26477
rect 7459 26398 7467 26432
rect 7501 26398 7511 26432
rect 7459 26367 7511 26398
rect 7905 26432 7957 26477
rect 7905 26398 7915 26432
rect 7949 26398 7957 26432
rect 7905 26367 7957 26398
rect 8011 26432 8063 26477
rect 8011 26398 8019 26432
rect 8053 26398 8063 26432
rect 8011 26367 8063 26398
rect 9009 26432 9061 26477
rect 9009 26398 9019 26432
rect 9053 26398 9061 26432
rect 9009 26367 9061 26398
rect 9115 26432 9167 26477
rect 9115 26398 9123 26432
rect 9157 26398 9167 26432
rect 9115 26367 9167 26398
rect 10113 26432 10165 26477
rect 10113 26398 10123 26432
rect 10157 26398 10165 26432
rect 10113 26367 10165 26398
rect 10219 26432 10271 26477
rect 10219 26398 10227 26432
rect 10261 26398 10271 26432
rect 10219 26367 10271 26398
rect 11217 26432 11269 26477
rect 11217 26398 11227 26432
rect 11261 26398 11269 26432
rect 11217 26367 11269 26398
rect 11323 26432 11375 26477
rect 11323 26398 11331 26432
rect 11365 26398 11375 26432
rect 11323 26367 11375 26398
rect 12321 26432 12373 26477
rect 12321 26398 12331 26432
rect 12365 26398 12373 26432
rect 12321 26367 12373 26398
rect 12611 26432 12663 26477
rect 12611 26398 12619 26432
rect 12653 26398 12663 26432
rect 12611 26367 12663 26398
rect 13057 26432 13109 26477
rect 13057 26398 13067 26432
rect 13101 26398 13109 26432
rect 13057 26367 13109 26398
rect 13163 26432 13215 26477
rect 13163 26398 13171 26432
rect 13205 26398 13215 26432
rect 13163 26367 13215 26398
rect 14161 26432 14213 26477
rect 14161 26398 14171 26432
rect 14205 26398 14213 26432
rect 14161 26367 14213 26398
rect 14267 26432 14319 26477
rect 14267 26398 14275 26432
rect 14309 26398 14319 26432
rect 14267 26367 14319 26398
rect 15265 26432 15317 26477
rect 15265 26398 15275 26432
rect 15309 26398 15317 26432
rect 15265 26367 15317 26398
rect 15371 26432 15423 26477
rect 15371 26398 15379 26432
rect 15413 26398 15423 26432
rect 15371 26367 15423 26398
rect 16369 26432 16421 26477
rect 16369 26398 16379 26432
rect 16413 26398 16421 26432
rect 16369 26367 16421 26398
rect 16475 26432 16527 26477
rect 16475 26398 16483 26432
rect 16517 26398 16527 26432
rect 16475 26367 16527 26398
rect 17473 26432 17525 26477
rect 17473 26398 17483 26432
rect 17517 26398 17525 26432
rect 17473 26367 17525 26398
rect 17763 26432 17815 26477
rect 17763 26398 17771 26432
rect 17805 26398 17815 26432
rect 17763 26367 17815 26398
rect 18761 26432 18813 26477
rect 18761 26398 18771 26432
rect 18805 26398 18813 26432
rect 18761 26367 18813 26398
rect 18867 26432 18919 26477
rect 18867 26398 18875 26432
rect 18909 26398 18919 26432
rect 18867 26367 18919 26398
rect 19865 26432 19917 26477
rect 19865 26398 19875 26432
rect 19909 26398 19917 26432
rect 19865 26367 19917 26398
rect 19971 26434 20023 26477
rect 19971 26400 19979 26434
rect 20013 26400 20023 26434
rect 19971 26367 20023 26400
rect 20141 26434 20193 26477
rect 20141 26400 20151 26434
rect 20185 26400 20193 26434
rect 20141 26367 20193 26400
rect 4975 26240 5027 26273
rect 4975 26206 4983 26240
rect 5017 26206 5027 26240
rect 4975 26163 5027 26206
rect 5145 26240 5197 26273
rect 5145 26206 5155 26240
rect 5189 26206 5197 26240
rect 5145 26163 5197 26206
rect 5435 26242 5487 26273
rect 5435 26208 5443 26242
rect 5477 26208 5487 26242
rect 5435 26163 5487 26208
rect 6433 26242 6485 26273
rect 6433 26208 6443 26242
rect 6477 26208 6485 26242
rect 6433 26163 6485 26208
rect 6539 26242 6591 26273
rect 6539 26208 6547 26242
rect 6581 26208 6591 26242
rect 6539 26163 6591 26208
rect 7537 26242 7589 26273
rect 7537 26208 7547 26242
rect 7581 26208 7589 26242
rect 7537 26163 7589 26208
rect 7643 26242 7695 26273
rect 7643 26208 7651 26242
rect 7685 26208 7695 26242
rect 7643 26163 7695 26208
rect 8641 26242 8693 26273
rect 8641 26208 8651 26242
rect 8685 26208 8693 26242
rect 8641 26163 8693 26208
rect 8747 26242 8799 26273
rect 8747 26208 8755 26242
rect 8789 26208 8799 26242
rect 8747 26163 8799 26208
rect 9745 26242 9797 26273
rect 9745 26208 9755 26242
rect 9789 26208 9797 26242
rect 9745 26163 9797 26208
rect 10035 26242 10087 26273
rect 10035 26208 10043 26242
rect 10077 26208 10087 26242
rect 10035 26163 10087 26208
rect 10481 26242 10533 26273
rect 10481 26208 10491 26242
rect 10525 26208 10533 26242
rect 10481 26163 10533 26208
rect 10587 26242 10639 26273
rect 10587 26208 10595 26242
rect 10629 26208 10639 26242
rect 10587 26163 10639 26208
rect 11585 26242 11637 26273
rect 11585 26208 11595 26242
rect 11629 26208 11637 26242
rect 11585 26163 11637 26208
rect 11691 26242 11743 26273
rect 11691 26208 11699 26242
rect 11733 26208 11743 26242
rect 11691 26163 11743 26208
rect 12689 26242 12741 26273
rect 12689 26208 12699 26242
rect 12733 26208 12741 26242
rect 12689 26163 12741 26208
rect 12795 26242 12847 26273
rect 12795 26208 12803 26242
rect 12837 26208 12847 26242
rect 12795 26163 12847 26208
rect 13793 26242 13845 26273
rect 13793 26208 13803 26242
rect 13837 26208 13845 26242
rect 13793 26163 13845 26208
rect 13899 26242 13951 26273
rect 13899 26208 13907 26242
rect 13941 26208 13951 26242
rect 13899 26163 13951 26208
rect 14897 26242 14949 26273
rect 14897 26208 14907 26242
rect 14941 26208 14949 26242
rect 14897 26163 14949 26208
rect 15187 26235 15239 26273
rect 15187 26201 15195 26235
rect 15229 26201 15239 26235
rect 15187 26163 15239 26201
rect 15449 26235 15501 26273
rect 15449 26201 15459 26235
rect 15493 26201 15501 26235
rect 15449 26163 15501 26201
rect 15555 26242 15607 26273
rect 15555 26208 15563 26242
rect 15597 26208 15607 26242
rect 15555 26163 15607 26208
rect 16553 26242 16605 26273
rect 16553 26208 16563 26242
rect 16597 26208 16605 26242
rect 16553 26163 16605 26208
rect 16659 26242 16711 26273
rect 16659 26208 16667 26242
rect 16701 26208 16711 26242
rect 16659 26163 16711 26208
rect 17657 26242 17709 26273
rect 17657 26208 17667 26242
rect 17701 26208 17709 26242
rect 17657 26163 17709 26208
rect 17763 26242 17815 26273
rect 17763 26208 17771 26242
rect 17805 26208 17815 26242
rect 17763 26163 17815 26208
rect 18761 26242 18813 26273
rect 18761 26208 18771 26242
rect 18805 26208 18813 26242
rect 18761 26163 18813 26208
rect 18867 26242 18919 26273
rect 18867 26208 18875 26242
rect 18909 26208 18919 26242
rect 18867 26163 18919 26208
rect 19865 26242 19917 26273
rect 19865 26208 19875 26242
rect 19909 26208 19917 26242
rect 19865 26163 19917 26208
rect 19971 26240 20023 26273
rect 19971 26206 19979 26240
rect 20013 26206 20023 26240
rect 19971 26163 20023 26206
rect 20141 26240 20193 26273
rect 20141 26206 20151 26240
rect 20185 26206 20193 26240
rect 20141 26163 20193 26206
rect 4975 25346 5027 25389
rect 4975 25312 4983 25346
rect 5017 25312 5027 25346
rect 4975 25279 5027 25312
rect 5145 25346 5197 25389
rect 5145 25312 5155 25346
rect 5189 25312 5197 25346
rect 5145 25279 5197 25312
rect 5435 25344 5487 25389
rect 5435 25310 5443 25344
rect 5477 25310 5487 25344
rect 5435 25279 5487 25310
rect 6065 25344 6117 25389
rect 6065 25310 6075 25344
rect 6109 25310 6117 25344
rect 6065 25279 6117 25310
rect 6171 25344 6223 25389
rect 6171 25310 6179 25344
rect 6213 25310 6223 25344
rect 6171 25279 6223 25310
rect 7169 25344 7221 25389
rect 7169 25310 7179 25344
rect 7213 25310 7221 25344
rect 7169 25279 7221 25310
rect 7459 25344 7511 25389
rect 7459 25310 7467 25344
rect 7501 25310 7511 25344
rect 7459 25279 7511 25310
rect 7905 25344 7957 25389
rect 7905 25310 7915 25344
rect 7949 25310 7957 25344
rect 7905 25279 7957 25310
rect 8011 25344 8063 25389
rect 8011 25310 8019 25344
rect 8053 25310 8063 25344
rect 8011 25279 8063 25310
rect 9009 25344 9061 25389
rect 9009 25310 9019 25344
rect 9053 25310 9061 25344
rect 9009 25279 9061 25310
rect 9115 25344 9167 25389
rect 9115 25310 9123 25344
rect 9157 25310 9167 25344
rect 9115 25279 9167 25310
rect 10113 25344 10165 25389
rect 10113 25310 10123 25344
rect 10157 25310 10165 25344
rect 10113 25279 10165 25310
rect 10219 25344 10271 25389
rect 10219 25310 10227 25344
rect 10261 25310 10271 25344
rect 10219 25279 10271 25310
rect 11217 25344 11269 25389
rect 11217 25310 11227 25344
rect 11261 25310 11269 25344
rect 11217 25279 11269 25310
rect 11323 25344 11375 25389
rect 11323 25310 11331 25344
rect 11365 25310 11375 25344
rect 11323 25279 11375 25310
rect 12321 25344 12373 25389
rect 12321 25310 12331 25344
rect 12365 25310 12373 25344
rect 12321 25279 12373 25310
rect 12611 25344 12663 25389
rect 12611 25310 12619 25344
rect 12653 25310 12663 25344
rect 12611 25279 12663 25310
rect 13057 25344 13109 25389
rect 13057 25310 13067 25344
rect 13101 25310 13109 25344
rect 13057 25279 13109 25310
rect 13163 25344 13215 25389
rect 13163 25310 13171 25344
rect 13205 25310 13215 25344
rect 13163 25279 13215 25310
rect 14161 25344 14213 25389
rect 14161 25310 14171 25344
rect 14205 25310 14213 25344
rect 14161 25279 14213 25310
rect 14267 25344 14319 25389
rect 14267 25310 14275 25344
rect 14309 25310 14319 25344
rect 14267 25279 14319 25310
rect 15265 25344 15317 25389
rect 15265 25310 15275 25344
rect 15309 25310 15317 25344
rect 15265 25279 15317 25310
rect 15371 25344 15423 25389
rect 15371 25310 15379 25344
rect 15413 25310 15423 25344
rect 15371 25279 15423 25310
rect 16369 25344 16421 25389
rect 16369 25310 16379 25344
rect 16413 25310 16421 25344
rect 16369 25279 16421 25310
rect 16475 25344 16527 25389
rect 16475 25310 16483 25344
rect 16517 25310 16527 25344
rect 16475 25279 16527 25310
rect 17473 25344 17525 25389
rect 17473 25310 17483 25344
rect 17517 25310 17525 25344
rect 17473 25279 17525 25310
rect 17763 25344 17815 25389
rect 17763 25310 17771 25344
rect 17805 25310 17815 25344
rect 17763 25279 17815 25310
rect 18761 25344 18813 25389
rect 18761 25310 18771 25344
rect 18805 25310 18813 25344
rect 18761 25279 18813 25310
rect 18867 25344 18919 25389
rect 18867 25310 18875 25344
rect 18909 25310 18919 25344
rect 18867 25279 18919 25310
rect 19865 25344 19917 25389
rect 19865 25310 19875 25344
rect 19909 25310 19917 25344
rect 19865 25279 19917 25310
rect 19971 25346 20023 25389
rect 19971 25312 19979 25346
rect 20013 25312 20023 25346
rect 19971 25279 20023 25312
rect 20141 25346 20193 25389
rect 20141 25312 20151 25346
rect 20185 25312 20193 25346
rect 20141 25279 20193 25312
rect 4975 25152 5027 25185
rect 4975 25118 4983 25152
rect 5017 25118 5027 25152
rect 4975 25075 5027 25118
rect 5145 25152 5197 25185
rect 5145 25118 5155 25152
rect 5189 25118 5197 25152
rect 5145 25075 5197 25118
rect 5435 25154 5487 25185
rect 5435 25120 5443 25154
rect 5477 25120 5487 25154
rect 5435 25075 5487 25120
rect 6433 25154 6485 25185
rect 6433 25120 6443 25154
rect 6477 25120 6485 25154
rect 6433 25075 6485 25120
rect 6539 25154 6591 25185
rect 6539 25120 6547 25154
rect 6581 25120 6591 25154
rect 6539 25075 6591 25120
rect 7537 25154 7589 25185
rect 7537 25120 7547 25154
rect 7581 25120 7589 25154
rect 7537 25075 7589 25120
rect 7643 25154 7695 25185
rect 7643 25120 7651 25154
rect 7685 25120 7695 25154
rect 7643 25075 7695 25120
rect 8641 25154 8693 25185
rect 8641 25120 8651 25154
rect 8685 25120 8693 25154
rect 8641 25075 8693 25120
rect 8747 25154 8799 25185
rect 8747 25120 8755 25154
rect 8789 25120 8799 25154
rect 8747 25075 8799 25120
rect 9745 25154 9797 25185
rect 9745 25120 9755 25154
rect 9789 25120 9797 25154
rect 9745 25075 9797 25120
rect 10035 25154 10087 25185
rect 10035 25120 10043 25154
rect 10077 25120 10087 25154
rect 10035 25075 10087 25120
rect 10481 25154 10533 25185
rect 10481 25120 10491 25154
rect 10525 25120 10533 25154
rect 10481 25075 10533 25120
rect 10587 25154 10639 25185
rect 10587 25120 10595 25154
rect 10629 25120 10639 25154
rect 10587 25075 10639 25120
rect 11585 25154 11637 25185
rect 11585 25120 11595 25154
rect 11629 25120 11637 25154
rect 11585 25075 11637 25120
rect 11691 25154 11743 25185
rect 11691 25120 11699 25154
rect 11733 25120 11743 25154
rect 11691 25075 11743 25120
rect 12689 25154 12741 25185
rect 12689 25120 12699 25154
rect 12733 25120 12741 25154
rect 12689 25075 12741 25120
rect 12795 25154 12847 25185
rect 12795 25120 12803 25154
rect 12837 25120 12847 25154
rect 12795 25075 12847 25120
rect 13793 25154 13845 25185
rect 13793 25120 13803 25154
rect 13837 25120 13845 25154
rect 13793 25075 13845 25120
rect 13899 25154 13951 25185
rect 13899 25120 13907 25154
rect 13941 25120 13951 25154
rect 13899 25075 13951 25120
rect 14897 25154 14949 25185
rect 14897 25120 14907 25154
rect 14941 25120 14949 25154
rect 14897 25075 14949 25120
rect 15187 25147 15239 25185
rect 15187 25113 15195 25147
rect 15229 25113 15239 25147
rect 15187 25075 15239 25113
rect 15449 25147 15501 25185
rect 15449 25113 15459 25147
rect 15493 25113 15501 25147
rect 15449 25075 15501 25113
rect 15555 25154 15607 25185
rect 15555 25120 15563 25154
rect 15597 25120 15607 25154
rect 15555 25075 15607 25120
rect 16553 25154 16605 25185
rect 16553 25120 16563 25154
rect 16597 25120 16605 25154
rect 16553 25075 16605 25120
rect 16659 25154 16711 25185
rect 16659 25120 16667 25154
rect 16701 25120 16711 25154
rect 16659 25075 16711 25120
rect 17657 25154 17709 25185
rect 17657 25120 17667 25154
rect 17701 25120 17709 25154
rect 17657 25075 17709 25120
rect 17763 25154 17815 25185
rect 17763 25120 17771 25154
rect 17805 25120 17815 25154
rect 17763 25075 17815 25120
rect 18761 25154 18813 25185
rect 18761 25120 18771 25154
rect 18805 25120 18813 25154
rect 18761 25075 18813 25120
rect 18867 25154 18919 25185
rect 18867 25120 18875 25154
rect 18909 25120 18919 25154
rect 18867 25075 18919 25120
rect 19865 25154 19917 25185
rect 19865 25120 19875 25154
rect 19909 25120 19917 25154
rect 19865 25075 19917 25120
rect 19971 25152 20023 25185
rect 19971 25118 19979 25152
rect 20013 25118 20023 25152
rect 19971 25075 20023 25118
rect 20141 25152 20193 25185
rect 20141 25118 20151 25152
rect 20185 25118 20193 25152
rect 20141 25075 20193 25118
rect 4975 24258 5027 24301
rect 4975 24224 4983 24258
rect 5017 24224 5027 24258
rect 4975 24191 5027 24224
rect 5145 24258 5197 24301
rect 5145 24224 5155 24258
rect 5189 24224 5197 24258
rect 5145 24191 5197 24224
rect 5435 24256 5487 24301
rect 5435 24222 5443 24256
rect 5477 24222 5487 24256
rect 5435 24191 5487 24222
rect 6065 24256 6117 24301
rect 6065 24222 6075 24256
rect 6109 24222 6117 24256
rect 6065 24191 6117 24222
rect 6171 24256 6223 24301
rect 6171 24222 6179 24256
rect 6213 24222 6223 24256
rect 6171 24191 6223 24222
rect 7169 24256 7221 24301
rect 7169 24222 7179 24256
rect 7213 24222 7221 24256
rect 7169 24191 7221 24222
rect 7459 24256 7511 24301
rect 7459 24222 7467 24256
rect 7501 24222 7511 24256
rect 7459 24191 7511 24222
rect 7905 24256 7957 24301
rect 7905 24222 7915 24256
rect 7949 24222 7957 24256
rect 7905 24191 7957 24222
rect 8011 24256 8063 24301
rect 8011 24222 8019 24256
rect 8053 24222 8063 24256
rect 8011 24191 8063 24222
rect 9009 24256 9061 24301
rect 9009 24222 9019 24256
rect 9053 24222 9061 24256
rect 9009 24191 9061 24222
rect 9115 24256 9167 24301
rect 9115 24222 9123 24256
rect 9157 24222 9167 24256
rect 9115 24191 9167 24222
rect 10113 24256 10165 24301
rect 10113 24222 10123 24256
rect 10157 24222 10165 24256
rect 10113 24191 10165 24222
rect 10219 24256 10271 24301
rect 10219 24222 10227 24256
rect 10261 24222 10271 24256
rect 10219 24191 10271 24222
rect 11217 24256 11269 24301
rect 11217 24222 11227 24256
rect 11261 24222 11269 24256
rect 11217 24191 11269 24222
rect 11323 24256 11375 24301
rect 11323 24222 11331 24256
rect 11365 24222 11375 24256
rect 11323 24191 11375 24222
rect 12321 24256 12373 24301
rect 12321 24222 12331 24256
rect 12365 24222 12373 24256
rect 12321 24191 12373 24222
rect 12611 24256 12663 24301
rect 12611 24222 12619 24256
rect 12653 24222 12663 24256
rect 12611 24191 12663 24222
rect 13057 24256 13109 24301
rect 13057 24222 13067 24256
rect 13101 24222 13109 24256
rect 13057 24191 13109 24222
rect 13163 24256 13215 24301
rect 13163 24222 13171 24256
rect 13205 24222 13215 24256
rect 13163 24191 13215 24222
rect 14161 24256 14213 24301
rect 14161 24222 14171 24256
rect 14205 24222 14213 24256
rect 14161 24191 14213 24222
rect 14267 24256 14319 24301
rect 14267 24222 14275 24256
rect 14309 24222 14319 24256
rect 14267 24191 14319 24222
rect 15265 24256 15317 24301
rect 15265 24222 15275 24256
rect 15309 24222 15317 24256
rect 15265 24191 15317 24222
rect 15371 24256 15423 24301
rect 15371 24222 15379 24256
rect 15413 24222 15423 24256
rect 15371 24191 15423 24222
rect 16369 24256 16421 24301
rect 16369 24222 16379 24256
rect 16413 24222 16421 24256
rect 16369 24191 16421 24222
rect 16475 24256 16527 24301
rect 16475 24222 16483 24256
rect 16517 24222 16527 24256
rect 16475 24191 16527 24222
rect 17473 24256 17525 24301
rect 17473 24222 17483 24256
rect 17517 24222 17525 24256
rect 17473 24191 17525 24222
rect 17763 24256 17815 24301
rect 17763 24222 17771 24256
rect 17805 24222 17815 24256
rect 17763 24191 17815 24222
rect 18761 24256 18813 24301
rect 18761 24222 18771 24256
rect 18805 24222 18813 24256
rect 18761 24191 18813 24222
rect 18867 24256 18919 24301
rect 18867 24222 18875 24256
rect 18909 24222 18919 24256
rect 18867 24191 18919 24222
rect 19865 24256 19917 24301
rect 19865 24222 19875 24256
rect 19909 24222 19917 24256
rect 19865 24191 19917 24222
rect 19971 24258 20023 24301
rect 19971 24224 19979 24258
rect 20013 24224 20023 24258
rect 19971 24191 20023 24224
rect 20141 24258 20193 24301
rect 20141 24224 20151 24258
rect 20185 24224 20193 24258
rect 20141 24191 20193 24224
rect 4975 24064 5027 24097
rect 4975 24030 4983 24064
rect 5017 24030 5027 24064
rect 4975 23987 5027 24030
rect 5145 24064 5197 24097
rect 5145 24030 5155 24064
rect 5189 24030 5197 24064
rect 5145 23987 5197 24030
rect 5435 24066 5487 24097
rect 5435 24032 5443 24066
rect 5477 24032 5487 24066
rect 5435 23987 5487 24032
rect 6433 24066 6485 24097
rect 6433 24032 6443 24066
rect 6477 24032 6485 24066
rect 6433 23987 6485 24032
rect 6539 24066 6591 24097
rect 6539 24032 6547 24066
rect 6581 24032 6591 24066
rect 6539 23987 6591 24032
rect 7537 24066 7589 24097
rect 7537 24032 7547 24066
rect 7581 24032 7589 24066
rect 7537 23987 7589 24032
rect 7643 24066 7695 24097
rect 7643 24032 7651 24066
rect 7685 24032 7695 24066
rect 7643 23987 7695 24032
rect 8641 24066 8693 24097
rect 8641 24032 8651 24066
rect 8685 24032 8693 24066
rect 8641 23987 8693 24032
rect 8747 24066 8799 24097
rect 8747 24032 8755 24066
rect 8789 24032 8799 24066
rect 8747 23987 8799 24032
rect 9745 24066 9797 24097
rect 9745 24032 9755 24066
rect 9789 24032 9797 24066
rect 9745 23987 9797 24032
rect 10035 24066 10087 24097
rect 10035 24032 10043 24066
rect 10077 24032 10087 24066
rect 10035 23987 10087 24032
rect 10481 24066 10533 24097
rect 10481 24032 10491 24066
rect 10525 24032 10533 24066
rect 10481 23987 10533 24032
rect 10587 24066 10639 24097
rect 10587 24032 10595 24066
rect 10629 24032 10639 24066
rect 10587 23987 10639 24032
rect 11585 24066 11637 24097
rect 11585 24032 11595 24066
rect 11629 24032 11637 24066
rect 11585 23987 11637 24032
rect 11691 24066 11743 24097
rect 11691 24032 11699 24066
rect 11733 24032 11743 24066
rect 11691 23987 11743 24032
rect 12689 24066 12741 24097
rect 12689 24032 12699 24066
rect 12733 24032 12741 24066
rect 12689 23987 12741 24032
rect 12795 24066 12847 24097
rect 12795 24032 12803 24066
rect 12837 24032 12847 24066
rect 12795 23987 12847 24032
rect 13793 24066 13845 24097
rect 13793 24032 13803 24066
rect 13837 24032 13845 24066
rect 13793 23987 13845 24032
rect 13899 24066 13951 24097
rect 13899 24032 13907 24066
rect 13941 24032 13951 24066
rect 13899 23987 13951 24032
rect 14897 24066 14949 24097
rect 14897 24032 14907 24066
rect 14941 24032 14949 24066
rect 14897 23987 14949 24032
rect 15187 24059 15239 24097
rect 15187 24025 15195 24059
rect 15229 24025 15239 24059
rect 15187 23987 15239 24025
rect 15449 24059 15501 24097
rect 15449 24025 15459 24059
rect 15493 24025 15501 24059
rect 15449 23987 15501 24025
rect 15555 24066 15607 24097
rect 15555 24032 15563 24066
rect 15597 24032 15607 24066
rect 15555 23987 15607 24032
rect 16553 24066 16605 24097
rect 16553 24032 16563 24066
rect 16597 24032 16605 24066
rect 16553 23987 16605 24032
rect 16659 24066 16711 24097
rect 16659 24032 16667 24066
rect 16701 24032 16711 24066
rect 16659 23987 16711 24032
rect 17657 24066 17709 24097
rect 17657 24032 17667 24066
rect 17701 24032 17709 24066
rect 17657 23987 17709 24032
rect 17763 24066 17815 24097
rect 17763 24032 17771 24066
rect 17805 24032 17815 24066
rect 17763 23987 17815 24032
rect 18761 24066 18813 24097
rect 18761 24032 18771 24066
rect 18805 24032 18813 24066
rect 18761 23987 18813 24032
rect 18867 24066 18919 24097
rect 18867 24032 18875 24066
rect 18909 24032 18919 24066
rect 18867 23987 18919 24032
rect 19865 24066 19917 24097
rect 19865 24032 19875 24066
rect 19909 24032 19917 24066
rect 19865 23987 19917 24032
rect 19971 24064 20023 24097
rect 19971 24030 19979 24064
rect 20013 24030 20023 24064
rect 19971 23987 20023 24030
rect 20141 24064 20193 24097
rect 20141 24030 20151 24064
rect 20185 24030 20193 24064
rect 20141 23987 20193 24030
rect 4975 23170 5027 23213
rect 4975 23136 4983 23170
rect 5017 23136 5027 23170
rect 4975 23103 5027 23136
rect 5145 23170 5197 23213
rect 5145 23136 5155 23170
rect 5189 23136 5197 23170
rect 5145 23103 5197 23136
rect 5435 23168 5487 23213
rect 5435 23134 5443 23168
rect 5477 23134 5487 23168
rect 5435 23103 5487 23134
rect 6065 23168 6117 23213
rect 6065 23134 6075 23168
rect 6109 23134 6117 23168
rect 6065 23103 6117 23134
rect 6171 23168 6223 23213
rect 6171 23134 6179 23168
rect 6213 23134 6223 23168
rect 6171 23103 6223 23134
rect 7169 23168 7221 23213
rect 7169 23134 7179 23168
rect 7213 23134 7221 23168
rect 7169 23103 7221 23134
rect 7459 23168 7511 23213
rect 7459 23134 7467 23168
rect 7501 23134 7511 23168
rect 7459 23103 7511 23134
rect 7905 23168 7957 23213
rect 7905 23134 7915 23168
rect 7949 23134 7957 23168
rect 7905 23103 7957 23134
rect 8011 23168 8063 23213
rect 8011 23134 8019 23168
rect 8053 23134 8063 23168
rect 8011 23103 8063 23134
rect 9009 23168 9061 23213
rect 9009 23134 9019 23168
rect 9053 23134 9061 23168
rect 9009 23103 9061 23134
rect 9115 23168 9167 23213
rect 9115 23134 9123 23168
rect 9157 23134 9167 23168
rect 9115 23103 9167 23134
rect 10113 23168 10165 23213
rect 10113 23134 10123 23168
rect 10157 23134 10165 23168
rect 10113 23103 10165 23134
rect 10219 23168 10271 23213
rect 10219 23134 10227 23168
rect 10261 23134 10271 23168
rect 10219 23103 10271 23134
rect 11217 23168 11269 23213
rect 11217 23134 11227 23168
rect 11261 23134 11269 23168
rect 11217 23103 11269 23134
rect 11323 23168 11375 23213
rect 11323 23134 11331 23168
rect 11365 23134 11375 23168
rect 11323 23103 11375 23134
rect 12321 23168 12373 23213
rect 12321 23134 12331 23168
rect 12365 23134 12373 23168
rect 12321 23103 12373 23134
rect 12611 23168 12663 23213
rect 12611 23134 12619 23168
rect 12653 23134 12663 23168
rect 12611 23103 12663 23134
rect 13057 23168 13109 23213
rect 13057 23134 13067 23168
rect 13101 23134 13109 23168
rect 13057 23103 13109 23134
rect 13163 23168 13215 23213
rect 13163 23134 13171 23168
rect 13205 23134 13215 23168
rect 13163 23103 13215 23134
rect 14161 23168 14213 23213
rect 14161 23134 14171 23168
rect 14205 23134 14213 23168
rect 14161 23103 14213 23134
rect 14267 23168 14319 23213
rect 14267 23134 14275 23168
rect 14309 23134 14319 23168
rect 14267 23103 14319 23134
rect 15265 23168 15317 23213
rect 15265 23134 15275 23168
rect 15309 23134 15317 23168
rect 15265 23103 15317 23134
rect 15371 23168 15423 23213
rect 15371 23134 15379 23168
rect 15413 23134 15423 23168
rect 15371 23103 15423 23134
rect 16369 23168 16421 23213
rect 16369 23134 16379 23168
rect 16413 23134 16421 23168
rect 16369 23103 16421 23134
rect 16475 23168 16527 23213
rect 16475 23134 16483 23168
rect 16517 23134 16527 23168
rect 16475 23103 16527 23134
rect 17473 23168 17525 23213
rect 17473 23134 17483 23168
rect 17517 23134 17525 23168
rect 17473 23103 17525 23134
rect 17763 23168 17815 23213
rect 17763 23134 17771 23168
rect 17805 23134 17815 23168
rect 17763 23103 17815 23134
rect 18761 23168 18813 23213
rect 18761 23134 18771 23168
rect 18805 23134 18813 23168
rect 18761 23103 18813 23134
rect 18867 23168 18919 23213
rect 18867 23134 18875 23168
rect 18909 23134 18919 23168
rect 18867 23103 18919 23134
rect 19865 23168 19917 23213
rect 19865 23134 19875 23168
rect 19909 23134 19917 23168
rect 19865 23103 19917 23134
rect 19971 23170 20023 23213
rect 19971 23136 19979 23170
rect 20013 23136 20023 23170
rect 19971 23103 20023 23136
rect 20141 23170 20193 23213
rect 20141 23136 20151 23170
rect 20185 23136 20193 23170
rect 20141 23103 20193 23136
rect 4975 22976 5027 23009
rect 4975 22942 4983 22976
rect 5017 22942 5027 22976
rect 4975 22899 5027 22942
rect 5145 22976 5197 23009
rect 5145 22942 5155 22976
rect 5189 22942 5197 22976
rect 5145 22899 5197 22942
rect 5435 22978 5487 23009
rect 5435 22944 5443 22978
rect 5477 22944 5487 22978
rect 5435 22899 5487 22944
rect 6433 22978 6485 23009
rect 6433 22944 6443 22978
rect 6477 22944 6485 22978
rect 6433 22899 6485 22944
rect 6539 22978 6591 23009
rect 6539 22944 6547 22978
rect 6581 22944 6591 22978
rect 6539 22899 6591 22944
rect 7537 22978 7589 23009
rect 7537 22944 7547 22978
rect 7581 22944 7589 22978
rect 7537 22899 7589 22944
rect 7643 22978 7695 23009
rect 7643 22944 7651 22978
rect 7685 22944 7695 22978
rect 7643 22899 7695 22944
rect 8641 22978 8693 23009
rect 8641 22944 8651 22978
rect 8685 22944 8693 22978
rect 8641 22899 8693 22944
rect 8747 22978 8799 23009
rect 8747 22944 8755 22978
rect 8789 22944 8799 22978
rect 8747 22899 8799 22944
rect 9745 22978 9797 23009
rect 9745 22944 9755 22978
rect 9789 22944 9797 22978
rect 9745 22899 9797 22944
rect 10035 22978 10087 23009
rect 10035 22944 10043 22978
rect 10077 22944 10087 22978
rect 10035 22899 10087 22944
rect 10481 22978 10533 23009
rect 10481 22944 10491 22978
rect 10525 22944 10533 22978
rect 10481 22899 10533 22944
rect 10587 22978 10639 23009
rect 10587 22944 10595 22978
rect 10629 22944 10639 22978
rect 10587 22899 10639 22944
rect 11585 22978 11637 23009
rect 11585 22944 11595 22978
rect 11629 22944 11637 22978
rect 11585 22899 11637 22944
rect 11691 22978 11743 23009
rect 11691 22944 11699 22978
rect 11733 22944 11743 22978
rect 11691 22899 11743 22944
rect 12689 22978 12741 23009
rect 12689 22944 12699 22978
rect 12733 22944 12741 22978
rect 12689 22899 12741 22944
rect 12795 22978 12847 23009
rect 12795 22944 12803 22978
rect 12837 22944 12847 22978
rect 12795 22899 12847 22944
rect 13793 22978 13845 23009
rect 13793 22944 13803 22978
rect 13837 22944 13845 22978
rect 13793 22899 13845 22944
rect 13899 22978 13951 23009
rect 13899 22944 13907 22978
rect 13941 22944 13951 22978
rect 13899 22899 13951 22944
rect 14897 22978 14949 23009
rect 14897 22944 14907 22978
rect 14941 22944 14949 22978
rect 14897 22899 14949 22944
rect 15187 22971 15239 23009
rect 15187 22937 15195 22971
rect 15229 22937 15239 22971
rect 15187 22899 15239 22937
rect 15449 22971 15501 23009
rect 15449 22937 15459 22971
rect 15493 22937 15501 22971
rect 15449 22899 15501 22937
rect 15555 22978 15607 23009
rect 15555 22944 15563 22978
rect 15597 22944 15607 22978
rect 15555 22899 15607 22944
rect 16553 22978 16605 23009
rect 16553 22944 16563 22978
rect 16597 22944 16605 22978
rect 16553 22899 16605 22944
rect 16659 22978 16711 23009
rect 16659 22944 16667 22978
rect 16701 22944 16711 22978
rect 16659 22899 16711 22944
rect 17657 22978 17709 23009
rect 17657 22944 17667 22978
rect 17701 22944 17709 22978
rect 17657 22899 17709 22944
rect 17763 22978 17815 23009
rect 17763 22944 17771 22978
rect 17805 22944 17815 22978
rect 17763 22899 17815 22944
rect 18761 22978 18813 23009
rect 18761 22944 18771 22978
rect 18805 22944 18813 22978
rect 18761 22899 18813 22944
rect 18867 22978 18919 23009
rect 18867 22944 18875 22978
rect 18909 22944 18919 22978
rect 18867 22899 18919 22944
rect 19865 22978 19917 23009
rect 19865 22944 19875 22978
rect 19909 22944 19917 22978
rect 19865 22899 19917 22944
rect 19971 22976 20023 23009
rect 19971 22942 19979 22976
rect 20013 22942 20023 22976
rect 19971 22899 20023 22942
rect 20141 22976 20193 23009
rect 20141 22942 20151 22976
rect 20185 22942 20193 22976
rect 20141 22899 20193 22942
rect 4975 22082 5027 22125
rect 4975 22048 4983 22082
rect 5017 22048 5027 22082
rect 4975 22015 5027 22048
rect 5145 22082 5197 22125
rect 5145 22048 5155 22082
rect 5189 22048 5197 22082
rect 5145 22015 5197 22048
rect 5435 22080 5487 22125
rect 5435 22046 5443 22080
rect 5477 22046 5487 22080
rect 5435 22015 5487 22046
rect 6065 22080 6117 22125
rect 6065 22046 6075 22080
rect 6109 22046 6117 22080
rect 6065 22015 6117 22046
rect 6171 22080 6223 22125
rect 6171 22046 6179 22080
rect 6213 22046 6223 22080
rect 6171 22015 6223 22046
rect 7169 22080 7221 22125
rect 7169 22046 7179 22080
rect 7213 22046 7221 22080
rect 7169 22015 7221 22046
rect 7459 22080 7511 22125
rect 7459 22046 7467 22080
rect 7501 22046 7511 22080
rect 7459 22015 7511 22046
rect 7905 22080 7957 22125
rect 7905 22046 7915 22080
rect 7949 22046 7957 22080
rect 7905 22015 7957 22046
rect 8011 22080 8063 22125
rect 8011 22046 8019 22080
rect 8053 22046 8063 22080
rect 8011 22015 8063 22046
rect 9009 22080 9061 22125
rect 9009 22046 9019 22080
rect 9053 22046 9061 22080
rect 9009 22015 9061 22046
rect 9115 22080 9167 22125
rect 9115 22046 9123 22080
rect 9157 22046 9167 22080
rect 9115 22015 9167 22046
rect 10113 22080 10165 22125
rect 10113 22046 10123 22080
rect 10157 22046 10165 22080
rect 10113 22015 10165 22046
rect 10219 22080 10271 22125
rect 10219 22046 10227 22080
rect 10261 22046 10271 22080
rect 10219 22015 10271 22046
rect 11217 22080 11269 22125
rect 11217 22046 11227 22080
rect 11261 22046 11269 22080
rect 11217 22015 11269 22046
rect 11323 22080 11375 22125
rect 11323 22046 11331 22080
rect 11365 22046 11375 22080
rect 11323 22015 11375 22046
rect 12321 22080 12373 22125
rect 12321 22046 12331 22080
rect 12365 22046 12373 22080
rect 12321 22015 12373 22046
rect 12611 22080 12663 22125
rect 12611 22046 12619 22080
rect 12653 22046 12663 22080
rect 12611 22015 12663 22046
rect 13057 22080 13109 22125
rect 13057 22046 13067 22080
rect 13101 22046 13109 22080
rect 13057 22015 13109 22046
rect 13163 22080 13215 22125
rect 13163 22046 13171 22080
rect 13205 22046 13215 22080
rect 13163 22015 13215 22046
rect 14161 22080 14213 22125
rect 14161 22046 14171 22080
rect 14205 22046 14213 22080
rect 14161 22015 14213 22046
rect 14267 22080 14319 22125
rect 14267 22046 14275 22080
rect 14309 22046 14319 22080
rect 14267 22015 14319 22046
rect 15265 22080 15317 22125
rect 15265 22046 15275 22080
rect 15309 22046 15317 22080
rect 15265 22015 15317 22046
rect 15371 22080 15423 22125
rect 15371 22046 15379 22080
rect 15413 22046 15423 22080
rect 15371 22015 15423 22046
rect 16369 22080 16421 22125
rect 16369 22046 16379 22080
rect 16413 22046 16421 22080
rect 16369 22015 16421 22046
rect 16475 22080 16527 22125
rect 16475 22046 16483 22080
rect 16517 22046 16527 22080
rect 16475 22015 16527 22046
rect 17473 22080 17525 22125
rect 17473 22046 17483 22080
rect 17517 22046 17525 22080
rect 17473 22015 17525 22046
rect 17763 22080 17815 22125
rect 17763 22046 17771 22080
rect 17805 22046 17815 22080
rect 17763 22015 17815 22046
rect 18761 22080 18813 22125
rect 18761 22046 18771 22080
rect 18805 22046 18813 22080
rect 18761 22015 18813 22046
rect 18867 22080 18919 22125
rect 18867 22046 18875 22080
rect 18909 22046 18919 22080
rect 18867 22015 18919 22046
rect 19865 22080 19917 22125
rect 19865 22046 19875 22080
rect 19909 22046 19917 22080
rect 19865 22015 19917 22046
rect 19971 22082 20023 22125
rect 19971 22048 19979 22082
rect 20013 22048 20023 22082
rect 19971 22015 20023 22048
rect 20141 22082 20193 22125
rect 20141 22048 20151 22082
rect 20185 22048 20193 22082
rect 20141 22015 20193 22048
rect 4975 21888 5027 21921
rect 4975 21854 4983 21888
rect 5017 21854 5027 21888
rect 4975 21811 5027 21854
rect 5145 21888 5197 21921
rect 5145 21854 5155 21888
rect 5189 21854 5197 21888
rect 5145 21811 5197 21854
rect 5435 21890 5487 21921
rect 5435 21856 5443 21890
rect 5477 21856 5487 21890
rect 5435 21811 5487 21856
rect 6433 21890 6485 21921
rect 6433 21856 6443 21890
rect 6477 21856 6485 21890
rect 6433 21811 6485 21856
rect 6539 21890 6591 21921
rect 6539 21856 6547 21890
rect 6581 21856 6591 21890
rect 6539 21811 6591 21856
rect 7537 21890 7589 21921
rect 7537 21856 7547 21890
rect 7581 21856 7589 21890
rect 7537 21811 7589 21856
rect 7643 21890 7695 21921
rect 7643 21856 7651 21890
rect 7685 21856 7695 21890
rect 7643 21811 7695 21856
rect 8641 21890 8693 21921
rect 8641 21856 8651 21890
rect 8685 21856 8693 21890
rect 8641 21811 8693 21856
rect 8747 21890 8799 21921
rect 8747 21856 8755 21890
rect 8789 21856 8799 21890
rect 8747 21811 8799 21856
rect 9745 21890 9797 21921
rect 9745 21856 9755 21890
rect 9789 21856 9797 21890
rect 9745 21811 9797 21856
rect 10035 21890 10087 21921
rect 10035 21856 10043 21890
rect 10077 21856 10087 21890
rect 10035 21811 10087 21856
rect 10481 21890 10533 21921
rect 10481 21856 10491 21890
rect 10525 21856 10533 21890
rect 10481 21811 10533 21856
rect 10587 21890 10639 21921
rect 10587 21856 10595 21890
rect 10629 21856 10639 21890
rect 10587 21811 10639 21856
rect 11585 21890 11637 21921
rect 11585 21856 11595 21890
rect 11629 21856 11637 21890
rect 11585 21811 11637 21856
rect 11691 21890 11743 21921
rect 11691 21856 11699 21890
rect 11733 21856 11743 21890
rect 11691 21811 11743 21856
rect 12689 21890 12741 21921
rect 12689 21856 12699 21890
rect 12733 21856 12741 21890
rect 12689 21811 12741 21856
rect 12795 21890 12847 21921
rect 12795 21856 12803 21890
rect 12837 21856 12847 21890
rect 12795 21811 12847 21856
rect 13793 21890 13845 21921
rect 13793 21856 13803 21890
rect 13837 21856 13845 21890
rect 13793 21811 13845 21856
rect 13899 21890 13951 21921
rect 13899 21856 13907 21890
rect 13941 21856 13951 21890
rect 13899 21811 13951 21856
rect 14897 21890 14949 21921
rect 14897 21856 14907 21890
rect 14941 21856 14949 21890
rect 14897 21811 14949 21856
rect 15187 21883 15239 21921
rect 15187 21849 15195 21883
rect 15229 21849 15239 21883
rect 15187 21811 15239 21849
rect 15449 21883 15501 21921
rect 15449 21849 15459 21883
rect 15493 21849 15501 21883
rect 15449 21811 15501 21849
rect 15555 21890 15607 21921
rect 15555 21856 15563 21890
rect 15597 21856 15607 21890
rect 15555 21811 15607 21856
rect 16553 21890 16605 21921
rect 16553 21856 16563 21890
rect 16597 21856 16605 21890
rect 16553 21811 16605 21856
rect 16659 21890 16711 21921
rect 16659 21856 16667 21890
rect 16701 21856 16711 21890
rect 16659 21811 16711 21856
rect 17657 21890 17709 21921
rect 17657 21856 17667 21890
rect 17701 21856 17709 21890
rect 17657 21811 17709 21856
rect 17763 21890 17815 21921
rect 17763 21856 17771 21890
rect 17805 21856 17815 21890
rect 17763 21811 17815 21856
rect 18761 21890 18813 21921
rect 18761 21856 18771 21890
rect 18805 21856 18813 21890
rect 18761 21811 18813 21856
rect 18867 21890 18919 21921
rect 18867 21856 18875 21890
rect 18909 21856 18919 21890
rect 18867 21811 18919 21856
rect 19865 21890 19917 21921
rect 19865 21856 19875 21890
rect 19909 21856 19917 21890
rect 19865 21811 19917 21856
rect 19971 21888 20023 21921
rect 19971 21854 19979 21888
rect 20013 21854 20023 21888
rect 19971 21811 20023 21854
rect 20141 21888 20193 21921
rect 20141 21854 20151 21888
rect 20185 21854 20193 21888
rect 20141 21811 20193 21854
rect 4975 20994 5027 21037
rect 4975 20960 4983 20994
rect 5017 20960 5027 20994
rect 4975 20927 5027 20960
rect 5145 20994 5197 21037
rect 5145 20960 5155 20994
rect 5189 20960 5197 20994
rect 5145 20927 5197 20960
rect 5435 20992 5487 21037
rect 5435 20958 5443 20992
rect 5477 20958 5487 20992
rect 5435 20927 5487 20958
rect 6065 20992 6117 21037
rect 6065 20958 6075 20992
rect 6109 20958 6117 20992
rect 6065 20927 6117 20958
rect 6171 20992 6223 21037
rect 6171 20958 6179 20992
rect 6213 20958 6223 20992
rect 6171 20927 6223 20958
rect 7169 20992 7221 21037
rect 7169 20958 7179 20992
rect 7213 20958 7221 20992
rect 7169 20927 7221 20958
rect 7459 20992 7511 21037
rect 7459 20958 7467 20992
rect 7501 20958 7511 20992
rect 7459 20927 7511 20958
rect 7905 20992 7957 21037
rect 7905 20958 7915 20992
rect 7949 20958 7957 20992
rect 7905 20927 7957 20958
rect 8011 20992 8063 21037
rect 8011 20958 8019 20992
rect 8053 20958 8063 20992
rect 8011 20927 8063 20958
rect 9009 20992 9061 21037
rect 9009 20958 9019 20992
rect 9053 20958 9061 20992
rect 9009 20927 9061 20958
rect 9115 20992 9167 21037
rect 9115 20958 9123 20992
rect 9157 20958 9167 20992
rect 9115 20927 9167 20958
rect 10113 20992 10165 21037
rect 10113 20958 10123 20992
rect 10157 20958 10165 20992
rect 10113 20927 10165 20958
rect 10219 20992 10271 21037
rect 10219 20958 10227 20992
rect 10261 20958 10271 20992
rect 10219 20927 10271 20958
rect 11217 20992 11269 21037
rect 11217 20958 11227 20992
rect 11261 20958 11269 20992
rect 11217 20927 11269 20958
rect 11323 20992 11375 21037
rect 11323 20958 11331 20992
rect 11365 20958 11375 20992
rect 11323 20927 11375 20958
rect 12321 20992 12373 21037
rect 12321 20958 12331 20992
rect 12365 20958 12373 20992
rect 12321 20927 12373 20958
rect 12611 20992 12663 21037
rect 12611 20958 12619 20992
rect 12653 20958 12663 20992
rect 12611 20927 12663 20958
rect 13057 20992 13109 21037
rect 13057 20958 13067 20992
rect 13101 20958 13109 20992
rect 13057 20927 13109 20958
rect 13163 20992 13215 21037
rect 13163 20958 13171 20992
rect 13205 20958 13215 20992
rect 13163 20927 13215 20958
rect 14161 20992 14213 21037
rect 14161 20958 14171 20992
rect 14205 20958 14213 20992
rect 14161 20927 14213 20958
rect 14267 20992 14319 21037
rect 14267 20958 14275 20992
rect 14309 20958 14319 20992
rect 14267 20927 14319 20958
rect 15265 20992 15317 21037
rect 15265 20958 15275 20992
rect 15309 20958 15317 20992
rect 15265 20927 15317 20958
rect 15371 20992 15423 21037
rect 15371 20958 15379 20992
rect 15413 20958 15423 20992
rect 15371 20927 15423 20958
rect 16369 20992 16421 21037
rect 16369 20958 16379 20992
rect 16413 20958 16421 20992
rect 16369 20927 16421 20958
rect 16475 20992 16527 21037
rect 16475 20958 16483 20992
rect 16517 20958 16527 20992
rect 16475 20927 16527 20958
rect 17473 20992 17525 21037
rect 17473 20958 17483 20992
rect 17517 20958 17525 20992
rect 17473 20927 17525 20958
rect 17763 20992 17815 21037
rect 17763 20958 17771 20992
rect 17805 20958 17815 20992
rect 17763 20927 17815 20958
rect 18761 20992 18813 21037
rect 18761 20958 18771 20992
rect 18805 20958 18813 20992
rect 18761 20927 18813 20958
rect 18867 20992 18919 21037
rect 18867 20958 18875 20992
rect 18909 20958 18919 20992
rect 18867 20927 18919 20958
rect 19865 20992 19917 21037
rect 19865 20958 19875 20992
rect 19909 20958 19917 20992
rect 19865 20927 19917 20958
rect 19971 20994 20023 21037
rect 19971 20960 19979 20994
rect 20013 20960 20023 20994
rect 19971 20927 20023 20960
rect 20141 20994 20193 21037
rect 20141 20960 20151 20994
rect 20185 20960 20193 20994
rect 20141 20927 20193 20960
rect 4975 20800 5027 20833
rect 4975 20766 4983 20800
rect 5017 20766 5027 20800
rect 4975 20723 5027 20766
rect 5145 20800 5197 20833
rect 5145 20766 5155 20800
rect 5189 20766 5197 20800
rect 5145 20723 5197 20766
rect 5435 20802 5487 20833
rect 5435 20768 5443 20802
rect 5477 20768 5487 20802
rect 5435 20723 5487 20768
rect 6433 20802 6485 20833
rect 6433 20768 6443 20802
rect 6477 20768 6485 20802
rect 6433 20723 6485 20768
rect 6539 20802 6591 20833
rect 6539 20768 6547 20802
rect 6581 20768 6591 20802
rect 6539 20723 6591 20768
rect 7537 20802 7589 20833
rect 7537 20768 7547 20802
rect 7581 20768 7589 20802
rect 7537 20723 7589 20768
rect 7643 20802 7695 20833
rect 7643 20768 7651 20802
rect 7685 20768 7695 20802
rect 7643 20723 7695 20768
rect 8641 20802 8693 20833
rect 8641 20768 8651 20802
rect 8685 20768 8693 20802
rect 8641 20723 8693 20768
rect 8747 20802 8799 20833
rect 8747 20768 8755 20802
rect 8789 20768 8799 20802
rect 8747 20723 8799 20768
rect 9745 20802 9797 20833
rect 9745 20768 9755 20802
rect 9789 20768 9797 20802
rect 9745 20723 9797 20768
rect 10035 20802 10087 20833
rect 10035 20768 10043 20802
rect 10077 20768 10087 20802
rect 10035 20723 10087 20768
rect 10481 20802 10533 20833
rect 10481 20768 10491 20802
rect 10525 20768 10533 20802
rect 10481 20723 10533 20768
rect 10587 20802 10639 20833
rect 10587 20768 10595 20802
rect 10629 20768 10639 20802
rect 10587 20723 10639 20768
rect 11585 20802 11637 20833
rect 11585 20768 11595 20802
rect 11629 20768 11637 20802
rect 11585 20723 11637 20768
rect 11691 20802 11743 20833
rect 11691 20768 11699 20802
rect 11733 20768 11743 20802
rect 11691 20723 11743 20768
rect 12689 20802 12741 20833
rect 12689 20768 12699 20802
rect 12733 20768 12741 20802
rect 12689 20723 12741 20768
rect 12795 20802 12847 20833
rect 12795 20768 12803 20802
rect 12837 20768 12847 20802
rect 12795 20723 12847 20768
rect 13793 20802 13845 20833
rect 13793 20768 13803 20802
rect 13837 20768 13845 20802
rect 13793 20723 13845 20768
rect 13899 20802 13951 20833
rect 13899 20768 13907 20802
rect 13941 20768 13951 20802
rect 13899 20723 13951 20768
rect 14897 20802 14949 20833
rect 14897 20768 14907 20802
rect 14941 20768 14949 20802
rect 14897 20723 14949 20768
rect 15187 20795 15239 20833
rect 15187 20761 15195 20795
rect 15229 20761 15239 20795
rect 15187 20723 15239 20761
rect 15449 20795 15501 20833
rect 15449 20761 15459 20795
rect 15493 20761 15501 20795
rect 15449 20723 15501 20761
rect 15555 20802 15607 20833
rect 15555 20768 15563 20802
rect 15597 20768 15607 20802
rect 15555 20723 15607 20768
rect 16553 20802 16605 20833
rect 16553 20768 16563 20802
rect 16597 20768 16605 20802
rect 16553 20723 16605 20768
rect 16659 20802 16711 20833
rect 16659 20768 16667 20802
rect 16701 20768 16711 20802
rect 16659 20723 16711 20768
rect 17657 20802 17709 20833
rect 17657 20768 17667 20802
rect 17701 20768 17709 20802
rect 17657 20723 17709 20768
rect 17763 20802 17815 20833
rect 17763 20768 17771 20802
rect 17805 20768 17815 20802
rect 17763 20723 17815 20768
rect 18761 20802 18813 20833
rect 18761 20768 18771 20802
rect 18805 20768 18813 20802
rect 18761 20723 18813 20768
rect 18867 20802 18919 20833
rect 18867 20768 18875 20802
rect 18909 20768 18919 20802
rect 18867 20723 18919 20768
rect 19865 20802 19917 20833
rect 19865 20768 19875 20802
rect 19909 20768 19917 20802
rect 19865 20723 19917 20768
rect 19971 20800 20023 20833
rect 19971 20766 19979 20800
rect 20013 20766 20023 20800
rect 19971 20723 20023 20766
rect 20141 20800 20193 20833
rect 20141 20766 20151 20800
rect 20185 20766 20193 20800
rect 20141 20723 20193 20766
rect 4975 19906 5027 19949
rect 4975 19872 4983 19906
rect 5017 19872 5027 19906
rect 4975 19839 5027 19872
rect 5145 19906 5197 19949
rect 5145 19872 5155 19906
rect 5189 19872 5197 19906
rect 5145 19839 5197 19872
rect 5435 19904 5487 19949
rect 5435 19870 5443 19904
rect 5477 19870 5487 19904
rect 5435 19839 5487 19870
rect 6065 19904 6117 19949
rect 6065 19870 6075 19904
rect 6109 19870 6117 19904
rect 6065 19839 6117 19870
rect 6171 19904 6223 19949
rect 6171 19870 6179 19904
rect 6213 19870 6223 19904
rect 6171 19839 6223 19870
rect 7169 19904 7221 19949
rect 7169 19870 7179 19904
rect 7213 19870 7221 19904
rect 7169 19839 7221 19870
rect 7459 19904 7511 19949
rect 7459 19870 7467 19904
rect 7501 19870 7511 19904
rect 7459 19839 7511 19870
rect 7905 19904 7957 19949
rect 7905 19870 7915 19904
rect 7949 19870 7957 19904
rect 7905 19839 7957 19870
rect 8011 19904 8063 19949
rect 8011 19870 8019 19904
rect 8053 19870 8063 19904
rect 8011 19839 8063 19870
rect 9009 19904 9061 19949
rect 9009 19870 9019 19904
rect 9053 19870 9061 19904
rect 9009 19839 9061 19870
rect 9115 19904 9167 19949
rect 9115 19870 9123 19904
rect 9157 19870 9167 19904
rect 9115 19839 9167 19870
rect 10113 19904 10165 19949
rect 10113 19870 10123 19904
rect 10157 19870 10165 19904
rect 10113 19839 10165 19870
rect 10219 19904 10271 19949
rect 10219 19870 10227 19904
rect 10261 19870 10271 19904
rect 10219 19839 10271 19870
rect 11217 19904 11269 19949
rect 11217 19870 11227 19904
rect 11261 19870 11269 19904
rect 11217 19839 11269 19870
rect 11323 19904 11375 19949
rect 11323 19870 11331 19904
rect 11365 19870 11375 19904
rect 11323 19839 11375 19870
rect 12321 19904 12373 19949
rect 12321 19870 12331 19904
rect 12365 19870 12373 19904
rect 12321 19839 12373 19870
rect 12611 19904 12663 19949
rect 12611 19870 12619 19904
rect 12653 19870 12663 19904
rect 12611 19839 12663 19870
rect 13057 19904 13109 19949
rect 13057 19870 13067 19904
rect 13101 19870 13109 19904
rect 13057 19839 13109 19870
rect 13163 19904 13215 19949
rect 13163 19870 13171 19904
rect 13205 19870 13215 19904
rect 13163 19839 13215 19870
rect 14161 19904 14213 19949
rect 14161 19870 14171 19904
rect 14205 19870 14213 19904
rect 14161 19839 14213 19870
rect 14267 19904 14319 19949
rect 14267 19870 14275 19904
rect 14309 19870 14319 19904
rect 14267 19839 14319 19870
rect 15265 19904 15317 19949
rect 15265 19870 15275 19904
rect 15309 19870 15317 19904
rect 15265 19839 15317 19870
rect 15371 19904 15423 19949
rect 15371 19870 15379 19904
rect 15413 19870 15423 19904
rect 15371 19839 15423 19870
rect 16369 19904 16421 19949
rect 16369 19870 16379 19904
rect 16413 19870 16421 19904
rect 16369 19839 16421 19870
rect 16475 19904 16527 19949
rect 16475 19870 16483 19904
rect 16517 19870 16527 19904
rect 16475 19839 16527 19870
rect 17473 19904 17525 19949
rect 17473 19870 17483 19904
rect 17517 19870 17525 19904
rect 17473 19839 17525 19870
rect 17763 19904 17815 19949
rect 17763 19870 17771 19904
rect 17805 19870 17815 19904
rect 17763 19839 17815 19870
rect 18761 19904 18813 19949
rect 18761 19870 18771 19904
rect 18805 19870 18813 19904
rect 18761 19839 18813 19870
rect 18867 19904 18919 19949
rect 18867 19870 18875 19904
rect 18909 19870 18919 19904
rect 18867 19839 18919 19870
rect 19865 19904 19917 19949
rect 19865 19870 19875 19904
rect 19909 19870 19917 19904
rect 19865 19839 19917 19870
rect 19971 19906 20023 19949
rect 19971 19872 19979 19906
rect 20013 19872 20023 19906
rect 19971 19839 20023 19872
rect 20141 19906 20193 19949
rect 20141 19872 20151 19906
rect 20185 19872 20193 19906
rect 20141 19839 20193 19872
rect 4975 19712 5027 19745
rect 4975 19678 4983 19712
rect 5017 19678 5027 19712
rect 4975 19635 5027 19678
rect 5145 19712 5197 19745
rect 5145 19678 5155 19712
rect 5189 19678 5197 19712
rect 5145 19635 5197 19678
rect 5435 19714 5487 19745
rect 5435 19680 5443 19714
rect 5477 19680 5487 19714
rect 5435 19635 5487 19680
rect 6433 19714 6485 19745
rect 6433 19680 6443 19714
rect 6477 19680 6485 19714
rect 6433 19635 6485 19680
rect 6539 19714 6591 19745
rect 6539 19680 6547 19714
rect 6581 19680 6591 19714
rect 6539 19635 6591 19680
rect 7537 19714 7589 19745
rect 7537 19680 7547 19714
rect 7581 19680 7589 19714
rect 7537 19635 7589 19680
rect 7643 19714 7695 19745
rect 7643 19680 7651 19714
rect 7685 19680 7695 19714
rect 7643 19635 7695 19680
rect 8641 19714 8693 19745
rect 8641 19680 8651 19714
rect 8685 19680 8693 19714
rect 8641 19635 8693 19680
rect 8747 19714 8799 19745
rect 8747 19680 8755 19714
rect 8789 19680 8799 19714
rect 8747 19635 8799 19680
rect 9745 19714 9797 19745
rect 9745 19680 9755 19714
rect 9789 19680 9797 19714
rect 9745 19635 9797 19680
rect 10035 19714 10087 19745
rect 10035 19680 10043 19714
rect 10077 19680 10087 19714
rect 10035 19635 10087 19680
rect 10481 19714 10533 19745
rect 10481 19680 10491 19714
rect 10525 19680 10533 19714
rect 10481 19635 10533 19680
rect 10587 19714 10639 19745
rect 10587 19680 10595 19714
rect 10629 19680 10639 19714
rect 10587 19635 10639 19680
rect 11585 19714 11637 19745
rect 11585 19680 11595 19714
rect 11629 19680 11637 19714
rect 11585 19635 11637 19680
rect 11691 19714 11743 19745
rect 11691 19680 11699 19714
rect 11733 19680 11743 19714
rect 11691 19635 11743 19680
rect 12689 19714 12741 19745
rect 12689 19680 12699 19714
rect 12733 19680 12741 19714
rect 12689 19635 12741 19680
rect 12795 19714 12847 19745
rect 12795 19680 12803 19714
rect 12837 19680 12847 19714
rect 12795 19635 12847 19680
rect 13793 19714 13845 19745
rect 13793 19680 13803 19714
rect 13837 19680 13845 19714
rect 13793 19635 13845 19680
rect 13899 19714 13951 19745
rect 13899 19680 13907 19714
rect 13941 19680 13951 19714
rect 13899 19635 13951 19680
rect 14897 19714 14949 19745
rect 14897 19680 14907 19714
rect 14941 19680 14949 19714
rect 14897 19635 14949 19680
rect 15187 19707 15239 19745
rect 15187 19673 15195 19707
rect 15229 19673 15239 19707
rect 15187 19635 15239 19673
rect 15449 19707 15501 19745
rect 15449 19673 15459 19707
rect 15493 19673 15501 19707
rect 15449 19635 15501 19673
rect 15555 19714 15607 19745
rect 15555 19680 15563 19714
rect 15597 19680 15607 19714
rect 15555 19635 15607 19680
rect 16553 19714 16605 19745
rect 16553 19680 16563 19714
rect 16597 19680 16605 19714
rect 16553 19635 16605 19680
rect 16659 19714 16711 19745
rect 16659 19680 16667 19714
rect 16701 19680 16711 19714
rect 16659 19635 16711 19680
rect 17657 19714 17709 19745
rect 17657 19680 17667 19714
rect 17701 19680 17709 19714
rect 17657 19635 17709 19680
rect 17763 19714 17815 19745
rect 17763 19680 17771 19714
rect 17805 19680 17815 19714
rect 17763 19635 17815 19680
rect 18761 19714 18813 19745
rect 18761 19680 18771 19714
rect 18805 19680 18813 19714
rect 18761 19635 18813 19680
rect 18867 19714 18919 19745
rect 18867 19680 18875 19714
rect 18909 19680 18919 19714
rect 18867 19635 18919 19680
rect 19865 19714 19917 19745
rect 19865 19680 19875 19714
rect 19909 19680 19917 19714
rect 19865 19635 19917 19680
rect 19971 19712 20023 19745
rect 19971 19678 19979 19712
rect 20013 19678 20023 19712
rect 19971 19635 20023 19678
rect 20141 19712 20193 19745
rect 20141 19678 20151 19712
rect 20185 19678 20193 19712
rect 20141 19635 20193 19678
rect 4975 18818 5027 18861
rect 4975 18784 4983 18818
rect 5017 18784 5027 18818
rect 4975 18751 5027 18784
rect 5145 18818 5197 18861
rect 5145 18784 5155 18818
rect 5189 18784 5197 18818
rect 5145 18751 5197 18784
rect 5435 18816 5487 18861
rect 5435 18782 5443 18816
rect 5477 18782 5487 18816
rect 5435 18751 5487 18782
rect 6065 18816 6117 18861
rect 6065 18782 6075 18816
rect 6109 18782 6117 18816
rect 6065 18751 6117 18782
rect 6171 18816 6223 18861
rect 6171 18782 6179 18816
rect 6213 18782 6223 18816
rect 6171 18751 6223 18782
rect 7169 18816 7221 18861
rect 7169 18782 7179 18816
rect 7213 18782 7221 18816
rect 7169 18751 7221 18782
rect 7459 18816 7511 18861
rect 7459 18782 7467 18816
rect 7501 18782 7511 18816
rect 7459 18751 7511 18782
rect 7905 18816 7957 18861
rect 7905 18782 7915 18816
rect 7949 18782 7957 18816
rect 7905 18751 7957 18782
rect 8011 18816 8063 18861
rect 8011 18782 8019 18816
rect 8053 18782 8063 18816
rect 8011 18751 8063 18782
rect 9009 18816 9061 18861
rect 9009 18782 9019 18816
rect 9053 18782 9061 18816
rect 9009 18751 9061 18782
rect 9115 18816 9167 18861
rect 9115 18782 9123 18816
rect 9157 18782 9167 18816
rect 9115 18751 9167 18782
rect 10113 18816 10165 18861
rect 10113 18782 10123 18816
rect 10157 18782 10165 18816
rect 10113 18751 10165 18782
rect 10219 18816 10271 18861
rect 10219 18782 10227 18816
rect 10261 18782 10271 18816
rect 10219 18751 10271 18782
rect 11217 18816 11269 18861
rect 11217 18782 11227 18816
rect 11261 18782 11269 18816
rect 11217 18751 11269 18782
rect 11323 18816 11375 18861
rect 11323 18782 11331 18816
rect 11365 18782 11375 18816
rect 11323 18751 11375 18782
rect 12321 18816 12373 18861
rect 12321 18782 12331 18816
rect 12365 18782 12373 18816
rect 12321 18751 12373 18782
rect 12611 18816 12663 18861
rect 12611 18782 12619 18816
rect 12653 18782 12663 18816
rect 12611 18751 12663 18782
rect 13057 18816 13109 18861
rect 13057 18782 13067 18816
rect 13101 18782 13109 18816
rect 13057 18751 13109 18782
rect 13163 18816 13215 18861
rect 13163 18782 13171 18816
rect 13205 18782 13215 18816
rect 13163 18751 13215 18782
rect 14161 18816 14213 18861
rect 14161 18782 14171 18816
rect 14205 18782 14213 18816
rect 14161 18751 14213 18782
rect 14267 18816 14319 18861
rect 14267 18782 14275 18816
rect 14309 18782 14319 18816
rect 14267 18751 14319 18782
rect 15265 18816 15317 18861
rect 15265 18782 15275 18816
rect 15309 18782 15317 18816
rect 15265 18751 15317 18782
rect 15371 18816 15423 18861
rect 15371 18782 15379 18816
rect 15413 18782 15423 18816
rect 15371 18751 15423 18782
rect 16369 18816 16421 18861
rect 16369 18782 16379 18816
rect 16413 18782 16421 18816
rect 16369 18751 16421 18782
rect 16475 18816 16527 18861
rect 16475 18782 16483 18816
rect 16517 18782 16527 18816
rect 16475 18751 16527 18782
rect 17473 18816 17525 18861
rect 17473 18782 17483 18816
rect 17517 18782 17525 18816
rect 17473 18751 17525 18782
rect 17763 18816 17815 18861
rect 17763 18782 17771 18816
rect 17805 18782 17815 18816
rect 17763 18751 17815 18782
rect 18761 18816 18813 18861
rect 18761 18782 18771 18816
rect 18805 18782 18813 18816
rect 18761 18751 18813 18782
rect 18867 18816 18919 18861
rect 18867 18782 18875 18816
rect 18909 18782 18919 18816
rect 18867 18751 18919 18782
rect 19865 18816 19917 18861
rect 19865 18782 19875 18816
rect 19909 18782 19917 18816
rect 19865 18751 19917 18782
rect 19971 18818 20023 18861
rect 19971 18784 19979 18818
rect 20013 18784 20023 18818
rect 19971 18751 20023 18784
rect 20141 18818 20193 18861
rect 20141 18784 20151 18818
rect 20185 18784 20193 18818
rect 20141 18751 20193 18784
rect 4975 18624 5027 18657
rect 4975 18590 4983 18624
rect 5017 18590 5027 18624
rect 4975 18547 5027 18590
rect 5145 18624 5197 18657
rect 5145 18590 5155 18624
rect 5189 18590 5197 18624
rect 5145 18547 5197 18590
rect 5435 18626 5487 18657
rect 5435 18592 5443 18626
rect 5477 18592 5487 18626
rect 5435 18547 5487 18592
rect 6433 18626 6485 18657
rect 6433 18592 6443 18626
rect 6477 18592 6485 18626
rect 6433 18547 6485 18592
rect 6539 18626 6591 18657
rect 6539 18592 6547 18626
rect 6581 18592 6591 18626
rect 6539 18547 6591 18592
rect 7537 18626 7589 18657
rect 7537 18592 7547 18626
rect 7581 18592 7589 18626
rect 7537 18547 7589 18592
rect 7643 18626 7695 18657
rect 7643 18592 7651 18626
rect 7685 18592 7695 18626
rect 7643 18547 7695 18592
rect 8641 18626 8693 18657
rect 8641 18592 8651 18626
rect 8685 18592 8693 18626
rect 8641 18547 8693 18592
rect 8747 18626 8799 18657
rect 8747 18592 8755 18626
rect 8789 18592 8799 18626
rect 8747 18547 8799 18592
rect 9745 18626 9797 18657
rect 9745 18592 9755 18626
rect 9789 18592 9797 18626
rect 9745 18547 9797 18592
rect 10035 18626 10087 18657
rect 10035 18592 10043 18626
rect 10077 18592 10087 18626
rect 10035 18547 10087 18592
rect 10481 18626 10533 18657
rect 10481 18592 10491 18626
rect 10525 18592 10533 18626
rect 10481 18547 10533 18592
rect 10587 18626 10639 18657
rect 10587 18592 10595 18626
rect 10629 18592 10639 18626
rect 10587 18547 10639 18592
rect 11585 18626 11637 18657
rect 11585 18592 11595 18626
rect 11629 18592 11637 18626
rect 11585 18547 11637 18592
rect 11691 18626 11743 18657
rect 11691 18592 11699 18626
rect 11733 18592 11743 18626
rect 11691 18547 11743 18592
rect 12689 18626 12741 18657
rect 12689 18592 12699 18626
rect 12733 18592 12741 18626
rect 12689 18547 12741 18592
rect 12795 18626 12847 18657
rect 12795 18592 12803 18626
rect 12837 18592 12847 18626
rect 12795 18547 12847 18592
rect 13793 18626 13845 18657
rect 13793 18592 13803 18626
rect 13837 18592 13845 18626
rect 13793 18547 13845 18592
rect 13899 18626 13951 18657
rect 13899 18592 13907 18626
rect 13941 18592 13951 18626
rect 13899 18547 13951 18592
rect 14897 18626 14949 18657
rect 14897 18592 14907 18626
rect 14941 18592 14949 18626
rect 14897 18547 14949 18592
rect 15187 18619 15239 18657
rect 15187 18585 15195 18619
rect 15229 18585 15239 18619
rect 15187 18547 15239 18585
rect 15449 18619 15501 18657
rect 15449 18585 15459 18619
rect 15493 18585 15501 18619
rect 15449 18547 15501 18585
rect 15555 18626 15607 18657
rect 15555 18592 15563 18626
rect 15597 18592 15607 18626
rect 15555 18547 15607 18592
rect 16553 18626 16605 18657
rect 16553 18592 16563 18626
rect 16597 18592 16605 18626
rect 16553 18547 16605 18592
rect 16659 18626 16711 18657
rect 16659 18592 16667 18626
rect 16701 18592 16711 18626
rect 16659 18547 16711 18592
rect 17657 18626 17709 18657
rect 17657 18592 17667 18626
rect 17701 18592 17709 18626
rect 17657 18547 17709 18592
rect 17763 18626 17815 18657
rect 17763 18592 17771 18626
rect 17805 18592 17815 18626
rect 17763 18547 17815 18592
rect 18761 18626 18813 18657
rect 18761 18592 18771 18626
rect 18805 18592 18813 18626
rect 18761 18547 18813 18592
rect 18867 18626 18919 18657
rect 18867 18592 18875 18626
rect 18909 18592 18919 18626
rect 18867 18547 18919 18592
rect 19865 18626 19917 18657
rect 19865 18592 19875 18626
rect 19909 18592 19917 18626
rect 19865 18547 19917 18592
rect 19971 18624 20023 18657
rect 19971 18590 19979 18624
rect 20013 18590 20023 18624
rect 19971 18547 20023 18590
rect 20141 18624 20193 18657
rect 20141 18590 20151 18624
rect 20185 18590 20193 18624
rect 20141 18547 20193 18590
rect 4975 17730 5027 17773
rect 4975 17696 4983 17730
rect 5017 17696 5027 17730
rect 4975 17663 5027 17696
rect 5145 17730 5197 17773
rect 5145 17696 5155 17730
rect 5189 17696 5197 17730
rect 5145 17663 5197 17696
rect 5435 17728 5487 17773
rect 5435 17694 5443 17728
rect 5477 17694 5487 17728
rect 5435 17663 5487 17694
rect 6065 17728 6117 17773
rect 6065 17694 6075 17728
rect 6109 17694 6117 17728
rect 6065 17663 6117 17694
rect 6171 17728 6223 17773
rect 6171 17694 6179 17728
rect 6213 17694 6223 17728
rect 6171 17663 6223 17694
rect 7169 17728 7221 17773
rect 7169 17694 7179 17728
rect 7213 17694 7221 17728
rect 7169 17663 7221 17694
rect 7459 17728 7511 17773
rect 7459 17694 7467 17728
rect 7501 17694 7511 17728
rect 7459 17663 7511 17694
rect 7905 17728 7957 17773
rect 7905 17694 7915 17728
rect 7949 17694 7957 17728
rect 7905 17663 7957 17694
rect 8011 17728 8063 17773
rect 8011 17694 8019 17728
rect 8053 17694 8063 17728
rect 8011 17663 8063 17694
rect 9009 17728 9061 17773
rect 9009 17694 9019 17728
rect 9053 17694 9061 17728
rect 9009 17663 9061 17694
rect 9115 17728 9167 17773
rect 9115 17694 9123 17728
rect 9157 17694 9167 17728
rect 9115 17663 9167 17694
rect 10113 17728 10165 17773
rect 10113 17694 10123 17728
rect 10157 17694 10165 17728
rect 10113 17663 10165 17694
rect 10219 17728 10271 17773
rect 10219 17694 10227 17728
rect 10261 17694 10271 17728
rect 10219 17663 10271 17694
rect 11217 17728 11269 17773
rect 11217 17694 11227 17728
rect 11261 17694 11269 17728
rect 11217 17663 11269 17694
rect 11323 17728 11375 17773
rect 11323 17694 11331 17728
rect 11365 17694 11375 17728
rect 11323 17663 11375 17694
rect 12321 17728 12373 17773
rect 12321 17694 12331 17728
rect 12365 17694 12373 17728
rect 12321 17663 12373 17694
rect 12611 17728 12663 17773
rect 12611 17694 12619 17728
rect 12653 17694 12663 17728
rect 12611 17663 12663 17694
rect 13057 17728 13109 17773
rect 13057 17694 13067 17728
rect 13101 17694 13109 17728
rect 13057 17663 13109 17694
rect 13163 17728 13215 17773
rect 13163 17694 13171 17728
rect 13205 17694 13215 17728
rect 13163 17663 13215 17694
rect 14161 17728 14213 17773
rect 14161 17694 14171 17728
rect 14205 17694 14213 17728
rect 14161 17663 14213 17694
rect 14267 17728 14319 17773
rect 14267 17694 14275 17728
rect 14309 17694 14319 17728
rect 14267 17663 14319 17694
rect 15265 17728 15317 17773
rect 15265 17694 15275 17728
rect 15309 17694 15317 17728
rect 15265 17663 15317 17694
rect 15371 17728 15423 17773
rect 15371 17694 15379 17728
rect 15413 17694 15423 17728
rect 15371 17663 15423 17694
rect 16369 17728 16421 17773
rect 16369 17694 16379 17728
rect 16413 17694 16421 17728
rect 16369 17663 16421 17694
rect 16475 17728 16527 17773
rect 16475 17694 16483 17728
rect 16517 17694 16527 17728
rect 16475 17663 16527 17694
rect 17473 17728 17525 17773
rect 17473 17694 17483 17728
rect 17517 17694 17525 17728
rect 17473 17663 17525 17694
rect 17763 17728 17815 17773
rect 17763 17694 17771 17728
rect 17805 17694 17815 17728
rect 17763 17663 17815 17694
rect 18761 17728 18813 17773
rect 18761 17694 18771 17728
rect 18805 17694 18813 17728
rect 18761 17663 18813 17694
rect 18867 17728 18919 17773
rect 18867 17694 18875 17728
rect 18909 17694 18919 17728
rect 18867 17663 18919 17694
rect 19865 17728 19917 17773
rect 19865 17694 19875 17728
rect 19909 17694 19917 17728
rect 19865 17663 19917 17694
rect 19971 17730 20023 17773
rect 19971 17696 19979 17730
rect 20013 17696 20023 17730
rect 19971 17663 20023 17696
rect 20141 17730 20193 17773
rect 20141 17696 20151 17730
rect 20185 17696 20193 17730
rect 20141 17663 20193 17696
rect 4975 17536 5027 17569
rect 4975 17502 4983 17536
rect 5017 17502 5027 17536
rect 4975 17459 5027 17502
rect 5145 17536 5197 17569
rect 5145 17502 5155 17536
rect 5189 17502 5197 17536
rect 5145 17459 5197 17502
rect 5435 17538 5487 17569
rect 5435 17504 5443 17538
rect 5477 17504 5487 17538
rect 5435 17459 5487 17504
rect 6433 17538 6485 17569
rect 6433 17504 6443 17538
rect 6477 17504 6485 17538
rect 6433 17459 6485 17504
rect 6539 17538 6591 17569
rect 6539 17504 6547 17538
rect 6581 17504 6591 17538
rect 6539 17459 6591 17504
rect 7537 17538 7589 17569
rect 7537 17504 7547 17538
rect 7581 17504 7589 17538
rect 7537 17459 7589 17504
rect 7643 17538 7695 17569
rect 7643 17504 7651 17538
rect 7685 17504 7695 17538
rect 7643 17459 7695 17504
rect 8641 17538 8693 17569
rect 8641 17504 8651 17538
rect 8685 17504 8693 17538
rect 8641 17459 8693 17504
rect 8747 17538 8799 17569
rect 8747 17504 8755 17538
rect 8789 17504 8799 17538
rect 8747 17459 8799 17504
rect 9745 17538 9797 17569
rect 9745 17504 9755 17538
rect 9789 17504 9797 17538
rect 9745 17459 9797 17504
rect 10035 17538 10087 17569
rect 10035 17504 10043 17538
rect 10077 17504 10087 17538
rect 10035 17459 10087 17504
rect 10481 17538 10533 17569
rect 10481 17504 10491 17538
rect 10525 17504 10533 17538
rect 10481 17459 10533 17504
rect 10587 17538 10639 17569
rect 10587 17504 10595 17538
rect 10629 17504 10639 17538
rect 10587 17459 10639 17504
rect 11585 17538 11637 17569
rect 11585 17504 11595 17538
rect 11629 17504 11637 17538
rect 11585 17459 11637 17504
rect 11691 17538 11743 17569
rect 11691 17504 11699 17538
rect 11733 17504 11743 17538
rect 11691 17459 11743 17504
rect 12689 17538 12741 17569
rect 12689 17504 12699 17538
rect 12733 17504 12741 17538
rect 12689 17459 12741 17504
rect 12795 17538 12847 17569
rect 12795 17504 12803 17538
rect 12837 17504 12847 17538
rect 12795 17459 12847 17504
rect 13793 17538 13845 17569
rect 13793 17504 13803 17538
rect 13837 17504 13845 17538
rect 13793 17459 13845 17504
rect 13899 17538 13951 17569
rect 13899 17504 13907 17538
rect 13941 17504 13951 17538
rect 13899 17459 13951 17504
rect 14897 17538 14949 17569
rect 14897 17504 14907 17538
rect 14941 17504 14949 17538
rect 14897 17459 14949 17504
rect 15187 17531 15239 17569
rect 15187 17497 15195 17531
rect 15229 17497 15239 17531
rect 15187 17459 15239 17497
rect 15449 17531 15501 17569
rect 15449 17497 15459 17531
rect 15493 17497 15501 17531
rect 15449 17459 15501 17497
rect 15555 17538 15607 17569
rect 15555 17504 15563 17538
rect 15597 17504 15607 17538
rect 15555 17459 15607 17504
rect 16553 17538 16605 17569
rect 16553 17504 16563 17538
rect 16597 17504 16605 17538
rect 16553 17459 16605 17504
rect 16659 17538 16711 17569
rect 16659 17504 16667 17538
rect 16701 17504 16711 17538
rect 16659 17459 16711 17504
rect 17657 17538 17709 17569
rect 17657 17504 17667 17538
rect 17701 17504 17709 17538
rect 17657 17459 17709 17504
rect 17763 17538 17815 17569
rect 17763 17504 17771 17538
rect 17805 17504 17815 17538
rect 17763 17459 17815 17504
rect 18761 17538 18813 17569
rect 18761 17504 18771 17538
rect 18805 17504 18813 17538
rect 18761 17459 18813 17504
rect 18867 17538 18919 17569
rect 18867 17504 18875 17538
rect 18909 17504 18919 17538
rect 18867 17459 18919 17504
rect 19865 17538 19917 17569
rect 19865 17504 19875 17538
rect 19909 17504 19917 17538
rect 19865 17459 19917 17504
rect 19971 17536 20023 17569
rect 19971 17502 19979 17536
rect 20013 17502 20023 17536
rect 19971 17459 20023 17502
rect 20141 17536 20193 17569
rect 20141 17502 20151 17536
rect 20185 17502 20193 17536
rect 20141 17459 20193 17502
rect 4975 16642 5027 16685
rect 4975 16608 4983 16642
rect 5017 16608 5027 16642
rect 4975 16575 5027 16608
rect 5145 16642 5197 16685
rect 5145 16608 5155 16642
rect 5189 16608 5197 16642
rect 5145 16575 5197 16608
rect 5435 16640 5487 16685
rect 5435 16606 5443 16640
rect 5477 16606 5487 16640
rect 5435 16575 5487 16606
rect 6065 16640 6117 16685
rect 6065 16606 6075 16640
rect 6109 16606 6117 16640
rect 6065 16575 6117 16606
rect 6171 16640 6223 16685
rect 6171 16606 6179 16640
rect 6213 16606 6223 16640
rect 6171 16575 6223 16606
rect 7169 16640 7221 16685
rect 7169 16606 7179 16640
rect 7213 16606 7221 16640
rect 7169 16575 7221 16606
rect 7459 16640 7511 16685
rect 7459 16606 7467 16640
rect 7501 16606 7511 16640
rect 7459 16575 7511 16606
rect 7905 16640 7957 16685
rect 7905 16606 7915 16640
rect 7949 16606 7957 16640
rect 7905 16575 7957 16606
rect 8011 16640 8063 16685
rect 8011 16606 8019 16640
rect 8053 16606 8063 16640
rect 8011 16575 8063 16606
rect 9009 16640 9061 16685
rect 9009 16606 9019 16640
rect 9053 16606 9061 16640
rect 9009 16575 9061 16606
rect 9115 16640 9167 16685
rect 9115 16606 9123 16640
rect 9157 16606 9167 16640
rect 9115 16575 9167 16606
rect 10113 16640 10165 16685
rect 10113 16606 10123 16640
rect 10157 16606 10165 16640
rect 10113 16575 10165 16606
rect 10219 16640 10271 16685
rect 10219 16606 10227 16640
rect 10261 16606 10271 16640
rect 10219 16575 10271 16606
rect 11217 16640 11269 16685
rect 11217 16606 11227 16640
rect 11261 16606 11269 16640
rect 11217 16575 11269 16606
rect 11323 16640 11375 16685
rect 11323 16606 11331 16640
rect 11365 16606 11375 16640
rect 11323 16575 11375 16606
rect 12321 16640 12373 16685
rect 12321 16606 12331 16640
rect 12365 16606 12373 16640
rect 12321 16575 12373 16606
rect 12611 16640 12663 16685
rect 12611 16606 12619 16640
rect 12653 16606 12663 16640
rect 12611 16575 12663 16606
rect 13057 16640 13109 16685
rect 13057 16606 13067 16640
rect 13101 16606 13109 16640
rect 13057 16575 13109 16606
rect 13163 16640 13215 16685
rect 13163 16606 13171 16640
rect 13205 16606 13215 16640
rect 13163 16575 13215 16606
rect 14161 16640 14213 16685
rect 14161 16606 14171 16640
rect 14205 16606 14213 16640
rect 14161 16575 14213 16606
rect 14267 16640 14319 16685
rect 14267 16606 14275 16640
rect 14309 16606 14319 16640
rect 14267 16575 14319 16606
rect 15265 16640 15317 16685
rect 15265 16606 15275 16640
rect 15309 16606 15317 16640
rect 15265 16575 15317 16606
rect 15371 16640 15423 16685
rect 15371 16606 15379 16640
rect 15413 16606 15423 16640
rect 15371 16575 15423 16606
rect 16369 16640 16421 16685
rect 16369 16606 16379 16640
rect 16413 16606 16421 16640
rect 16369 16575 16421 16606
rect 16475 16640 16527 16685
rect 16475 16606 16483 16640
rect 16517 16606 16527 16640
rect 16475 16575 16527 16606
rect 17473 16640 17525 16685
rect 17473 16606 17483 16640
rect 17517 16606 17525 16640
rect 17473 16575 17525 16606
rect 17763 16640 17815 16685
rect 17763 16606 17771 16640
rect 17805 16606 17815 16640
rect 17763 16575 17815 16606
rect 18761 16640 18813 16685
rect 18761 16606 18771 16640
rect 18805 16606 18813 16640
rect 18761 16575 18813 16606
rect 18867 16640 18919 16685
rect 18867 16606 18875 16640
rect 18909 16606 18919 16640
rect 18867 16575 18919 16606
rect 19865 16640 19917 16685
rect 19865 16606 19875 16640
rect 19909 16606 19917 16640
rect 19865 16575 19917 16606
rect 19971 16642 20023 16685
rect 19971 16608 19979 16642
rect 20013 16608 20023 16642
rect 19971 16575 20023 16608
rect 20141 16642 20193 16685
rect 20141 16608 20151 16642
rect 20185 16608 20193 16642
rect 20141 16575 20193 16608
rect 4975 16448 5027 16481
rect 4975 16414 4983 16448
rect 5017 16414 5027 16448
rect 4975 16371 5027 16414
rect 5145 16448 5197 16481
rect 5145 16414 5155 16448
rect 5189 16414 5197 16448
rect 5145 16371 5197 16414
rect 5435 16450 5487 16481
rect 5435 16416 5443 16450
rect 5477 16416 5487 16450
rect 5435 16371 5487 16416
rect 6433 16450 6485 16481
rect 6433 16416 6443 16450
rect 6477 16416 6485 16450
rect 6433 16371 6485 16416
rect 6539 16450 6591 16481
rect 6539 16416 6547 16450
rect 6581 16416 6591 16450
rect 6539 16371 6591 16416
rect 7537 16450 7589 16481
rect 7537 16416 7547 16450
rect 7581 16416 7589 16450
rect 7537 16371 7589 16416
rect 7643 16450 7695 16481
rect 7643 16416 7651 16450
rect 7685 16416 7695 16450
rect 7643 16371 7695 16416
rect 8641 16450 8693 16481
rect 8641 16416 8651 16450
rect 8685 16416 8693 16450
rect 8641 16371 8693 16416
rect 8747 16450 8799 16481
rect 8747 16416 8755 16450
rect 8789 16416 8799 16450
rect 8747 16371 8799 16416
rect 9745 16450 9797 16481
rect 9745 16416 9755 16450
rect 9789 16416 9797 16450
rect 9745 16371 9797 16416
rect 10035 16450 10087 16481
rect 10035 16416 10043 16450
rect 10077 16416 10087 16450
rect 10035 16371 10087 16416
rect 10481 16450 10533 16481
rect 10481 16416 10491 16450
rect 10525 16416 10533 16450
rect 10481 16371 10533 16416
rect 10587 16450 10639 16481
rect 10587 16416 10595 16450
rect 10629 16416 10639 16450
rect 10587 16371 10639 16416
rect 11585 16450 11637 16481
rect 11585 16416 11595 16450
rect 11629 16416 11637 16450
rect 11585 16371 11637 16416
rect 11691 16450 11743 16481
rect 11691 16416 11699 16450
rect 11733 16416 11743 16450
rect 11691 16371 11743 16416
rect 12689 16450 12741 16481
rect 12689 16416 12699 16450
rect 12733 16416 12741 16450
rect 12689 16371 12741 16416
rect 12795 16450 12847 16481
rect 12795 16416 12803 16450
rect 12837 16416 12847 16450
rect 12795 16371 12847 16416
rect 13793 16450 13845 16481
rect 13793 16416 13803 16450
rect 13837 16416 13845 16450
rect 13793 16371 13845 16416
rect 13899 16450 13951 16481
rect 13899 16416 13907 16450
rect 13941 16416 13951 16450
rect 13899 16371 13951 16416
rect 14897 16450 14949 16481
rect 14897 16416 14907 16450
rect 14941 16416 14949 16450
rect 14897 16371 14949 16416
rect 15187 16443 15239 16481
rect 15187 16409 15195 16443
rect 15229 16409 15239 16443
rect 15187 16371 15239 16409
rect 15449 16443 15501 16481
rect 15449 16409 15459 16443
rect 15493 16409 15501 16443
rect 15449 16371 15501 16409
rect 15555 16450 15607 16481
rect 15555 16416 15563 16450
rect 15597 16416 15607 16450
rect 15555 16371 15607 16416
rect 16553 16450 16605 16481
rect 16553 16416 16563 16450
rect 16597 16416 16605 16450
rect 16553 16371 16605 16416
rect 16659 16450 16711 16481
rect 16659 16416 16667 16450
rect 16701 16416 16711 16450
rect 16659 16371 16711 16416
rect 17657 16450 17709 16481
rect 17657 16416 17667 16450
rect 17701 16416 17709 16450
rect 17657 16371 17709 16416
rect 17763 16450 17815 16481
rect 17763 16416 17771 16450
rect 17805 16416 17815 16450
rect 17763 16371 17815 16416
rect 18761 16450 18813 16481
rect 18761 16416 18771 16450
rect 18805 16416 18813 16450
rect 18761 16371 18813 16416
rect 18867 16450 18919 16481
rect 18867 16416 18875 16450
rect 18909 16416 18919 16450
rect 18867 16371 18919 16416
rect 19865 16450 19917 16481
rect 19865 16416 19875 16450
rect 19909 16416 19917 16450
rect 19865 16371 19917 16416
rect 19971 16448 20023 16481
rect 19971 16414 19979 16448
rect 20013 16414 20023 16448
rect 19971 16371 20023 16414
rect 20141 16448 20193 16481
rect 20141 16414 20151 16448
rect 20185 16414 20193 16448
rect 20141 16371 20193 16414
rect 4975 15554 5027 15597
rect 4975 15520 4983 15554
rect 5017 15520 5027 15554
rect 4975 15487 5027 15520
rect 5145 15554 5197 15597
rect 5145 15520 5155 15554
rect 5189 15520 5197 15554
rect 5145 15487 5197 15520
rect 5435 15552 5487 15597
rect 5435 15518 5443 15552
rect 5477 15518 5487 15552
rect 5435 15487 5487 15518
rect 6065 15552 6117 15597
rect 6065 15518 6075 15552
rect 6109 15518 6117 15552
rect 6065 15487 6117 15518
rect 6171 15552 6223 15597
rect 6171 15518 6179 15552
rect 6213 15518 6223 15552
rect 6171 15487 6223 15518
rect 7169 15552 7221 15597
rect 7169 15518 7179 15552
rect 7213 15518 7221 15552
rect 7169 15487 7221 15518
rect 7459 15552 7511 15597
rect 7459 15518 7467 15552
rect 7501 15518 7511 15552
rect 7459 15487 7511 15518
rect 7905 15552 7957 15597
rect 7905 15518 7915 15552
rect 7949 15518 7957 15552
rect 7905 15487 7957 15518
rect 8011 15552 8063 15597
rect 8011 15518 8019 15552
rect 8053 15518 8063 15552
rect 8011 15487 8063 15518
rect 9009 15552 9061 15597
rect 9009 15518 9019 15552
rect 9053 15518 9061 15552
rect 9009 15487 9061 15518
rect 9115 15552 9167 15597
rect 9115 15518 9123 15552
rect 9157 15518 9167 15552
rect 9115 15487 9167 15518
rect 10113 15552 10165 15597
rect 10113 15518 10123 15552
rect 10157 15518 10165 15552
rect 10113 15487 10165 15518
rect 10219 15552 10271 15597
rect 10219 15518 10227 15552
rect 10261 15518 10271 15552
rect 10219 15487 10271 15518
rect 11217 15552 11269 15597
rect 11217 15518 11227 15552
rect 11261 15518 11269 15552
rect 11217 15487 11269 15518
rect 11323 15552 11375 15597
rect 11323 15518 11331 15552
rect 11365 15518 11375 15552
rect 11323 15487 11375 15518
rect 12321 15552 12373 15597
rect 12321 15518 12331 15552
rect 12365 15518 12373 15552
rect 12321 15487 12373 15518
rect 12611 15552 12663 15597
rect 12611 15518 12619 15552
rect 12653 15518 12663 15552
rect 12611 15487 12663 15518
rect 13057 15552 13109 15597
rect 13057 15518 13067 15552
rect 13101 15518 13109 15552
rect 13057 15487 13109 15518
rect 13163 15552 13215 15597
rect 13163 15518 13171 15552
rect 13205 15518 13215 15552
rect 13163 15487 13215 15518
rect 14161 15552 14213 15597
rect 14161 15518 14171 15552
rect 14205 15518 14213 15552
rect 14161 15487 14213 15518
rect 14267 15552 14319 15597
rect 14267 15518 14275 15552
rect 14309 15518 14319 15552
rect 14267 15487 14319 15518
rect 15265 15552 15317 15597
rect 15265 15518 15275 15552
rect 15309 15518 15317 15552
rect 15265 15487 15317 15518
rect 15371 15552 15423 15597
rect 15371 15518 15379 15552
rect 15413 15518 15423 15552
rect 15371 15487 15423 15518
rect 16369 15552 16421 15597
rect 16369 15518 16379 15552
rect 16413 15518 16421 15552
rect 16369 15487 16421 15518
rect 16475 15552 16527 15597
rect 16475 15518 16483 15552
rect 16517 15518 16527 15552
rect 16475 15487 16527 15518
rect 17473 15552 17525 15597
rect 17473 15518 17483 15552
rect 17517 15518 17525 15552
rect 17473 15487 17525 15518
rect 17763 15552 17815 15597
rect 17763 15518 17771 15552
rect 17805 15518 17815 15552
rect 17763 15487 17815 15518
rect 18761 15552 18813 15597
rect 18761 15518 18771 15552
rect 18805 15518 18813 15552
rect 18761 15487 18813 15518
rect 18867 15552 18919 15597
rect 18867 15518 18875 15552
rect 18909 15518 18919 15552
rect 18867 15487 18919 15518
rect 19865 15552 19917 15597
rect 19865 15518 19875 15552
rect 19909 15518 19917 15552
rect 19865 15487 19917 15518
rect 19971 15554 20023 15597
rect 19971 15520 19979 15554
rect 20013 15520 20023 15554
rect 19971 15487 20023 15520
rect 20141 15554 20193 15597
rect 20141 15520 20151 15554
rect 20185 15520 20193 15554
rect 20141 15487 20193 15520
rect 4975 15360 5027 15393
rect 4975 15326 4983 15360
rect 5017 15326 5027 15360
rect 4975 15283 5027 15326
rect 5145 15360 5197 15393
rect 5145 15326 5155 15360
rect 5189 15326 5197 15360
rect 5145 15283 5197 15326
rect 5435 15362 5487 15393
rect 5435 15328 5443 15362
rect 5477 15328 5487 15362
rect 5435 15283 5487 15328
rect 6433 15362 6485 15393
rect 6433 15328 6443 15362
rect 6477 15328 6485 15362
rect 6433 15283 6485 15328
rect 6539 15362 6591 15393
rect 6539 15328 6547 15362
rect 6581 15328 6591 15362
rect 6539 15283 6591 15328
rect 7537 15362 7589 15393
rect 7537 15328 7547 15362
rect 7581 15328 7589 15362
rect 7537 15283 7589 15328
rect 7643 15362 7695 15393
rect 7643 15328 7651 15362
rect 7685 15328 7695 15362
rect 7643 15283 7695 15328
rect 8641 15362 8693 15393
rect 8641 15328 8651 15362
rect 8685 15328 8693 15362
rect 8641 15283 8693 15328
rect 8747 15362 8799 15393
rect 8747 15328 8755 15362
rect 8789 15328 8799 15362
rect 8747 15283 8799 15328
rect 9745 15362 9797 15393
rect 9745 15328 9755 15362
rect 9789 15328 9797 15362
rect 9745 15283 9797 15328
rect 10035 15362 10087 15393
rect 10035 15328 10043 15362
rect 10077 15328 10087 15362
rect 10035 15283 10087 15328
rect 10481 15362 10533 15393
rect 10481 15328 10491 15362
rect 10525 15328 10533 15362
rect 10481 15283 10533 15328
rect 10587 15362 10639 15393
rect 10587 15328 10595 15362
rect 10629 15328 10639 15362
rect 10587 15283 10639 15328
rect 11585 15362 11637 15393
rect 11585 15328 11595 15362
rect 11629 15328 11637 15362
rect 11585 15283 11637 15328
rect 11691 15362 11743 15393
rect 11691 15328 11699 15362
rect 11733 15328 11743 15362
rect 11691 15283 11743 15328
rect 12689 15362 12741 15393
rect 12689 15328 12699 15362
rect 12733 15328 12741 15362
rect 12689 15283 12741 15328
rect 12817 15355 12869 15393
rect 12817 15321 12825 15355
rect 12859 15321 12869 15355
rect 12817 15309 12869 15321
rect 12899 15381 12953 15393
rect 12899 15347 12909 15381
rect 12943 15347 12953 15381
rect 12899 15309 12953 15347
rect 13053 15355 13105 15393
rect 13053 15321 13063 15355
rect 13097 15321 13105 15355
rect 13053 15309 13105 15321
rect 13159 15355 13211 15393
rect 13159 15321 13167 15355
rect 13201 15321 13211 15355
rect 13159 15309 13211 15321
rect 13311 15381 13376 15393
rect 13311 15347 13326 15381
rect 13360 15347 13376 15381
rect 13311 15309 13376 15347
rect 13326 15263 13376 15309
rect 13406 15355 13458 15393
rect 13406 15321 13416 15355
rect 13450 15321 13458 15355
rect 13406 15263 13458 15321
rect 13531 15355 13583 15393
rect 13531 15321 13539 15355
rect 13573 15321 13583 15355
rect 13531 15283 13583 15321
rect 13793 15355 13845 15393
rect 13793 15321 13803 15355
rect 13837 15321 13845 15355
rect 13793 15283 13845 15321
rect 13899 15362 13951 15393
rect 13899 15328 13907 15362
rect 13941 15328 13951 15362
rect 13899 15283 13951 15328
rect 14897 15362 14949 15393
rect 14897 15328 14907 15362
rect 14941 15328 14949 15362
rect 14897 15283 14949 15328
rect 15095 15360 15147 15393
rect 15095 15326 15103 15360
rect 15137 15326 15147 15360
rect 15095 15283 15147 15326
rect 15265 15360 15317 15393
rect 15265 15326 15275 15360
rect 15309 15326 15317 15360
rect 15265 15283 15317 15326
rect 15393 15355 15445 15393
rect 15393 15321 15401 15355
rect 15435 15321 15445 15355
rect 15393 15309 15445 15321
rect 15475 15381 15529 15393
rect 15475 15347 15485 15381
rect 15519 15347 15529 15381
rect 15475 15309 15529 15347
rect 15629 15355 15681 15393
rect 15629 15321 15639 15355
rect 15673 15321 15681 15355
rect 15629 15309 15681 15321
rect 15735 15355 15787 15393
rect 15735 15321 15743 15355
rect 15777 15321 15787 15355
rect 15735 15309 15787 15321
rect 15887 15381 15952 15393
rect 15887 15347 15902 15381
rect 15936 15347 15952 15381
rect 15887 15309 15952 15347
rect 15902 15263 15952 15309
rect 15982 15355 16034 15393
rect 15982 15321 15992 15355
rect 16026 15321 16034 15355
rect 15982 15263 16034 15321
rect 16107 15362 16159 15393
rect 16107 15328 16115 15362
rect 16149 15328 16159 15362
rect 16107 15283 16159 15328
rect 16553 15362 16605 15393
rect 16553 15328 16563 15362
rect 16597 15328 16605 15362
rect 16553 15283 16605 15328
rect 16659 15362 16711 15393
rect 16659 15328 16667 15362
rect 16701 15328 16711 15362
rect 16659 15283 16711 15328
rect 17657 15362 17709 15393
rect 17657 15328 17667 15362
rect 17701 15328 17709 15362
rect 17657 15283 17709 15328
rect 17763 15362 17815 15393
rect 17763 15328 17771 15362
rect 17805 15328 17815 15362
rect 17763 15283 17815 15328
rect 18761 15362 18813 15393
rect 18761 15328 18771 15362
rect 18805 15328 18813 15362
rect 18761 15283 18813 15328
rect 18867 15362 18919 15393
rect 18867 15328 18875 15362
rect 18909 15328 18919 15362
rect 18867 15283 18919 15328
rect 19865 15362 19917 15393
rect 19865 15328 19875 15362
rect 19909 15328 19917 15362
rect 19865 15283 19917 15328
rect 19971 15360 20023 15393
rect 19971 15326 19979 15360
rect 20013 15326 20023 15360
rect 19971 15283 20023 15326
rect 20141 15360 20193 15393
rect 20141 15326 20151 15360
rect 20185 15326 20193 15360
rect 20141 15283 20193 15326
rect 4975 14466 5027 14509
rect 4975 14432 4983 14466
rect 5017 14432 5027 14466
rect 4975 14399 5027 14432
rect 5145 14466 5197 14509
rect 5145 14432 5155 14466
rect 5189 14432 5197 14466
rect 5145 14399 5197 14432
rect 5435 14464 5487 14509
rect 5435 14430 5443 14464
rect 5477 14430 5487 14464
rect 5435 14399 5487 14430
rect 6065 14464 6117 14509
rect 6065 14430 6075 14464
rect 6109 14430 6117 14464
rect 6065 14399 6117 14430
rect 6171 14464 6223 14509
rect 6171 14430 6179 14464
rect 6213 14430 6223 14464
rect 6171 14399 6223 14430
rect 7169 14464 7221 14509
rect 7169 14430 7179 14464
rect 7213 14430 7221 14464
rect 7169 14399 7221 14430
rect 7367 14464 7419 14509
rect 7367 14430 7375 14464
rect 7409 14430 7419 14464
rect 7367 14399 7419 14430
rect 8365 14464 8417 14509
rect 8365 14430 8375 14464
rect 8409 14430 8417 14464
rect 8365 14399 8417 14430
rect 8471 14464 8523 14509
rect 8471 14430 8479 14464
rect 8513 14430 8523 14464
rect 8471 14399 8523 14430
rect 9469 14464 9521 14509
rect 9469 14430 9479 14464
rect 9513 14430 9521 14464
rect 9469 14399 9521 14430
rect 9575 14464 9627 14509
rect 9575 14430 9583 14464
rect 9617 14430 9627 14464
rect 9575 14399 9627 14430
rect 10573 14464 10625 14509
rect 11319 14483 11371 14529
rect 10573 14430 10583 14464
rect 10617 14430 10625 14464
rect 10573 14399 10625 14430
rect 10725 14460 10777 14483
rect 10725 14426 10733 14460
rect 10767 14426 10777 14460
rect 10725 14399 10777 14426
rect 10807 14460 10945 14483
rect 10807 14426 10817 14460
rect 10851 14426 10885 14460
rect 10919 14426 10945 14460
rect 10807 14399 10945 14426
rect 10975 14399 11041 14483
rect 11071 14460 11166 14483
rect 11071 14426 11120 14460
rect 11154 14426 11166 14460
rect 11071 14399 11166 14426
rect 11196 14399 11262 14483
rect 11292 14445 11371 14483
rect 11292 14411 11327 14445
rect 11361 14411 11371 14445
rect 11292 14399 11371 14411
rect 11401 14464 11453 14529
rect 11401 14430 11411 14464
rect 11445 14430 11453 14464
rect 11401 14399 11453 14430
rect 11691 14464 11743 14509
rect 11691 14430 11699 14464
rect 11733 14430 11743 14464
rect 11691 14399 11743 14430
rect 12321 14464 12373 14509
rect 12321 14430 12331 14464
rect 12365 14430 12373 14464
rect 12321 14399 12373 14430
rect 13343 14483 13395 14529
rect 12749 14460 12801 14483
rect 12749 14426 12757 14460
rect 12791 14426 12801 14460
rect 12749 14399 12801 14426
rect 12831 14460 12969 14483
rect 12831 14426 12841 14460
rect 12875 14426 12909 14460
rect 12943 14426 12969 14460
rect 12831 14399 12969 14426
rect 12999 14399 13065 14483
rect 13095 14460 13190 14483
rect 13095 14426 13144 14460
rect 13178 14426 13190 14460
rect 13095 14399 13190 14426
rect 13220 14399 13286 14483
rect 13316 14445 13395 14483
rect 13316 14411 13351 14445
rect 13385 14411 13395 14445
rect 13316 14399 13395 14411
rect 13425 14464 13477 14529
rect 13425 14430 13435 14464
rect 13469 14430 13477 14464
rect 13425 14399 13477 14430
rect 13531 14464 13583 14509
rect 13531 14430 13539 14464
rect 13573 14430 13583 14464
rect 13531 14399 13583 14430
rect 14161 14464 14213 14509
rect 14161 14430 14171 14464
rect 14205 14430 14213 14464
rect 14161 14399 14213 14430
rect 14267 14458 14319 14503
rect 14267 14424 14275 14458
rect 14309 14424 14319 14458
rect 14267 14399 14319 14424
rect 14349 14445 14407 14503
rect 14349 14411 14361 14445
rect 14395 14411 14407 14445
rect 14349 14399 14407 14411
rect 14437 14475 14489 14503
rect 14437 14441 14447 14475
rect 14481 14441 14489 14475
rect 14437 14399 14489 14441
rect 14543 14495 14595 14529
rect 14543 14461 14551 14495
rect 14585 14461 14595 14495
rect 14543 14399 14595 14461
rect 14625 14483 14675 14529
rect 14625 14445 14697 14483
rect 14625 14411 14635 14445
rect 14669 14411 14697 14445
rect 14625 14399 14697 14411
rect 14751 14461 14803 14483
rect 14751 14427 14759 14461
rect 14793 14427 14803 14461
rect 14751 14399 14803 14427
rect 14833 14399 14894 14483
rect 14924 14441 15043 14483
rect 14924 14407 14977 14441
rect 15011 14407 15043 14441
rect 14924 14399 15043 14407
rect 15073 14471 15123 14483
rect 15293 14471 15347 14527
rect 15073 14399 15139 14471
rect 15169 14445 15248 14471
rect 15169 14411 15189 14445
rect 15223 14411 15248 14445
rect 15169 14399 15248 14411
rect 15278 14441 15347 14471
rect 15278 14407 15299 14441
rect 15333 14407 15347 14441
rect 15278 14399 15347 14407
rect 15377 14483 15427 14527
rect 15377 14445 15479 14483
rect 15377 14411 15411 14445
rect 15445 14411 15479 14445
rect 15377 14399 15479 14411
rect 15509 14399 15551 14483
rect 15581 14471 15699 14483
rect 15858 14471 15908 14483
rect 15581 14399 15717 14471
rect 15747 14447 15813 14471
rect 15747 14413 15757 14447
rect 15791 14413 15813 14447
rect 15747 14399 15813 14413
rect 15843 14447 15908 14471
rect 15843 14413 15864 14447
rect 15898 14413 15908 14447
rect 15843 14399 15908 14413
rect 15938 14441 16043 14483
rect 15938 14407 15997 14441
rect 16031 14407 16043 14441
rect 15938 14399 16043 14407
rect 16111 14471 16163 14483
rect 16111 14437 16119 14471
rect 16153 14437 16163 14471
rect 16111 14399 16163 14437
rect 16193 14445 16247 14483
rect 16193 14411 16203 14445
rect 16237 14411 16247 14445
rect 16193 14399 16247 14411
rect 16277 14471 16329 14483
rect 16277 14437 16287 14471
rect 16321 14437 16329 14471
rect 16277 14399 16329 14437
rect 16475 14464 16527 14509
rect 16475 14430 16483 14464
rect 16517 14430 16527 14464
rect 16475 14399 16527 14430
rect 17473 14464 17525 14509
rect 17473 14430 17483 14464
rect 17517 14430 17525 14464
rect 17473 14399 17525 14430
rect 17763 14464 17815 14509
rect 17763 14430 17771 14464
rect 17805 14430 17815 14464
rect 17763 14399 17815 14430
rect 18761 14464 18813 14509
rect 18761 14430 18771 14464
rect 18805 14430 18813 14464
rect 18761 14399 18813 14430
rect 18867 14464 18919 14509
rect 18867 14430 18875 14464
rect 18909 14430 18919 14464
rect 18867 14399 18919 14430
rect 19865 14464 19917 14509
rect 19865 14430 19875 14464
rect 19909 14430 19917 14464
rect 19865 14399 19917 14430
rect 19971 14466 20023 14509
rect 19971 14432 19979 14466
rect 20013 14432 20023 14466
rect 19971 14399 20023 14432
rect 20141 14466 20193 14509
rect 20141 14432 20151 14466
rect 20185 14432 20193 14466
rect 20141 14399 20193 14432
rect 4975 14272 5027 14305
rect 4975 14238 4983 14272
rect 5017 14238 5027 14272
rect 4975 14195 5027 14238
rect 5145 14272 5197 14305
rect 5145 14238 5155 14272
rect 5189 14238 5197 14272
rect 5145 14195 5197 14238
rect 5435 14274 5487 14305
rect 5435 14240 5443 14274
rect 5477 14240 5487 14274
rect 5435 14195 5487 14240
rect 6433 14274 6485 14305
rect 6433 14240 6443 14274
rect 6477 14240 6485 14274
rect 6433 14195 6485 14240
rect 6539 14274 6591 14305
rect 6539 14240 6547 14274
rect 6581 14240 6591 14274
rect 6539 14195 6591 14240
rect 7537 14274 7589 14305
rect 7537 14240 7547 14274
rect 7581 14240 7589 14274
rect 7537 14195 7589 14240
rect 7643 14274 7695 14305
rect 7643 14240 7651 14274
rect 7685 14240 7695 14274
rect 7643 14195 7695 14240
rect 8641 14274 8693 14305
rect 8641 14240 8651 14274
rect 8685 14240 8693 14274
rect 8641 14195 8693 14240
rect 8747 14274 8799 14305
rect 8747 14240 8755 14274
rect 8789 14240 8799 14274
rect 8747 14195 8799 14240
rect 9745 14274 9797 14305
rect 9745 14240 9755 14274
rect 9789 14240 9797 14274
rect 9745 14195 9797 14240
rect 10127 14243 10179 14305
rect 10127 14209 10135 14243
rect 10169 14209 10179 14243
rect 10127 14175 10179 14209
rect 10209 14293 10281 14305
rect 10209 14259 10219 14293
rect 10253 14259 10281 14293
rect 10209 14221 10281 14259
rect 10335 14277 10387 14305
rect 10335 14243 10343 14277
rect 10377 14243 10387 14277
rect 10335 14221 10387 14243
rect 10417 14221 10478 14305
rect 10508 14297 10627 14305
rect 10508 14263 10561 14297
rect 10595 14263 10627 14297
rect 10508 14221 10627 14263
rect 10657 14233 10723 14305
rect 10753 14293 10832 14305
rect 10753 14259 10773 14293
rect 10807 14259 10832 14293
rect 10753 14233 10832 14259
rect 10862 14297 10931 14305
rect 10862 14263 10883 14297
rect 10917 14263 10931 14297
rect 10862 14233 10931 14263
rect 10657 14221 10707 14233
rect 10209 14175 10259 14221
rect 10877 14177 10931 14233
rect 10961 14293 11063 14305
rect 10961 14259 10995 14293
rect 11029 14259 11063 14293
rect 10961 14221 11063 14259
rect 11093 14221 11135 14305
rect 11165 14233 11301 14305
rect 11331 14291 11397 14305
rect 11331 14257 11341 14291
rect 11375 14257 11397 14291
rect 11331 14233 11397 14257
rect 11427 14291 11492 14305
rect 11427 14257 11448 14291
rect 11482 14257 11492 14291
rect 11427 14233 11492 14257
rect 11165 14221 11283 14233
rect 10961 14177 11011 14221
rect 11442 14221 11492 14233
rect 11522 14297 11627 14305
rect 11522 14263 11581 14297
rect 11615 14263 11627 14297
rect 11522 14221 11627 14263
rect 11695 14267 11747 14305
rect 11695 14233 11703 14267
rect 11737 14233 11747 14267
rect 11695 14221 11747 14233
rect 11777 14293 11831 14305
rect 11777 14259 11787 14293
rect 11821 14259 11831 14293
rect 11777 14221 11831 14259
rect 11861 14267 11913 14305
rect 11861 14233 11871 14267
rect 11905 14233 11913 14267
rect 11861 14221 11913 14233
rect 11967 14263 12019 14305
rect 11967 14229 11975 14263
rect 12009 14229 12019 14263
rect 11967 14201 12019 14229
rect 12049 14293 12107 14305
rect 12049 14259 12061 14293
rect 12095 14259 12107 14293
rect 12049 14201 12107 14259
rect 12137 14280 12189 14305
rect 12137 14246 12147 14280
rect 12181 14246 12189 14280
rect 12137 14201 12189 14246
rect 12260 14289 12313 14305
rect 12260 14255 12268 14289
rect 12302 14255 12313 14289
rect 12260 14221 12313 14255
rect 12343 14280 12399 14305
rect 12343 14246 12354 14280
rect 12388 14246 12399 14280
rect 12343 14221 12399 14246
rect 12429 14289 12485 14305
rect 12429 14255 12440 14289
rect 12474 14255 12485 14289
rect 12429 14221 12485 14255
rect 12515 14280 12571 14305
rect 12515 14246 12526 14280
rect 12560 14246 12571 14280
rect 12515 14221 12571 14246
rect 12601 14289 12657 14305
rect 12601 14255 12612 14289
rect 12646 14255 12657 14289
rect 12601 14221 12657 14255
rect 12687 14280 12743 14305
rect 12687 14246 12698 14280
rect 12732 14246 12743 14280
rect 12687 14221 12743 14246
rect 12773 14289 12829 14305
rect 12773 14255 12784 14289
rect 12818 14255 12829 14289
rect 12773 14221 12829 14255
rect 12859 14280 12915 14305
rect 12859 14246 12870 14280
rect 12904 14246 12915 14280
rect 12859 14221 12915 14246
rect 12945 14289 13000 14305
rect 12945 14255 12955 14289
rect 12989 14255 13000 14289
rect 12945 14221 13000 14255
rect 13030 14280 13086 14305
rect 13030 14246 13041 14280
rect 13075 14246 13086 14280
rect 13030 14221 13086 14246
rect 13116 14289 13172 14305
rect 13116 14255 13127 14289
rect 13161 14255 13172 14289
rect 13116 14221 13172 14255
rect 13202 14280 13258 14305
rect 13202 14246 13213 14280
rect 13247 14246 13258 14280
rect 13202 14221 13258 14246
rect 13288 14289 13344 14305
rect 13288 14255 13299 14289
rect 13333 14255 13344 14289
rect 13288 14221 13344 14255
rect 13374 14280 13430 14305
rect 13374 14246 13385 14280
rect 13419 14246 13430 14280
rect 13374 14221 13430 14246
rect 13460 14289 13516 14305
rect 13460 14255 13471 14289
rect 13505 14255 13516 14289
rect 13460 14221 13516 14255
rect 13546 14280 13602 14305
rect 13546 14246 13557 14280
rect 13591 14246 13602 14280
rect 13546 14221 13602 14246
rect 13632 14280 13688 14305
rect 13632 14246 13643 14280
rect 13677 14246 13688 14280
rect 13632 14221 13688 14246
rect 13718 14280 13774 14305
rect 13718 14246 13729 14280
rect 13763 14246 13774 14280
rect 13718 14221 13774 14246
rect 13804 14280 13860 14305
rect 13804 14246 13815 14280
rect 13849 14246 13860 14280
rect 13804 14221 13860 14246
rect 13890 14280 13946 14305
rect 13890 14246 13901 14280
rect 13935 14246 13946 14280
rect 13890 14221 13946 14246
rect 13976 14293 14029 14305
rect 13976 14259 13987 14293
rect 14021 14259 14029 14293
rect 13976 14221 14029 14259
rect 14289 14267 14341 14305
rect 14289 14233 14297 14267
rect 14331 14233 14341 14267
rect 14289 14221 14341 14233
rect 14371 14293 14425 14305
rect 14371 14259 14381 14293
rect 14415 14259 14425 14293
rect 14371 14221 14425 14259
rect 14525 14267 14577 14305
rect 14525 14233 14535 14267
rect 14569 14233 14577 14267
rect 14525 14221 14577 14233
rect 14631 14267 14683 14305
rect 14631 14233 14639 14267
rect 14673 14233 14683 14267
rect 14631 14221 14683 14233
rect 14783 14293 14848 14305
rect 14783 14259 14798 14293
rect 14832 14259 14848 14293
rect 14783 14221 14848 14259
rect 14798 14175 14848 14221
rect 14878 14267 14930 14305
rect 14878 14233 14888 14267
rect 14922 14233 14930 14267
rect 14878 14175 14930 14233
rect 15187 14274 15239 14305
rect 15187 14240 15195 14274
rect 15229 14240 15239 14274
rect 15187 14175 15239 14240
rect 15269 14293 15348 14305
rect 15269 14259 15279 14293
rect 15313 14259 15348 14293
rect 15269 14221 15348 14259
rect 15378 14221 15444 14305
rect 15474 14278 15569 14305
rect 15474 14244 15486 14278
rect 15520 14244 15569 14278
rect 15474 14221 15569 14244
rect 15599 14221 15665 14305
rect 15695 14278 15833 14305
rect 15695 14244 15721 14278
rect 15755 14244 15789 14278
rect 15823 14244 15833 14278
rect 15695 14221 15833 14244
rect 15863 14278 15915 14305
rect 15863 14244 15873 14278
rect 15907 14244 15915 14278
rect 15863 14221 15915 14244
rect 16015 14263 16067 14305
rect 16015 14229 16023 14263
rect 16057 14229 16067 14263
rect 15269 14175 15321 14221
rect 16015 14201 16067 14229
rect 16097 14293 16155 14305
rect 16097 14259 16109 14293
rect 16143 14259 16155 14293
rect 16097 14201 16155 14259
rect 16185 14280 16237 14305
rect 16185 14246 16195 14280
rect 16229 14246 16237 14280
rect 16185 14201 16237 14246
rect 16291 14263 16343 14305
rect 16291 14229 16299 14263
rect 16333 14229 16343 14263
rect 16291 14201 16343 14229
rect 16373 14293 16431 14305
rect 16373 14259 16385 14293
rect 16419 14259 16431 14293
rect 16373 14201 16431 14259
rect 16461 14280 16513 14305
rect 16461 14246 16471 14280
rect 16505 14246 16513 14280
rect 16461 14201 16513 14246
rect 16659 14274 16711 14305
rect 16659 14240 16667 14274
rect 16701 14240 16711 14274
rect 16659 14195 16711 14240
rect 17657 14274 17709 14305
rect 17657 14240 17667 14274
rect 17701 14240 17709 14274
rect 17657 14195 17709 14240
rect 17763 14274 17815 14305
rect 17763 14240 17771 14274
rect 17805 14240 17815 14274
rect 17763 14195 17815 14240
rect 18761 14274 18813 14305
rect 18761 14240 18771 14274
rect 18805 14240 18813 14274
rect 18761 14195 18813 14240
rect 18867 14274 18919 14305
rect 18867 14240 18875 14274
rect 18909 14240 18919 14274
rect 18867 14195 18919 14240
rect 19865 14274 19917 14305
rect 19865 14240 19875 14274
rect 19909 14240 19917 14274
rect 19865 14195 19917 14240
rect 19971 14272 20023 14305
rect 19971 14238 19979 14272
rect 20013 14238 20023 14272
rect 19971 14195 20023 14238
rect 20141 14272 20193 14305
rect 20141 14238 20151 14272
rect 20185 14238 20193 14272
rect 20141 14195 20193 14238
rect 4975 13378 5027 13421
rect 4975 13344 4983 13378
rect 5017 13344 5027 13378
rect 4975 13311 5027 13344
rect 5145 13378 5197 13421
rect 5145 13344 5155 13378
rect 5189 13344 5197 13378
rect 5145 13311 5197 13344
rect 5435 13376 5487 13421
rect 5435 13342 5443 13376
rect 5477 13342 5487 13376
rect 5435 13311 5487 13342
rect 6065 13376 6117 13421
rect 6065 13342 6075 13376
rect 6109 13342 6117 13376
rect 6065 13311 6117 13342
rect 6171 13376 6223 13421
rect 6171 13342 6179 13376
rect 6213 13342 6223 13376
rect 6171 13311 6223 13342
rect 7169 13376 7221 13421
rect 7169 13342 7179 13376
rect 7213 13342 7221 13376
rect 7169 13311 7221 13342
rect 7459 13376 7511 13421
rect 7459 13342 7467 13376
rect 7501 13342 7511 13376
rect 7459 13311 7511 13342
rect 8457 13376 8509 13421
rect 8457 13342 8467 13376
rect 8501 13342 8509 13376
rect 8457 13311 8509 13342
rect 8563 13376 8615 13421
rect 8563 13342 8571 13376
rect 8605 13342 8615 13376
rect 8563 13311 8615 13342
rect 9561 13376 9613 13421
rect 9561 13342 9571 13376
rect 9605 13342 9613 13376
rect 9561 13311 9613 13342
rect 9667 13370 9719 13415
rect 9667 13336 9675 13370
rect 9709 13336 9719 13370
rect 9667 13311 9719 13336
rect 9749 13357 9807 13415
rect 9749 13323 9761 13357
rect 9795 13323 9807 13357
rect 9749 13311 9807 13323
rect 9837 13387 9889 13415
rect 9837 13353 9847 13387
rect 9881 13353 9889 13387
rect 9837 13311 9889 13353
rect 9960 13361 10013 13395
rect 9960 13327 9968 13361
rect 10002 13327 10013 13361
rect 9960 13311 10013 13327
rect 10043 13370 10099 13395
rect 10043 13336 10054 13370
rect 10088 13336 10099 13370
rect 10043 13311 10099 13336
rect 10129 13361 10185 13395
rect 10129 13327 10140 13361
rect 10174 13327 10185 13361
rect 10129 13311 10185 13327
rect 10215 13370 10271 13395
rect 10215 13336 10226 13370
rect 10260 13336 10271 13370
rect 10215 13311 10271 13336
rect 10301 13361 10357 13395
rect 10301 13327 10312 13361
rect 10346 13327 10357 13361
rect 10301 13311 10357 13327
rect 10387 13370 10443 13395
rect 10387 13336 10398 13370
rect 10432 13336 10443 13370
rect 10387 13311 10443 13336
rect 10473 13361 10529 13395
rect 10473 13327 10484 13361
rect 10518 13327 10529 13361
rect 10473 13311 10529 13327
rect 10559 13370 10615 13395
rect 10559 13336 10570 13370
rect 10604 13336 10615 13370
rect 10559 13311 10615 13336
rect 10645 13361 10700 13395
rect 10645 13327 10655 13361
rect 10689 13327 10700 13361
rect 10645 13311 10700 13327
rect 10730 13370 10786 13395
rect 10730 13336 10741 13370
rect 10775 13336 10786 13370
rect 10730 13311 10786 13336
rect 10816 13361 10872 13395
rect 10816 13327 10827 13361
rect 10861 13327 10872 13361
rect 10816 13311 10872 13327
rect 10902 13370 10958 13395
rect 10902 13336 10913 13370
rect 10947 13336 10958 13370
rect 10902 13311 10958 13336
rect 10988 13361 11044 13395
rect 10988 13327 10999 13361
rect 11033 13327 11044 13361
rect 10988 13311 11044 13327
rect 11074 13370 11130 13395
rect 11074 13336 11085 13370
rect 11119 13336 11130 13370
rect 11074 13311 11130 13336
rect 11160 13361 11216 13395
rect 11160 13327 11171 13361
rect 11205 13327 11216 13361
rect 11160 13311 11216 13327
rect 11246 13370 11302 13395
rect 11246 13336 11257 13370
rect 11291 13336 11302 13370
rect 11246 13311 11302 13336
rect 11332 13370 11388 13395
rect 11332 13336 11343 13370
rect 11377 13336 11388 13370
rect 11332 13311 11388 13336
rect 11418 13370 11474 13395
rect 11418 13336 11429 13370
rect 11463 13336 11474 13370
rect 11418 13311 11474 13336
rect 11504 13370 11560 13395
rect 11504 13336 11515 13370
rect 11549 13336 11560 13370
rect 11504 13311 11560 13336
rect 11590 13370 11646 13395
rect 11590 13336 11601 13370
rect 11635 13336 11646 13370
rect 11590 13311 11646 13336
rect 11676 13357 11729 13395
rect 11676 13323 11687 13357
rect 11721 13323 11729 13357
rect 11676 13311 11729 13323
rect 11875 13376 11927 13421
rect 11875 13342 11883 13376
rect 11917 13342 11927 13376
rect 11875 13311 11927 13342
rect 12321 13376 12373 13421
rect 12321 13342 12331 13376
rect 12365 13342 12373 13376
rect 12321 13311 12373 13342
rect 12519 13387 12571 13415
rect 12519 13353 12527 13387
rect 12561 13353 12571 13387
rect 12519 13311 12571 13353
rect 12601 13357 12659 13415
rect 12601 13323 12613 13357
rect 12647 13323 12659 13357
rect 12601 13311 12659 13323
rect 12689 13370 12741 13415
rect 12689 13336 12699 13370
rect 12733 13336 12741 13370
rect 12689 13311 12741 13336
rect 12887 13407 12939 13441
rect 12887 13373 12895 13407
rect 12929 13373 12939 13407
rect 12887 13311 12939 13373
rect 12969 13395 13019 13441
rect 12969 13357 13041 13395
rect 12969 13323 12979 13357
rect 13013 13323 13041 13357
rect 12969 13311 13041 13323
rect 13095 13373 13147 13395
rect 13095 13339 13103 13373
rect 13137 13339 13147 13373
rect 13095 13311 13147 13339
rect 13177 13311 13238 13395
rect 13268 13353 13387 13395
rect 13268 13319 13321 13353
rect 13355 13319 13387 13353
rect 13268 13311 13387 13319
rect 13417 13383 13467 13395
rect 13637 13383 13691 13439
rect 13417 13311 13483 13383
rect 13513 13357 13592 13383
rect 13513 13323 13533 13357
rect 13567 13323 13592 13357
rect 13513 13311 13592 13323
rect 13622 13353 13691 13383
rect 13622 13319 13643 13353
rect 13677 13319 13691 13353
rect 13622 13311 13691 13319
rect 13721 13395 13771 13439
rect 13721 13357 13823 13395
rect 13721 13323 13755 13357
rect 13789 13323 13823 13357
rect 13721 13311 13823 13323
rect 13853 13311 13895 13395
rect 13925 13383 14043 13395
rect 14202 13383 14252 13395
rect 13925 13311 14061 13383
rect 14091 13359 14157 13383
rect 14091 13325 14101 13359
rect 14135 13325 14157 13359
rect 14091 13311 14157 13325
rect 14187 13359 14252 13383
rect 14187 13325 14208 13359
rect 14242 13325 14252 13359
rect 14187 13311 14252 13325
rect 14282 13353 14387 13395
rect 14282 13319 14341 13353
rect 14375 13319 14387 13353
rect 14282 13311 14387 13319
rect 14455 13383 14507 13395
rect 14455 13349 14463 13383
rect 14497 13349 14507 13383
rect 14455 13311 14507 13349
rect 14537 13357 14591 13395
rect 14537 13323 14547 13357
rect 14581 13323 14591 13357
rect 14537 13311 14591 13323
rect 14621 13383 14673 13395
rect 14621 13349 14631 13383
rect 14665 13349 14673 13383
rect 14621 13311 14673 13349
rect 14727 13357 14780 13395
rect 14727 13323 14735 13357
rect 14769 13323 14780 13357
rect 14727 13311 14780 13323
rect 14810 13370 14866 13395
rect 14810 13336 14821 13370
rect 14855 13336 14866 13370
rect 14810 13311 14866 13336
rect 14896 13370 14952 13395
rect 14896 13336 14907 13370
rect 14941 13336 14952 13370
rect 14896 13311 14952 13336
rect 14982 13370 15038 13395
rect 14982 13336 14993 13370
rect 15027 13336 15038 13370
rect 14982 13311 15038 13336
rect 15068 13370 15124 13395
rect 15068 13336 15079 13370
rect 15113 13336 15124 13370
rect 15068 13311 15124 13336
rect 15154 13370 15210 13395
rect 15154 13336 15165 13370
rect 15199 13336 15210 13370
rect 15154 13311 15210 13336
rect 15240 13361 15296 13395
rect 15240 13327 15251 13361
rect 15285 13327 15296 13361
rect 15240 13311 15296 13327
rect 15326 13370 15382 13395
rect 15326 13336 15337 13370
rect 15371 13336 15382 13370
rect 15326 13311 15382 13336
rect 15412 13361 15468 13395
rect 15412 13327 15423 13361
rect 15457 13327 15468 13361
rect 15412 13311 15468 13327
rect 15498 13370 15554 13395
rect 15498 13336 15509 13370
rect 15543 13336 15554 13370
rect 15498 13311 15554 13336
rect 15584 13361 15640 13395
rect 15584 13327 15595 13361
rect 15629 13327 15640 13361
rect 15584 13311 15640 13327
rect 15670 13370 15726 13395
rect 15670 13336 15681 13370
rect 15715 13336 15726 13370
rect 15670 13311 15726 13336
rect 15756 13361 15811 13395
rect 15756 13327 15767 13361
rect 15801 13327 15811 13361
rect 15756 13311 15811 13327
rect 15841 13370 15897 13395
rect 15841 13336 15852 13370
rect 15886 13336 15897 13370
rect 15841 13311 15897 13336
rect 15927 13361 15983 13395
rect 15927 13327 15938 13361
rect 15972 13327 15983 13361
rect 15927 13311 15983 13327
rect 16013 13370 16069 13395
rect 16013 13336 16024 13370
rect 16058 13336 16069 13370
rect 16013 13311 16069 13336
rect 16099 13361 16155 13395
rect 16099 13327 16110 13361
rect 16144 13327 16155 13361
rect 16099 13311 16155 13327
rect 16185 13370 16241 13395
rect 16185 13336 16196 13370
rect 16230 13336 16241 13370
rect 16185 13311 16241 13336
rect 16271 13361 16327 13395
rect 16271 13327 16282 13361
rect 16316 13327 16327 13361
rect 16271 13311 16327 13327
rect 16357 13370 16413 13395
rect 16357 13336 16368 13370
rect 16402 13336 16413 13370
rect 16357 13311 16413 13336
rect 16443 13361 16496 13395
rect 16443 13327 16454 13361
rect 16488 13327 16496 13361
rect 16443 13311 16496 13327
rect 16567 13376 16619 13441
rect 16567 13342 16575 13376
rect 16609 13342 16619 13376
rect 16567 13311 16619 13342
rect 16649 13395 16701 13441
rect 16649 13357 16728 13395
rect 16649 13323 16659 13357
rect 16693 13323 16728 13357
rect 16649 13311 16728 13323
rect 16758 13311 16824 13395
rect 16854 13372 16949 13395
rect 16854 13338 16866 13372
rect 16900 13338 16949 13372
rect 16854 13311 16949 13338
rect 16979 13311 17045 13395
rect 17075 13372 17213 13395
rect 17075 13338 17101 13372
rect 17135 13338 17169 13372
rect 17203 13338 17213 13372
rect 17075 13311 17213 13338
rect 17243 13372 17295 13395
rect 17243 13338 17253 13372
rect 17287 13338 17295 13372
rect 17243 13311 17295 13338
rect 17763 13376 17815 13421
rect 17763 13342 17771 13376
rect 17805 13342 17815 13376
rect 17763 13311 17815 13342
rect 18761 13376 18813 13421
rect 18761 13342 18771 13376
rect 18805 13342 18813 13376
rect 18761 13311 18813 13342
rect 18867 13376 18919 13421
rect 18867 13342 18875 13376
rect 18909 13342 18919 13376
rect 18867 13311 18919 13342
rect 19865 13376 19917 13421
rect 19865 13342 19875 13376
rect 19909 13342 19917 13376
rect 19865 13311 19917 13342
rect 19971 13378 20023 13421
rect 19971 13344 19979 13378
rect 20013 13344 20023 13378
rect 19971 13311 20023 13344
rect 20141 13378 20193 13421
rect 20141 13344 20151 13378
rect 20185 13344 20193 13378
rect 20141 13311 20193 13344
rect 4975 13184 5027 13217
rect 4975 13150 4983 13184
rect 5017 13150 5027 13184
rect 4975 13107 5027 13150
rect 5145 13184 5197 13217
rect 5145 13150 5155 13184
rect 5189 13150 5197 13184
rect 5145 13107 5197 13150
rect 5251 13186 5303 13217
rect 5251 13152 5259 13186
rect 5293 13152 5303 13186
rect 5251 13107 5303 13152
rect 5697 13186 5749 13217
rect 5697 13152 5707 13186
rect 5741 13152 5749 13186
rect 5697 13107 5749 13152
rect 5803 13186 5855 13217
rect 5803 13152 5811 13186
rect 5845 13152 5855 13186
rect 5803 13107 5855 13152
rect 6801 13186 6853 13217
rect 6801 13152 6811 13186
rect 6845 13152 6853 13186
rect 6801 13107 6853 13152
rect 6907 13186 6959 13217
rect 6907 13152 6915 13186
rect 6949 13152 6959 13186
rect 6907 13107 6959 13152
rect 7905 13186 7957 13217
rect 7905 13152 7915 13186
rect 7949 13152 7957 13186
rect 7905 13107 7957 13152
rect 8011 13186 8063 13217
rect 8011 13152 8019 13186
rect 8053 13152 8063 13186
rect 8011 13107 8063 13152
rect 9009 13186 9061 13217
rect 9009 13152 9019 13186
rect 9053 13152 9061 13186
rect 9009 13107 9061 13152
rect 9137 13179 9189 13217
rect 9137 13145 9145 13179
rect 9179 13145 9189 13179
rect 9137 13133 9189 13145
rect 9219 13205 9273 13217
rect 9219 13171 9229 13205
rect 9263 13171 9273 13205
rect 9219 13133 9273 13171
rect 9373 13179 9425 13217
rect 9373 13145 9383 13179
rect 9417 13145 9425 13179
rect 9373 13133 9425 13145
rect 9479 13179 9531 13217
rect 9479 13145 9487 13179
rect 9521 13145 9531 13179
rect 9479 13133 9531 13145
rect 9631 13205 9696 13217
rect 9631 13171 9646 13205
rect 9680 13171 9696 13205
rect 9631 13133 9696 13171
rect 9646 13087 9696 13133
rect 9726 13179 9778 13217
rect 9726 13145 9736 13179
rect 9770 13145 9778 13179
rect 9726 13087 9778 13145
rect 10035 13179 10087 13217
rect 10035 13145 10043 13179
rect 10077 13145 10087 13179
rect 10035 13107 10087 13145
rect 10297 13179 10349 13217
rect 10297 13145 10307 13179
rect 10341 13145 10349 13179
rect 10297 13107 10349 13145
rect 10403 13155 10455 13217
rect 10403 13121 10411 13155
rect 10445 13121 10455 13155
rect 10403 13087 10455 13121
rect 10485 13205 10557 13217
rect 10485 13171 10495 13205
rect 10529 13171 10557 13205
rect 10485 13133 10557 13171
rect 10611 13189 10663 13217
rect 10611 13155 10619 13189
rect 10653 13155 10663 13189
rect 10611 13133 10663 13155
rect 10693 13133 10754 13217
rect 10784 13209 10903 13217
rect 10784 13175 10837 13209
rect 10871 13175 10903 13209
rect 10784 13133 10903 13175
rect 10933 13145 10999 13217
rect 11029 13205 11108 13217
rect 11029 13171 11049 13205
rect 11083 13171 11108 13205
rect 11029 13145 11108 13171
rect 11138 13209 11207 13217
rect 11138 13175 11159 13209
rect 11193 13175 11207 13209
rect 11138 13145 11207 13175
rect 10933 13133 10983 13145
rect 10485 13087 10535 13133
rect 11153 13089 11207 13145
rect 11237 13205 11339 13217
rect 11237 13171 11271 13205
rect 11305 13171 11339 13205
rect 11237 13133 11339 13171
rect 11369 13133 11411 13217
rect 11441 13145 11577 13217
rect 11607 13203 11673 13217
rect 11607 13169 11617 13203
rect 11651 13169 11673 13203
rect 11607 13145 11673 13169
rect 11703 13203 11768 13217
rect 11703 13169 11724 13203
rect 11758 13169 11768 13203
rect 11703 13145 11768 13169
rect 11441 13133 11559 13145
rect 11237 13089 11287 13133
rect 11718 13133 11768 13145
rect 11798 13209 11903 13217
rect 11798 13175 11857 13209
rect 11891 13175 11903 13209
rect 11798 13133 11903 13175
rect 11971 13179 12023 13217
rect 11971 13145 11979 13179
rect 12013 13145 12023 13179
rect 11971 13133 12023 13145
rect 12053 13205 12107 13217
rect 12053 13171 12063 13205
rect 12097 13171 12107 13205
rect 12053 13133 12107 13171
rect 12137 13179 12189 13217
rect 12137 13145 12147 13179
rect 12181 13145 12189 13179
rect 12137 13133 12189 13145
rect 12243 13179 12295 13217
rect 12243 13145 12251 13179
rect 12285 13145 12295 13179
rect 12243 13133 12295 13145
rect 12325 13205 12379 13217
rect 12325 13171 12335 13205
rect 12369 13171 12379 13205
rect 12325 13133 12379 13171
rect 12409 13179 12461 13217
rect 12409 13145 12419 13179
rect 12453 13145 12461 13179
rect 12409 13133 12461 13145
rect 12529 13209 12634 13217
rect 12529 13175 12541 13209
rect 12575 13175 12634 13209
rect 12529 13133 12634 13175
rect 12664 13203 12729 13217
rect 12664 13169 12674 13203
rect 12708 13169 12729 13203
rect 12664 13145 12729 13169
rect 12759 13203 12825 13217
rect 12759 13169 12781 13203
rect 12815 13169 12825 13203
rect 12759 13145 12825 13169
rect 12855 13145 12991 13217
rect 12664 13133 12714 13145
rect 12873 13133 12991 13145
rect 13021 13133 13063 13217
rect 13093 13205 13195 13217
rect 13093 13171 13127 13205
rect 13161 13171 13195 13205
rect 13093 13133 13195 13171
rect 13145 13089 13195 13133
rect 13225 13209 13294 13217
rect 13225 13175 13239 13209
rect 13273 13175 13294 13209
rect 13225 13145 13294 13175
rect 13324 13205 13403 13217
rect 13324 13171 13349 13205
rect 13383 13171 13403 13205
rect 13324 13145 13403 13171
rect 13433 13145 13499 13217
rect 13225 13089 13279 13145
rect 13449 13133 13499 13145
rect 13529 13209 13648 13217
rect 13529 13175 13561 13209
rect 13595 13175 13648 13209
rect 13529 13133 13648 13175
rect 13678 13133 13739 13217
rect 13769 13189 13821 13217
rect 13769 13155 13779 13189
rect 13813 13155 13821 13189
rect 13769 13133 13821 13155
rect 13875 13205 13947 13217
rect 13875 13171 13903 13205
rect 13937 13171 13947 13205
rect 13875 13133 13947 13171
rect 13897 13087 13947 13133
rect 13977 13155 14029 13217
rect 13977 13121 13987 13155
rect 14021 13121 14029 13155
rect 13977 13087 14029 13121
rect 14083 13186 14135 13217
rect 14083 13152 14091 13186
rect 14125 13152 14135 13186
rect 14083 13087 14135 13152
rect 14165 13205 14244 13217
rect 14165 13171 14175 13205
rect 14209 13171 14244 13205
rect 14165 13133 14244 13171
rect 14274 13133 14340 13217
rect 14370 13190 14465 13217
rect 14370 13156 14382 13190
rect 14416 13156 14465 13190
rect 14370 13133 14465 13156
rect 14495 13133 14561 13217
rect 14591 13190 14729 13217
rect 14591 13156 14617 13190
rect 14651 13156 14685 13190
rect 14719 13156 14729 13190
rect 14591 13133 14729 13156
rect 14759 13190 14811 13217
rect 14759 13156 14769 13190
rect 14803 13156 14811 13190
rect 14759 13133 14811 13156
rect 14165 13087 14217 13133
rect 15095 13155 15147 13217
rect 15095 13121 15103 13155
rect 15137 13121 15147 13155
rect 15095 13087 15147 13121
rect 15177 13205 15249 13217
rect 15177 13171 15187 13205
rect 15221 13171 15249 13205
rect 15177 13133 15249 13171
rect 15303 13189 15355 13217
rect 15303 13155 15311 13189
rect 15345 13155 15355 13189
rect 15303 13133 15355 13155
rect 15385 13133 15446 13217
rect 15476 13209 15595 13217
rect 15476 13175 15529 13209
rect 15563 13175 15595 13209
rect 15476 13133 15595 13175
rect 15625 13145 15691 13217
rect 15721 13205 15800 13217
rect 15721 13171 15741 13205
rect 15775 13171 15800 13205
rect 15721 13145 15800 13171
rect 15830 13209 15899 13217
rect 15830 13175 15851 13209
rect 15885 13175 15899 13209
rect 15830 13145 15899 13175
rect 15625 13133 15675 13145
rect 15177 13087 15227 13133
rect 15845 13089 15899 13145
rect 15929 13205 16031 13217
rect 15929 13171 15963 13205
rect 15997 13171 16031 13205
rect 15929 13133 16031 13171
rect 16061 13133 16103 13217
rect 16133 13145 16269 13217
rect 16299 13203 16365 13217
rect 16299 13169 16309 13203
rect 16343 13169 16365 13203
rect 16299 13145 16365 13169
rect 16395 13203 16460 13217
rect 16395 13169 16416 13203
rect 16450 13169 16460 13203
rect 16395 13145 16460 13169
rect 16133 13133 16251 13145
rect 15929 13089 15979 13133
rect 16410 13133 16460 13145
rect 16490 13209 16595 13217
rect 16490 13175 16549 13209
rect 16583 13175 16595 13209
rect 16490 13133 16595 13175
rect 16663 13179 16715 13217
rect 16663 13145 16671 13179
rect 16705 13145 16715 13179
rect 16663 13133 16715 13145
rect 16745 13205 16799 13217
rect 16745 13171 16755 13205
rect 16789 13171 16799 13205
rect 16745 13133 16799 13171
rect 16829 13179 16881 13217
rect 16829 13145 16839 13179
rect 16873 13145 16881 13179
rect 16829 13133 16881 13145
rect 16954 13179 17006 13217
rect 16954 13145 16962 13179
rect 16996 13145 17006 13179
rect 16954 13087 17006 13145
rect 17036 13205 17101 13217
rect 17036 13171 17052 13205
rect 17086 13171 17101 13205
rect 17036 13133 17101 13171
rect 17201 13179 17253 13217
rect 17201 13145 17211 13179
rect 17245 13145 17253 13179
rect 17201 13133 17253 13145
rect 17307 13179 17359 13217
rect 17307 13145 17315 13179
rect 17349 13145 17359 13179
rect 17307 13133 17359 13145
rect 17459 13205 17513 13217
rect 17459 13171 17469 13205
rect 17503 13171 17513 13205
rect 17459 13133 17513 13171
rect 17543 13179 17595 13217
rect 17543 13145 17553 13179
rect 17587 13145 17595 13179
rect 17543 13133 17595 13145
rect 17763 13186 17815 13217
rect 17763 13152 17771 13186
rect 17805 13152 17815 13186
rect 17036 13087 17086 13133
rect 17763 13107 17815 13152
rect 18761 13186 18813 13217
rect 18761 13152 18771 13186
rect 18805 13152 18813 13186
rect 18761 13107 18813 13152
rect 18867 13186 18919 13217
rect 18867 13152 18875 13186
rect 18909 13152 18919 13186
rect 18867 13107 18919 13152
rect 19865 13186 19917 13217
rect 19865 13152 19875 13186
rect 19909 13152 19917 13186
rect 19865 13107 19917 13152
rect 19971 13184 20023 13217
rect 19971 13150 19979 13184
rect 20013 13150 20023 13184
rect 19971 13107 20023 13150
rect 20141 13184 20193 13217
rect 20141 13150 20151 13184
rect 20185 13150 20193 13184
rect 20141 13107 20193 13150
rect 4975 12290 5027 12333
rect 4975 12256 4983 12290
rect 5017 12256 5027 12290
rect 4975 12223 5027 12256
rect 5145 12290 5197 12333
rect 5145 12256 5155 12290
rect 5189 12256 5197 12290
rect 5145 12223 5197 12256
rect 5619 12288 5671 12333
rect 5619 12254 5627 12288
rect 5661 12254 5671 12288
rect 5619 12223 5671 12254
rect 6617 12288 6669 12333
rect 6617 12254 6627 12288
rect 6661 12254 6669 12288
rect 6617 12223 6669 12254
rect 6725 12273 6783 12307
rect 6725 12239 6738 12273
rect 6772 12239 6783 12273
rect 6725 12223 6783 12239
rect 6813 12295 6869 12307
rect 6813 12261 6824 12295
rect 6858 12261 6869 12295
rect 6813 12223 6869 12261
rect 6899 12273 6955 12307
rect 6899 12239 6910 12273
rect 6944 12239 6955 12273
rect 6899 12223 6955 12239
rect 6985 12295 7041 12307
rect 6985 12261 6996 12295
rect 7030 12261 7041 12295
rect 6985 12223 7041 12261
rect 7071 12273 7138 12307
rect 7071 12239 7093 12273
rect 7127 12239 7138 12273
rect 7071 12223 7138 12239
rect 7168 12277 7221 12307
rect 7168 12243 7179 12277
rect 7213 12243 7221 12277
rect 7168 12223 7221 12243
rect 7367 12295 7419 12333
rect 7367 12261 7375 12295
rect 7409 12261 7419 12295
rect 7367 12223 7419 12261
rect 7629 12295 7681 12333
rect 7629 12261 7639 12295
rect 7673 12261 7681 12295
rect 7629 12223 7681 12261
rect 7735 12288 7787 12333
rect 7735 12254 7743 12288
rect 7777 12254 7787 12288
rect 7735 12223 7787 12254
rect 8733 12288 8785 12333
rect 8733 12254 8743 12288
rect 8777 12254 8785 12288
rect 8733 12223 8785 12254
rect 8841 12273 8899 12307
rect 8841 12239 8854 12273
rect 8888 12239 8899 12273
rect 8841 12223 8899 12239
rect 8929 12295 8985 12307
rect 8929 12261 8940 12295
rect 8974 12261 8985 12295
rect 8929 12223 8985 12261
rect 9015 12273 9071 12307
rect 9015 12239 9026 12273
rect 9060 12239 9071 12273
rect 9015 12223 9071 12239
rect 9101 12295 9157 12307
rect 9101 12261 9112 12295
rect 9146 12261 9157 12295
rect 9101 12223 9157 12261
rect 9187 12273 9254 12307
rect 9187 12239 9209 12273
rect 9243 12239 9254 12273
rect 9187 12223 9254 12239
rect 9284 12277 9337 12307
rect 9284 12243 9295 12277
rect 9329 12243 9337 12277
rect 9284 12223 9337 12243
rect 9483 12295 9535 12333
rect 9483 12261 9491 12295
rect 9525 12261 9535 12295
rect 9483 12223 9535 12261
rect 9745 12295 9797 12333
rect 9745 12261 9755 12295
rect 9789 12261 9797 12295
rect 9745 12223 9797 12261
rect 9945 12273 10003 12307
rect 9945 12239 9958 12273
rect 9992 12239 10003 12273
rect 9945 12223 10003 12239
rect 10033 12295 10089 12307
rect 10033 12261 10044 12295
rect 10078 12261 10089 12295
rect 10033 12223 10089 12261
rect 10119 12273 10175 12307
rect 10119 12239 10130 12273
rect 10164 12239 10175 12273
rect 10119 12223 10175 12239
rect 10205 12295 10261 12307
rect 10205 12261 10216 12295
rect 10250 12261 10261 12295
rect 10205 12223 10261 12261
rect 10291 12273 10358 12307
rect 10291 12239 10313 12273
rect 10347 12239 10358 12273
rect 10291 12223 10358 12239
rect 10388 12277 10441 12307
rect 10388 12243 10399 12277
rect 10433 12243 10441 12277
rect 10388 12223 10441 12243
rect 10495 12288 10547 12353
rect 10495 12254 10503 12288
rect 10537 12254 10547 12288
rect 10495 12223 10547 12254
rect 10577 12307 10629 12353
rect 12055 12307 12107 12353
rect 10577 12269 10656 12307
rect 10577 12235 10587 12269
rect 10621 12235 10656 12269
rect 10577 12223 10656 12235
rect 10686 12223 10752 12307
rect 10782 12284 10877 12307
rect 10782 12250 10794 12284
rect 10828 12250 10877 12284
rect 10782 12223 10877 12250
rect 10907 12223 10973 12307
rect 11003 12284 11141 12307
rect 11003 12250 11029 12284
rect 11063 12250 11097 12284
rect 11131 12250 11141 12284
rect 11003 12223 11141 12250
rect 11171 12284 11223 12307
rect 11171 12250 11181 12284
rect 11215 12250 11223 12284
rect 11171 12223 11223 12250
rect 11461 12284 11513 12307
rect 11461 12250 11469 12284
rect 11503 12250 11513 12284
rect 11461 12223 11513 12250
rect 11543 12284 11681 12307
rect 11543 12250 11553 12284
rect 11587 12250 11621 12284
rect 11655 12250 11681 12284
rect 11543 12223 11681 12250
rect 11711 12223 11777 12307
rect 11807 12284 11902 12307
rect 11807 12250 11856 12284
rect 11890 12250 11902 12284
rect 11807 12223 11902 12250
rect 11932 12223 11998 12307
rect 12028 12269 12107 12307
rect 12028 12235 12063 12269
rect 12097 12235 12107 12269
rect 12028 12223 12107 12235
rect 12137 12288 12189 12353
rect 12137 12254 12147 12288
rect 12181 12254 12189 12288
rect 12137 12223 12189 12254
rect 12705 12273 12763 12307
rect 12705 12239 12718 12273
rect 12752 12239 12763 12273
rect 12705 12223 12763 12239
rect 12793 12295 12849 12307
rect 12793 12261 12804 12295
rect 12838 12261 12849 12295
rect 12793 12223 12849 12261
rect 12879 12273 12935 12307
rect 12879 12239 12890 12273
rect 12924 12239 12935 12273
rect 12879 12223 12935 12239
rect 12965 12295 13021 12307
rect 12965 12261 12976 12295
rect 13010 12261 13021 12295
rect 12965 12223 13021 12261
rect 13051 12273 13118 12307
rect 13051 12239 13073 12273
rect 13107 12239 13118 12273
rect 13051 12223 13118 12239
rect 13148 12277 13201 12307
rect 13148 12243 13159 12277
rect 13193 12243 13201 12277
rect 13148 12223 13201 12243
rect 13255 12277 13308 12307
rect 13255 12243 13263 12277
rect 13297 12243 13308 12277
rect 13255 12223 13308 12243
rect 13338 12273 13405 12307
rect 13338 12239 13349 12273
rect 13383 12239 13405 12273
rect 13338 12223 13405 12239
rect 13435 12295 13491 12307
rect 13435 12261 13446 12295
rect 13480 12261 13491 12295
rect 13435 12223 13491 12261
rect 13521 12273 13577 12307
rect 13521 12239 13532 12273
rect 13566 12239 13577 12273
rect 13521 12223 13577 12239
rect 13607 12295 13663 12307
rect 13607 12261 13618 12295
rect 13652 12261 13663 12295
rect 13607 12223 13663 12261
rect 13693 12273 13751 12307
rect 13693 12239 13704 12273
rect 13738 12239 13751 12273
rect 13693 12223 13751 12239
rect 13807 12282 13859 12327
rect 13807 12248 13815 12282
rect 13849 12248 13859 12282
rect 13807 12223 13859 12248
rect 13889 12269 13947 12327
rect 13889 12235 13901 12269
rect 13935 12235 13947 12269
rect 13889 12223 13947 12235
rect 13977 12299 14029 12327
rect 14614 12307 14664 12353
rect 13977 12265 13987 12299
rect 14021 12265 14029 12299
rect 13977 12223 14029 12265
rect 14105 12295 14157 12307
rect 14105 12261 14113 12295
rect 14147 12261 14157 12295
rect 14105 12223 14157 12261
rect 14187 12269 14241 12307
rect 14187 12235 14197 12269
rect 14231 12235 14241 12269
rect 14187 12223 14241 12235
rect 14341 12295 14393 12307
rect 14341 12261 14351 12295
rect 14385 12261 14393 12295
rect 14341 12223 14393 12261
rect 14447 12295 14499 12307
rect 14447 12261 14455 12295
rect 14489 12261 14499 12295
rect 14447 12223 14499 12261
rect 14599 12269 14664 12307
rect 14599 12235 14614 12269
rect 14648 12235 14664 12269
rect 14599 12223 14664 12235
rect 14694 12295 14746 12353
rect 14694 12261 14704 12295
rect 14738 12261 14746 12295
rect 14694 12223 14746 12261
rect 15095 12295 15147 12307
rect 15095 12261 15103 12295
rect 15137 12261 15147 12295
rect 15095 12223 15147 12261
rect 15177 12269 15231 12307
rect 15177 12235 15187 12269
rect 15221 12235 15231 12269
rect 15177 12223 15231 12235
rect 15261 12295 15313 12307
rect 15261 12261 15271 12295
rect 15305 12261 15313 12295
rect 15261 12223 15313 12261
rect 15381 12265 15486 12307
rect 15381 12231 15393 12265
rect 15427 12231 15486 12265
rect 15381 12223 15486 12231
rect 15516 12295 15566 12307
rect 15997 12307 16047 12351
rect 15725 12295 15843 12307
rect 15516 12271 15581 12295
rect 15516 12237 15526 12271
rect 15560 12237 15581 12271
rect 15516 12223 15581 12237
rect 15611 12271 15677 12295
rect 15611 12237 15633 12271
rect 15667 12237 15677 12271
rect 15611 12223 15677 12237
rect 15707 12223 15843 12295
rect 15873 12223 15915 12307
rect 15945 12269 16047 12307
rect 15945 12235 15979 12269
rect 16013 12235 16047 12269
rect 15945 12223 16047 12235
rect 16077 12295 16131 12351
rect 16749 12307 16799 12353
rect 16301 12295 16351 12307
rect 16077 12265 16146 12295
rect 16077 12231 16091 12265
rect 16125 12231 16146 12265
rect 16077 12223 16146 12231
rect 16176 12269 16255 12295
rect 16176 12235 16201 12269
rect 16235 12235 16255 12269
rect 16176 12223 16255 12235
rect 16285 12223 16351 12295
rect 16381 12265 16500 12307
rect 16381 12231 16413 12265
rect 16447 12231 16500 12265
rect 16381 12223 16500 12231
rect 16530 12223 16591 12307
rect 16621 12285 16673 12307
rect 16621 12251 16631 12285
rect 16665 12251 16673 12285
rect 16621 12223 16673 12251
rect 16727 12269 16799 12307
rect 16727 12235 16755 12269
rect 16789 12235 16799 12269
rect 16727 12223 16799 12235
rect 16829 12319 16881 12353
rect 16829 12285 16839 12319
rect 16873 12285 16881 12319
rect 16829 12223 16881 12285
rect 17027 12277 17080 12307
rect 17027 12243 17035 12277
rect 17069 12243 17080 12277
rect 17027 12223 17080 12243
rect 17110 12273 17177 12307
rect 17110 12239 17121 12273
rect 17155 12239 17177 12273
rect 17110 12223 17177 12239
rect 17207 12295 17263 12307
rect 17207 12261 17218 12295
rect 17252 12261 17263 12295
rect 17207 12223 17263 12261
rect 17293 12273 17349 12307
rect 17293 12239 17304 12273
rect 17338 12239 17349 12273
rect 17293 12223 17349 12239
rect 17379 12295 17435 12307
rect 17379 12261 17390 12295
rect 17424 12261 17435 12295
rect 17379 12223 17435 12261
rect 17465 12273 17523 12307
rect 17465 12239 17476 12273
rect 17510 12239 17523 12273
rect 17763 12288 17815 12333
rect 17763 12254 17771 12288
rect 17805 12254 17815 12288
rect 17465 12223 17523 12239
rect 17763 12223 17815 12254
rect 18209 12288 18261 12333
rect 18209 12254 18219 12288
rect 18253 12254 18261 12288
rect 18209 12223 18261 12254
rect 18315 12288 18367 12333
rect 18315 12254 18323 12288
rect 18357 12254 18367 12288
rect 18315 12223 18367 12254
rect 19313 12288 19365 12333
rect 19313 12254 19323 12288
rect 19357 12254 19365 12288
rect 19313 12223 19365 12254
rect 19419 12277 19472 12307
rect 19419 12243 19427 12277
rect 19461 12243 19472 12277
rect 19419 12223 19472 12243
rect 19502 12273 19569 12307
rect 19502 12239 19513 12273
rect 19547 12239 19569 12273
rect 19502 12223 19569 12239
rect 19599 12295 19655 12307
rect 19599 12261 19610 12295
rect 19644 12261 19655 12295
rect 19599 12223 19655 12261
rect 19685 12273 19741 12307
rect 19685 12239 19696 12273
rect 19730 12239 19741 12273
rect 19685 12223 19741 12239
rect 19771 12295 19827 12307
rect 19771 12261 19782 12295
rect 19816 12261 19827 12295
rect 19771 12223 19827 12261
rect 19857 12273 19915 12307
rect 19857 12239 19868 12273
rect 19902 12239 19915 12273
rect 19857 12223 19915 12239
rect 19971 12290 20023 12333
rect 19971 12256 19979 12290
rect 20013 12256 20023 12290
rect 19971 12223 20023 12256
rect 20141 12290 20193 12333
rect 20141 12256 20151 12290
rect 20185 12256 20193 12290
rect 20141 12223 20193 12256
rect 29860 4546 29918 4558
rect 29860 4370 29872 4546
rect 29906 4370 29918 4546
rect 29860 4358 29918 4370
rect 30118 4546 30176 4558
rect 30118 4370 30130 4546
rect 30164 4370 30176 4546
rect 30118 4358 30176 4370
rect 30240 4546 30298 4558
rect 30240 4370 30252 4546
rect 30286 4370 30298 4546
rect 30240 4358 30298 4370
rect 30498 4546 30556 4558
rect 30498 4370 30510 4546
rect 30544 4370 30556 4546
rect 30498 4358 30556 4370
rect 30640 4546 30698 4558
rect 30640 4370 30652 4546
rect 30686 4370 30698 4546
rect 30640 4358 30698 4370
rect 30898 4546 30956 4558
rect 30898 4370 30910 4546
rect 30944 4370 30956 4546
rect 30898 4358 30956 4370
rect 31020 4546 31078 4558
rect 31020 4370 31032 4546
rect 31066 4370 31078 4546
rect 31020 4358 31078 4370
rect 31278 4546 31336 4558
rect 31278 4370 31290 4546
rect 31324 4370 31336 4546
rect 31278 4358 31336 4370
rect 31536 4546 31594 4558
rect 31536 4370 31548 4546
rect 31582 4370 31594 4546
rect 31536 4358 31594 4370
rect 31794 4546 31852 4558
rect 31794 4370 31806 4546
rect 31840 4370 31852 4546
rect 31794 4358 31852 4370
rect 32052 4546 32110 4558
rect 32052 4370 32064 4546
rect 32098 4370 32110 4546
rect 32052 4358 32110 4370
rect 32310 4546 32368 4558
rect 32310 4370 32322 4546
rect 32356 4370 32368 4546
rect 32310 4358 32368 4370
rect 32568 4546 32626 4558
rect 32568 4370 32580 4546
rect 32614 4370 32626 4546
rect 32568 4358 32626 4370
rect 32826 4546 32884 4558
rect 32826 4370 32838 4546
rect 32872 4370 32884 4546
rect 32826 4358 32884 4370
rect 33084 4546 33142 4558
rect 33084 4370 33096 4546
rect 33130 4370 33142 4546
rect 33084 4358 33142 4370
rect 33342 4546 33400 4558
rect 33342 4370 33354 4546
rect 33388 4370 33400 4546
rect 33342 4358 33400 4370
rect 33460 4546 33518 4558
rect 33460 4370 33472 4546
rect 33506 4370 33518 4546
rect 33460 4358 33518 4370
rect 33718 4546 33776 4558
rect 33718 4370 33730 4546
rect 33764 4370 33776 4546
rect 33718 4358 33776 4370
rect 1430 2696 1488 2708
rect 1430 1720 1442 2696
rect 1476 1720 1488 2696
rect 1430 1708 1488 1720
rect 1518 2696 1576 2708
rect 1518 1720 1530 2696
rect 1564 1720 1576 2696
rect 1630 2696 1688 2708
rect 1630 2520 1642 2696
rect 1676 2520 1688 2696
rect 1630 2508 1688 2520
rect 1718 2696 1776 2708
rect 1718 2520 1730 2696
rect 1764 2520 1776 2696
rect 1718 2508 1776 2520
rect 1843 2689 1905 2701
rect 1518 1708 1576 1720
rect 1843 1713 1855 2689
rect 1889 1713 1905 2689
rect 1843 1701 1905 1713
rect 1935 2689 2001 2701
rect 1935 1713 1951 2689
rect 1985 1713 2001 2689
rect 1935 1701 2001 1713
rect 2031 2689 2097 2701
rect 2031 1713 2047 2689
rect 2081 1713 2097 2689
rect 2031 1701 2097 1713
rect 2127 2689 2193 2701
rect 2127 1713 2143 2689
rect 2177 1713 2193 2689
rect 2127 1701 2193 1713
rect 2223 2689 2289 2701
rect 2223 1713 2239 2689
rect 2273 1713 2289 2689
rect 2223 1701 2289 1713
rect 2319 2689 2385 2701
rect 2319 1713 2335 2689
rect 2369 1713 2385 2689
rect 2319 1701 2385 1713
rect 2415 2689 2481 2701
rect 2415 1713 2431 2689
rect 2465 1713 2481 2689
rect 2415 1701 2481 1713
rect 2511 2689 2577 2701
rect 2511 1713 2527 2689
rect 2561 1713 2577 2689
rect 2511 1701 2577 1713
rect 2607 2689 2673 2701
rect 2607 1713 2623 2689
rect 2657 1713 2673 2689
rect 2607 1701 2673 1713
rect 2703 2689 2769 2701
rect 2703 1713 2719 2689
rect 2753 1713 2769 2689
rect 2703 1701 2769 1713
rect 2799 2689 2865 2701
rect 2799 1713 2815 2689
rect 2849 1713 2865 2689
rect 2799 1701 2865 1713
rect 2895 2689 2961 2701
rect 2895 1713 2911 2689
rect 2945 1713 2961 2689
rect 2895 1701 2961 1713
rect 2991 2689 3053 2701
rect 2991 1713 3007 2689
rect 3041 1713 3053 2689
rect 2991 1701 3053 1713
rect 3110 2696 3168 2708
rect 3110 1720 3122 2696
rect 3156 1720 3168 2696
rect 3110 1708 3168 1720
rect 3198 2696 3256 2708
rect 3198 1720 3210 2696
rect 3244 1720 3256 2696
rect 3198 1708 3256 1720
rect 4730 2696 4788 2708
rect 4730 1720 4742 2696
rect 4776 1720 4788 2696
rect 4730 1708 4788 1720
rect 4818 2696 4876 2708
rect 4818 1720 4830 2696
rect 4864 1720 4876 2696
rect 4930 2696 4988 2708
rect 4930 2520 4942 2696
rect 4976 2520 4988 2696
rect 4930 2508 4988 2520
rect 5018 2696 5076 2708
rect 5018 2520 5030 2696
rect 5064 2520 5076 2696
rect 5018 2508 5076 2520
rect 5143 2689 5205 2701
rect 4818 1708 4876 1720
rect 5143 1713 5155 2689
rect 5189 1713 5205 2689
rect 5143 1701 5205 1713
rect 5235 2689 5301 2701
rect 5235 1713 5251 2689
rect 5285 1713 5301 2689
rect 5235 1701 5301 1713
rect 5331 2689 5397 2701
rect 5331 1713 5347 2689
rect 5381 1713 5397 2689
rect 5331 1701 5397 1713
rect 5427 2689 5493 2701
rect 5427 1713 5443 2689
rect 5477 1713 5493 2689
rect 5427 1701 5493 1713
rect 5523 2689 5589 2701
rect 5523 1713 5539 2689
rect 5573 1713 5589 2689
rect 5523 1701 5589 1713
rect 5619 2689 5685 2701
rect 5619 1713 5635 2689
rect 5669 1713 5685 2689
rect 5619 1701 5685 1713
rect 5715 2689 5781 2701
rect 5715 1713 5731 2689
rect 5765 1713 5781 2689
rect 5715 1701 5781 1713
rect 5811 2689 5877 2701
rect 5811 1713 5827 2689
rect 5861 1713 5877 2689
rect 5811 1701 5877 1713
rect 5907 2689 5973 2701
rect 5907 1713 5923 2689
rect 5957 1713 5973 2689
rect 5907 1701 5973 1713
rect 6003 2689 6069 2701
rect 6003 1713 6019 2689
rect 6053 1713 6069 2689
rect 6003 1701 6069 1713
rect 6099 2689 6165 2701
rect 6099 1713 6115 2689
rect 6149 1713 6165 2689
rect 6099 1701 6165 1713
rect 6195 2689 6261 2701
rect 6195 1713 6211 2689
rect 6245 1713 6261 2689
rect 6195 1701 6261 1713
rect 6291 2689 6353 2701
rect 6291 1713 6307 2689
rect 6341 1713 6353 2689
rect 6291 1701 6353 1713
rect 6410 2696 6468 2708
rect 6410 1720 6422 2696
rect 6456 1720 6468 2696
rect 6410 1708 6468 1720
rect 6498 2696 6556 2708
rect 6498 1720 6510 2696
rect 6544 1720 6556 2696
rect 6498 1708 6556 1720
rect 8030 2696 8088 2708
rect 8030 1720 8042 2696
rect 8076 1720 8088 2696
rect 8030 1708 8088 1720
rect 8118 2696 8176 2708
rect 8118 1720 8130 2696
rect 8164 1720 8176 2696
rect 8230 2696 8288 2708
rect 8230 2520 8242 2696
rect 8276 2520 8288 2696
rect 8230 2508 8288 2520
rect 8318 2696 8376 2708
rect 8318 2520 8330 2696
rect 8364 2520 8376 2696
rect 8318 2508 8376 2520
rect 8443 2689 8505 2701
rect 8118 1708 8176 1720
rect 8443 1713 8455 2689
rect 8489 1713 8505 2689
rect 8443 1701 8505 1713
rect 8535 2689 8601 2701
rect 8535 1713 8551 2689
rect 8585 1713 8601 2689
rect 8535 1701 8601 1713
rect 8631 2689 8697 2701
rect 8631 1713 8647 2689
rect 8681 1713 8697 2689
rect 8631 1701 8697 1713
rect 8727 2689 8793 2701
rect 8727 1713 8743 2689
rect 8777 1713 8793 2689
rect 8727 1701 8793 1713
rect 8823 2689 8889 2701
rect 8823 1713 8839 2689
rect 8873 1713 8889 2689
rect 8823 1701 8889 1713
rect 8919 2689 8985 2701
rect 8919 1713 8935 2689
rect 8969 1713 8985 2689
rect 8919 1701 8985 1713
rect 9015 2689 9081 2701
rect 9015 1713 9031 2689
rect 9065 1713 9081 2689
rect 9015 1701 9081 1713
rect 9111 2689 9177 2701
rect 9111 1713 9127 2689
rect 9161 1713 9177 2689
rect 9111 1701 9177 1713
rect 9207 2689 9273 2701
rect 9207 1713 9223 2689
rect 9257 1713 9273 2689
rect 9207 1701 9273 1713
rect 9303 2689 9369 2701
rect 9303 1713 9319 2689
rect 9353 1713 9369 2689
rect 9303 1701 9369 1713
rect 9399 2689 9465 2701
rect 9399 1713 9415 2689
rect 9449 1713 9465 2689
rect 9399 1701 9465 1713
rect 9495 2689 9561 2701
rect 9495 1713 9511 2689
rect 9545 1713 9561 2689
rect 9495 1701 9561 1713
rect 9591 2689 9653 2701
rect 9591 1713 9607 2689
rect 9641 1713 9653 2689
rect 9591 1701 9653 1713
rect 9710 2696 9768 2708
rect 9710 1720 9722 2696
rect 9756 1720 9768 2696
rect 9710 1708 9768 1720
rect 9798 2696 9856 2708
rect 9798 1720 9810 2696
rect 9844 1720 9856 2696
rect 9798 1708 9856 1720
rect 11330 2696 11388 2708
rect 11330 1720 11342 2696
rect 11376 1720 11388 2696
rect 11330 1708 11388 1720
rect 11418 2696 11476 2708
rect 11418 1720 11430 2696
rect 11464 1720 11476 2696
rect 11530 2696 11588 2708
rect 11530 2520 11542 2696
rect 11576 2520 11588 2696
rect 11530 2508 11588 2520
rect 11618 2696 11676 2708
rect 11618 2520 11630 2696
rect 11664 2520 11676 2696
rect 11618 2508 11676 2520
rect 11743 2689 11805 2701
rect 11418 1708 11476 1720
rect 11743 1713 11755 2689
rect 11789 1713 11805 2689
rect 11743 1701 11805 1713
rect 11835 2689 11901 2701
rect 11835 1713 11851 2689
rect 11885 1713 11901 2689
rect 11835 1701 11901 1713
rect 11931 2689 11997 2701
rect 11931 1713 11947 2689
rect 11981 1713 11997 2689
rect 11931 1701 11997 1713
rect 12027 2689 12093 2701
rect 12027 1713 12043 2689
rect 12077 1713 12093 2689
rect 12027 1701 12093 1713
rect 12123 2689 12189 2701
rect 12123 1713 12139 2689
rect 12173 1713 12189 2689
rect 12123 1701 12189 1713
rect 12219 2689 12285 2701
rect 12219 1713 12235 2689
rect 12269 1713 12285 2689
rect 12219 1701 12285 1713
rect 12315 2689 12381 2701
rect 12315 1713 12331 2689
rect 12365 1713 12381 2689
rect 12315 1701 12381 1713
rect 12411 2689 12477 2701
rect 12411 1713 12427 2689
rect 12461 1713 12477 2689
rect 12411 1701 12477 1713
rect 12507 2689 12573 2701
rect 12507 1713 12523 2689
rect 12557 1713 12573 2689
rect 12507 1701 12573 1713
rect 12603 2689 12669 2701
rect 12603 1713 12619 2689
rect 12653 1713 12669 2689
rect 12603 1701 12669 1713
rect 12699 2689 12765 2701
rect 12699 1713 12715 2689
rect 12749 1713 12765 2689
rect 12699 1701 12765 1713
rect 12795 2689 12861 2701
rect 12795 1713 12811 2689
rect 12845 1713 12861 2689
rect 12795 1701 12861 1713
rect 12891 2689 12953 2701
rect 12891 1713 12907 2689
rect 12941 1713 12953 2689
rect 12891 1701 12953 1713
rect 13010 2696 13068 2708
rect 13010 1720 13022 2696
rect 13056 1720 13068 2696
rect 13010 1708 13068 1720
rect 13098 2696 13156 2708
rect 13098 1720 13110 2696
rect 13144 1720 13156 2696
rect 13098 1708 13156 1720
rect 14930 2696 14988 2708
rect 14930 1720 14942 2696
rect 14976 1720 14988 2696
rect 14930 1708 14988 1720
rect 15018 2696 15076 2708
rect 15018 1720 15030 2696
rect 15064 1720 15076 2696
rect 15130 2696 15188 2708
rect 15130 2520 15142 2696
rect 15176 2520 15188 2696
rect 15130 2508 15188 2520
rect 15218 2696 15276 2708
rect 15218 2520 15230 2696
rect 15264 2520 15276 2696
rect 15218 2508 15276 2520
rect 15343 2689 15405 2701
rect 15018 1708 15076 1720
rect 15343 1713 15355 2689
rect 15389 1713 15405 2689
rect 15343 1701 15405 1713
rect 15435 2689 15501 2701
rect 15435 1713 15451 2689
rect 15485 1713 15501 2689
rect 15435 1701 15501 1713
rect 15531 2689 15597 2701
rect 15531 1713 15547 2689
rect 15581 1713 15597 2689
rect 15531 1701 15597 1713
rect 15627 2689 15693 2701
rect 15627 1713 15643 2689
rect 15677 1713 15693 2689
rect 15627 1701 15693 1713
rect 15723 2689 15789 2701
rect 15723 1713 15739 2689
rect 15773 1713 15789 2689
rect 15723 1701 15789 1713
rect 15819 2689 15885 2701
rect 15819 1713 15835 2689
rect 15869 1713 15885 2689
rect 15819 1701 15885 1713
rect 15915 2689 15981 2701
rect 15915 1713 15931 2689
rect 15965 1713 15981 2689
rect 15915 1701 15981 1713
rect 16011 2689 16077 2701
rect 16011 1713 16027 2689
rect 16061 1713 16077 2689
rect 16011 1701 16077 1713
rect 16107 2689 16173 2701
rect 16107 1713 16123 2689
rect 16157 1713 16173 2689
rect 16107 1701 16173 1713
rect 16203 2689 16269 2701
rect 16203 1713 16219 2689
rect 16253 1713 16269 2689
rect 16203 1701 16269 1713
rect 16299 2689 16365 2701
rect 16299 1713 16315 2689
rect 16349 1713 16365 2689
rect 16299 1701 16365 1713
rect 16395 2689 16461 2701
rect 16395 1713 16411 2689
rect 16445 1713 16461 2689
rect 16395 1701 16461 1713
rect 16491 2689 16553 2701
rect 16491 1713 16507 2689
rect 16541 1713 16553 2689
rect 16491 1701 16553 1713
rect 16610 2696 16668 2708
rect 16610 1720 16622 2696
rect 16656 1720 16668 2696
rect 16610 1708 16668 1720
rect 16698 2696 16756 2708
rect 16698 1720 16710 2696
rect 16744 1720 16756 2696
rect 16698 1708 16756 1720
rect 18430 2696 18488 2708
rect 18430 1720 18442 2696
rect 18476 1720 18488 2696
rect 18430 1708 18488 1720
rect 18518 2696 18576 2708
rect 18518 1720 18530 2696
rect 18564 1720 18576 2696
rect 18630 2696 18688 2708
rect 18630 2520 18642 2696
rect 18676 2520 18688 2696
rect 18630 2508 18688 2520
rect 18718 2696 18776 2708
rect 18718 2520 18730 2696
rect 18764 2520 18776 2696
rect 18718 2508 18776 2520
rect 18843 2689 18905 2701
rect 18518 1708 18576 1720
rect 18843 1713 18855 2689
rect 18889 1713 18905 2689
rect 18843 1701 18905 1713
rect 18935 2689 19001 2701
rect 18935 1713 18951 2689
rect 18985 1713 19001 2689
rect 18935 1701 19001 1713
rect 19031 2689 19097 2701
rect 19031 1713 19047 2689
rect 19081 1713 19097 2689
rect 19031 1701 19097 1713
rect 19127 2689 19193 2701
rect 19127 1713 19143 2689
rect 19177 1713 19193 2689
rect 19127 1701 19193 1713
rect 19223 2689 19289 2701
rect 19223 1713 19239 2689
rect 19273 1713 19289 2689
rect 19223 1701 19289 1713
rect 19319 2689 19385 2701
rect 19319 1713 19335 2689
rect 19369 1713 19385 2689
rect 19319 1701 19385 1713
rect 19415 2689 19481 2701
rect 19415 1713 19431 2689
rect 19465 1713 19481 2689
rect 19415 1701 19481 1713
rect 19511 2689 19577 2701
rect 19511 1713 19527 2689
rect 19561 1713 19577 2689
rect 19511 1701 19577 1713
rect 19607 2689 19673 2701
rect 19607 1713 19623 2689
rect 19657 1713 19673 2689
rect 19607 1701 19673 1713
rect 19703 2689 19769 2701
rect 19703 1713 19719 2689
rect 19753 1713 19769 2689
rect 19703 1701 19769 1713
rect 19799 2689 19865 2701
rect 19799 1713 19815 2689
rect 19849 1713 19865 2689
rect 19799 1701 19865 1713
rect 19895 2689 19961 2701
rect 19895 1713 19911 2689
rect 19945 1713 19961 2689
rect 19895 1701 19961 1713
rect 19991 2689 20053 2701
rect 19991 1713 20007 2689
rect 20041 1713 20053 2689
rect 19991 1701 20053 1713
rect 20110 2696 20168 2708
rect 20110 1720 20122 2696
rect 20156 1720 20168 2696
rect 20110 1708 20168 1720
rect 20198 2696 20256 2708
rect 20198 1720 20210 2696
rect 20244 1720 20256 2696
rect 20198 1708 20256 1720
rect 22130 2696 22188 2708
rect 22130 1720 22142 2696
rect 22176 1720 22188 2696
rect 22130 1708 22188 1720
rect 22218 2696 22276 2708
rect 22218 1720 22230 2696
rect 22264 1720 22276 2696
rect 22330 2696 22388 2708
rect 22330 2520 22342 2696
rect 22376 2520 22388 2696
rect 22330 2508 22388 2520
rect 22418 2696 22476 2708
rect 22418 2520 22430 2696
rect 22464 2520 22476 2696
rect 22418 2508 22476 2520
rect 22543 2689 22605 2701
rect 22218 1708 22276 1720
rect 22543 1713 22555 2689
rect 22589 1713 22605 2689
rect 22543 1701 22605 1713
rect 22635 2689 22701 2701
rect 22635 1713 22651 2689
rect 22685 1713 22701 2689
rect 22635 1701 22701 1713
rect 22731 2689 22797 2701
rect 22731 1713 22747 2689
rect 22781 1713 22797 2689
rect 22731 1701 22797 1713
rect 22827 2689 22893 2701
rect 22827 1713 22843 2689
rect 22877 1713 22893 2689
rect 22827 1701 22893 1713
rect 22923 2689 22989 2701
rect 22923 1713 22939 2689
rect 22973 1713 22989 2689
rect 22923 1701 22989 1713
rect 23019 2689 23085 2701
rect 23019 1713 23035 2689
rect 23069 1713 23085 2689
rect 23019 1701 23085 1713
rect 23115 2689 23181 2701
rect 23115 1713 23131 2689
rect 23165 1713 23181 2689
rect 23115 1701 23181 1713
rect 23211 2689 23277 2701
rect 23211 1713 23227 2689
rect 23261 1713 23277 2689
rect 23211 1701 23277 1713
rect 23307 2689 23373 2701
rect 23307 1713 23323 2689
rect 23357 1713 23373 2689
rect 23307 1701 23373 1713
rect 23403 2689 23469 2701
rect 23403 1713 23419 2689
rect 23453 1713 23469 2689
rect 23403 1701 23469 1713
rect 23499 2689 23565 2701
rect 23499 1713 23515 2689
rect 23549 1713 23565 2689
rect 23499 1701 23565 1713
rect 23595 2689 23661 2701
rect 23595 1713 23611 2689
rect 23645 1713 23661 2689
rect 23595 1701 23661 1713
rect 23691 2689 23753 2701
rect 23691 1713 23707 2689
rect 23741 1713 23753 2689
rect 23691 1701 23753 1713
rect 23810 2696 23868 2708
rect 23810 1720 23822 2696
rect 23856 1720 23868 2696
rect 23810 1708 23868 1720
rect 23898 2696 23956 2708
rect 23898 1720 23910 2696
rect 23944 1720 23956 2696
rect 23898 1708 23956 1720
rect 25930 2696 25988 2708
rect 25930 1720 25942 2696
rect 25976 1720 25988 2696
rect 25930 1708 25988 1720
rect 26018 2696 26076 2708
rect 26018 1720 26030 2696
rect 26064 1720 26076 2696
rect 26130 2696 26188 2708
rect 26130 2520 26142 2696
rect 26176 2520 26188 2696
rect 26130 2508 26188 2520
rect 26218 2696 26276 2708
rect 26218 2520 26230 2696
rect 26264 2520 26276 2696
rect 26218 2508 26276 2520
rect 26343 2689 26405 2701
rect 26018 1708 26076 1720
rect 26343 1713 26355 2689
rect 26389 1713 26405 2689
rect 26343 1701 26405 1713
rect 26435 2689 26501 2701
rect 26435 1713 26451 2689
rect 26485 1713 26501 2689
rect 26435 1701 26501 1713
rect 26531 2689 26597 2701
rect 26531 1713 26547 2689
rect 26581 1713 26597 2689
rect 26531 1701 26597 1713
rect 26627 2689 26693 2701
rect 26627 1713 26643 2689
rect 26677 1713 26693 2689
rect 26627 1701 26693 1713
rect 26723 2689 26789 2701
rect 26723 1713 26739 2689
rect 26773 1713 26789 2689
rect 26723 1701 26789 1713
rect 26819 2689 26885 2701
rect 26819 1713 26835 2689
rect 26869 1713 26885 2689
rect 26819 1701 26885 1713
rect 26915 2689 26981 2701
rect 26915 1713 26931 2689
rect 26965 1713 26981 2689
rect 26915 1701 26981 1713
rect 27011 2689 27077 2701
rect 27011 1713 27027 2689
rect 27061 1713 27077 2689
rect 27011 1701 27077 1713
rect 27107 2689 27173 2701
rect 27107 1713 27123 2689
rect 27157 1713 27173 2689
rect 27107 1701 27173 1713
rect 27203 2689 27269 2701
rect 27203 1713 27219 2689
rect 27253 1713 27269 2689
rect 27203 1701 27269 1713
rect 27299 2689 27365 2701
rect 27299 1713 27315 2689
rect 27349 1713 27365 2689
rect 27299 1701 27365 1713
rect 27395 2689 27461 2701
rect 27395 1713 27411 2689
rect 27445 1713 27461 2689
rect 27395 1701 27461 1713
rect 27491 2689 27553 2701
rect 27491 1713 27507 2689
rect 27541 1713 27553 2689
rect 27491 1701 27553 1713
rect 27610 2696 27668 2708
rect 27610 1720 27622 2696
rect 27656 1720 27668 2696
rect 27610 1708 27668 1720
rect 27698 2696 27756 2708
rect 27698 1720 27710 2696
rect 27744 1720 27756 2696
rect 27698 1708 27756 1720
<< pdiff >>
rect 4975 27052 5027 27085
rect 4975 27018 4983 27052
rect 5017 27018 5027 27052
rect 4975 26957 5027 27018
rect 4975 26923 4983 26957
rect 5017 26923 5027 26957
rect 4975 26911 5027 26923
rect 5145 27052 5197 27085
rect 5145 27018 5155 27052
rect 5189 27018 5197 27052
rect 5145 26957 5197 27018
rect 5145 26923 5155 26957
rect 5189 26923 5197 26957
rect 5145 26911 5197 26923
rect 5251 27052 5303 27085
rect 5251 27018 5259 27052
rect 5293 27018 5303 27052
rect 5251 26957 5303 27018
rect 5251 26923 5259 26957
rect 5293 26923 5303 26957
rect 5251 26911 5303 26923
rect 5421 27052 5473 27085
rect 5421 27018 5431 27052
rect 5465 27018 5473 27052
rect 5421 26957 5473 27018
rect 5421 26923 5431 26957
rect 5465 26923 5473 26957
rect 5421 26911 5473 26923
rect 5528 27039 5588 27111
rect 5528 27005 5543 27039
rect 5577 27005 5588 27039
rect 5528 26971 5588 27005
rect 5528 26937 5543 26971
rect 5577 26937 5588 26971
rect 5528 26911 5588 26937
rect 5618 27101 5674 27111
rect 5618 27067 5629 27101
rect 5663 27067 5674 27101
rect 5618 27033 5674 27067
rect 5618 26999 5629 27033
rect 5663 26999 5674 27033
rect 5618 26965 5674 26999
rect 5618 26931 5629 26965
rect 5663 26931 5674 26965
rect 5618 26911 5674 26931
rect 5704 26957 5760 27111
rect 5704 26923 5715 26957
rect 5749 26923 5760 26957
rect 5704 26911 5760 26923
rect 5790 26992 5846 27111
rect 5790 26958 5801 26992
rect 5835 26958 5846 26992
rect 5790 26911 5846 26958
rect 5876 27025 5942 27111
rect 5876 26991 5897 27025
rect 5931 26991 5942 27025
rect 5876 26957 5942 26991
rect 5876 26923 5897 26957
rect 5931 26923 5942 26957
rect 5876 26911 5942 26923
rect 5972 27087 6025 27111
rect 5972 27053 5983 27087
rect 6017 27053 6025 27087
rect 5972 26965 6025 27053
rect 5972 26931 5983 26965
rect 6017 26931 6025 26965
rect 5972 26911 6025 26931
rect 6171 26957 6223 27085
rect 6171 26923 6179 26957
rect 6213 26923 6223 26957
rect 6171 26911 6223 26923
rect 7169 26957 7221 27085
rect 7169 26923 7179 26957
rect 7213 26923 7221 26957
rect 7367 27052 7419 27085
rect 7367 27018 7375 27052
rect 7409 27018 7419 27052
rect 7367 26957 7419 27018
rect 7169 26911 7221 26923
rect 7367 26923 7375 26957
rect 7409 26923 7419 26957
rect 7367 26911 7419 26923
rect 7537 27052 7589 27085
rect 7537 27018 7547 27052
rect 7581 27018 7589 27052
rect 7537 26957 7589 27018
rect 7537 26923 7547 26957
rect 7581 26923 7589 26957
rect 7537 26911 7589 26923
rect 7643 26957 7695 27085
rect 7643 26923 7651 26957
rect 7685 26923 7695 26957
rect 7643 26911 7695 26923
rect 8641 26957 8693 27085
rect 8641 26923 8651 26957
rect 8685 26923 8693 26957
rect 8641 26911 8693 26923
rect 8747 26957 8799 27085
rect 8747 26923 8755 26957
rect 8789 26923 8799 26957
rect 8747 26911 8799 26923
rect 9745 26957 9797 27085
rect 9745 26923 9755 26957
rect 9789 26923 9797 26957
rect 10127 27033 10179 27069
rect 10127 26999 10135 27033
rect 10169 26999 10179 27033
rect 10127 26965 10179 26999
rect 10127 26931 10135 26965
rect 10169 26931 10179 26965
rect 9745 26911 9797 26923
rect 10127 26911 10179 26931
rect 10209 27033 10267 27069
rect 10209 26999 10221 27033
rect 10255 26999 10267 27033
rect 10209 26965 10267 26999
rect 10209 26931 10221 26965
rect 10255 26931 10267 26965
rect 10209 26911 10267 26931
rect 10297 27046 10349 27069
rect 10297 27012 10307 27046
rect 10341 27012 10349 27046
rect 10297 26965 10349 27012
rect 10297 26931 10307 26965
rect 10341 26931 10349 26965
rect 10297 26911 10349 26931
rect 10587 27059 10639 27085
rect 10587 27025 10595 27059
rect 10629 27025 10639 27059
rect 10587 26957 10639 27025
rect 10587 26923 10595 26957
rect 10629 26923 10639 26957
rect 10587 26911 10639 26923
rect 11217 27059 11269 27085
rect 11217 27025 11227 27059
rect 11261 27025 11269 27059
rect 11217 26957 11269 27025
rect 11217 26923 11227 26957
rect 11261 26923 11269 26957
rect 11217 26911 11269 26923
rect 11323 26957 11375 27085
rect 11323 26923 11331 26957
rect 11365 26923 11375 26957
rect 11323 26911 11375 26923
rect 12321 26957 12373 27085
rect 12321 26923 12331 26957
rect 12365 26923 12373 26957
rect 12519 27052 12571 27085
rect 12519 27018 12527 27052
rect 12561 27018 12571 27052
rect 12519 26957 12571 27018
rect 12321 26911 12373 26923
rect 12519 26923 12527 26957
rect 12561 26923 12571 26957
rect 12519 26911 12571 26923
rect 12689 27052 12741 27085
rect 12689 27018 12699 27052
rect 12733 27018 12741 27052
rect 12689 26957 12741 27018
rect 12689 26923 12699 26957
rect 12733 26923 12741 26957
rect 12689 26911 12741 26923
rect 12795 26957 12847 27085
rect 12795 26923 12803 26957
rect 12837 26923 12847 26957
rect 12795 26911 12847 26923
rect 13793 26957 13845 27085
rect 13793 26923 13803 26957
rect 13837 26923 13845 26957
rect 13793 26911 13845 26923
rect 13899 26957 13951 27085
rect 13899 26923 13907 26957
rect 13941 26923 13951 26957
rect 13899 26911 13951 26923
rect 14897 26957 14949 27085
rect 14897 26923 14907 26957
rect 14941 26923 14949 26957
rect 15095 27052 15147 27085
rect 15095 27018 15103 27052
rect 15137 27018 15147 27052
rect 15095 26957 15147 27018
rect 14897 26911 14949 26923
rect 15095 26923 15103 26957
rect 15137 26923 15147 26957
rect 15095 26911 15147 26923
rect 15265 27052 15317 27085
rect 15265 27018 15275 27052
rect 15309 27018 15317 27052
rect 15265 26957 15317 27018
rect 15265 26923 15275 26957
rect 15309 26923 15317 26957
rect 15265 26911 15317 26923
rect 15371 26957 15423 27085
rect 15371 26923 15379 26957
rect 15413 26923 15423 26957
rect 15371 26911 15423 26923
rect 16369 26957 16421 27085
rect 16369 26923 16379 26957
rect 16413 26923 16421 26957
rect 16369 26911 16421 26923
rect 16475 26957 16527 27085
rect 16475 26923 16483 26957
rect 16517 26923 16527 26957
rect 16475 26911 16527 26923
rect 17473 26957 17525 27085
rect 17473 26923 17483 26957
rect 17517 26923 17525 26957
rect 17763 27059 17815 27085
rect 17763 27025 17771 27059
rect 17805 27025 17815 27059
rect 17763 26957 17815 27025
rect 17473 26911 17525 26923
rect 17763 26923 17771 26957
rect 17805 26923 17815 26957
rect 17763 26911 17815 26923
rect 18393 27059 18445 27085
rect 18393 27025 18403 27059
rect 18437 27025 18445 27059
rect 18393 26957 18445 27025
rect 18393 26923 18403 26957
rect 18437 26923 18445 26957
rect 18393 26911 18445 26923
rect 18500 27039 18560 27111
rect 18500 27005 18515 27039
rect 18549 27005 18560 27039
rect 18500 26971 18560 27005
rect 18500 26937 18515 26971
rect 18549 26937 18560 26971
rect 18500 26911 18560 26937
rect 18590 27101 18646 27111
rect 18590 27067 18601 27101
rect 18635 27067 18646 27101
rect 18590 27033 18646 27067
rect 18590 26999 18601 27033
rect 18635 26999 18646 27033
rect 18590 26965 18646 26999
rect 18590 26931 18601 26965
rect 18635 26931 18646 26965
rect 18590 26911 18646 26931
rect 18676 26957 18732 27111
rect 18676 26923 18687 26957
rect 18721 26923 18732 26957
rect 18676 26911 18732 26923
rect 18762 26992 18818 27111
rect 18762 26958 18773 26992
rect 18807 26958 18818 26992
rect 18762 26911 18818 26958
rect 18848 27025 18914 27111
rect 18848 26991 18869 27025
rect 18903 26991 18914 27025
rect 18848 26957 18914 26991
rect 18848 26923 18869 26957
rect 18903 26923 18914 26957
rect 18848 26911 18914 26923
rect 18944 27087 18997 27111
rect 18944 27053 18955 27087
rect 18989 27053 18997 27087
rect 18944 26965 18997 27053
rect 18944 26931 18955 26965
rect 18989 26931 18997 26965
rect 18944 26911 18997 26931
rect 19235 27059 19287 27085
rect 19235 27025 19243 27059
rect 19277 27025 19287 27059
rect 19235 26957 19287 27025
rect 19235 26923 19243 26957
rect 19277 26923 19287 26957
rect 19235 26911 19287 26923
rect 19865 27059 19917 27085
rect 19865 27025 19875 27059
rect 19909 27025 19917 27059
rect 19865 26957 19917 27025
rect 19865 26923 19875 26957
rect 19909 26923 19917 26957
rect 19865 26911 19917 26923
rect 19971 27052 20023 27085
rect 19971 27018 19979 27052
rect 20013 27018 20023 27052
rect 19971 26957 20023 27018
rect 19971 26923 19979 26957
rect 20013 26923 20023 26957
rect 19971 26911 20023 26923
rect 20141 27052 20193 27085
rect 20141 27018 20151 27052
rect 20185 27018 20193 27052
rect 20141 26957 20193 27018
rect 20141 26923 20151 26957
rect 20185 26923 20193 26957
rect 20141 26911 20193 26923
rect 4975 26805 5027 26817
rect 4975 26771 4983 26805
rect 5017 26771 5027 26805
rect 4975 26710 5027 26771
rect 4975 26676 4983 26710
rect 5017 26676 5027 26710
rect 4975 26643 5027 26676
rect 5145 26805 5197 26817
rect 5145 26771 5155 26805
rect 5189 26771 5197 26805
rect 5145 26710 5197 26771
rect 5145 26676 5155 26710
rect 5189 26676 5197 26710
rect 5145 26643 5197 26676
rect 5435 26805 5487 26817
rect 5435 26771 5443 26805
rect 5477 26771 5487 26805
rect 5435 26703 5487 26771
rect 5435 26669 5443 26703
rect 5477 26669 5487 26703
rect 5435 26643 5487 26669
rect 6065 26805 6117 26817
rect 6065 26771 6075 26805
rect 6109 26771 6117 26805
rect 6065 26703 6117 26771
rect 6065 26669 6075 26703
rect 6109 26669 6117 26703
rect 6065 26643 6117 26669
rect 6171 26805 6223 26817
rect 6171 26771 6179 26805
rect 6213 26771 6223 26805
rect 6171 26643 6223 26771
rect 7169 26805 7221 26817
rect 7169 26771 7179 26805
rect 7213 26771 7221 26805
rect 7459 26805 7511 26817
rect 7169 26643 7221 26771
rect 7459 26771 7467 26805
rect 7501 26771 7511 26805
rect 7459 26703 7511 26771
rect 7459 26669 7467 26703
rect 7501 26669 7511 26703
rect 7459 26643 7511 26669
rect 7905 26805 7957 26817
rect 7905 26771 7915 26805
rect 7949 26771 7957 26805
rect 7905 26703 7957 26771
rect 7905 26669 7915 26703
rect 7949 26669 7957 26703
rect 7905 26643 7957 26669
rect 8011 26805 8063 26817
rect 8011 26771 8019 26805
rect 8053 26771 8063 26805
rect 8011 26643 8063 26771
rect 9009 26805 9061 26817
rect 9009 26771 9019 26805
rect 9053 26771 9061 26805
rect 9009 26643 9061 26771
rect 9115 26805 9167 26817
rect 9115 26771 9123 26805
rect 9157 26771 9167 26805
rect 9115 26643 9167 26771
rect 10113 26805 10165 26817
rect 10113 26771 10123 26805
rect 10157 26771 10165 26805
rect 10113 26643 10165 26771
rect 10219 26805 10271 26817
rect 10219 26771 10227 26805
rect 10261 26771 10271 26805
rect 10219 26643 10271 26771
rect 11217 26805 11269 26817
rect 11217 26771 11227 26805
rect 11261 26771 11269 26805
rect 11217 26643 11269 26771
rect 11323 26805 11375 26817
rect 11323 26771 11331 26805
rect 11365 26771 11375 26805
rect 11323 26643 11375 26771
rect 12321 26805 12373 26817
rect 12321 26771 12331 26805
rect 12365 26771 12373 26805
rect 12611 26805 12663 26817
rect 12321 26643 12373 26771
rect 12611 26771 12619 26805
rect 12653 26771 12663 26805
rect 12611 26703 12663 26771
rect 12611 26669 12619 26703
rect 12653 26669 12663 26703
rect 12611 26643 12663 26669
rect 13057 26805 13109 26817
rect 13057 26771 13067 26805
rect 13101 26771 13109 26805
rect 13057 26703 13109 26771
rect 13057 26669 13067 26703
rect 13101 26669 13109 26703
rect 13057 26643 13109 26669
rect 13163 26805 13215 26817
rect 13163 26771 13171 26805
rect 13205 26771 13215 26805
rect 13163 26643 13215 26771
rect 14161 26805 14213 26817
rect 14161 26771 14171 26805
rect 14205 26771 14213 26805
rect 14161 26643 14213 26771
rect 14267 26805 14319 26817
rect 14267 26771 14275 26805
rect 14309 26771 14319 26805
rect 14267 26643 14319 26771
rect 15265 26805 15317 26817
rect 15265 26771 15275 26805
rect 15309 26771 15317 26805
rect 15265 26643 15317 26771
rect 15371 26805 15423 26817
rect 15371 26771 15379 26805
rect 15413 26771 15423 26805
rect 15371 26643 15423 26771
rect 16369 26805 16421 26817
rect 16369 26771 16379 26805
rect 16413 26771 16421 26805
rect 16369 26643 16421 26771
rect 16475 26805 16527 26817
rect 16475 26771 16483 26805
rect 16517 26771 16527 26805
rect 16475 26643 16527 26771
rect 17473 26805 17525 26817
rect 17473 26771 17483 26805
rect 17517 26771 17525 26805
rect 17763 26805 17815 26817
rect 17473 26643 17525 26771
rect 17763 26771 17771 26805
rect 17805 26771 17815 26805
rect 17763 26643 17815 26771
rect 18761 26805 18813 26817
rect 18761 26771 18771 26805
rect 18805 26771 18813 26805
rect 18761 26643 18813 26771
rect 18867 26805 18919 26817
rect 18867 26771 18875 26805
rect 18909 26771 18919 26805
rect 18867 26643 18919 26771
rect 19865 26805 19917 26817
rect 19865 26771 19875 26805
rect 19909 26771 19917 26805
rect 19865 26643 19917 26771
rect 19971 26805 20023 26817
rect 19971 26771 19979 26805
rect 20013 26771 20023 26805
rect 19971 26710 20023 26771
rect 19971 26676 19979 26710
rect 20013 26676 20023 26710
rect 19971 26643 20023 26676
rect 20141 26805 20193 26817
rect 20141 26771 20151 26805
rect 20185 26771 20193 26805
rect 20141 26710 20193 26771
rect 20141 26676 20151 26710
rect 20185 26676 20193 26710
rect 20141 26643 20193 26676
rect 4975 25964 5027 25997
rect 4975 25930 4983 25964
rect 5017 25930 5027 25964
rect 4975 25869 5027 25930
rect 4975 25835 4983 25869
rect 5017 25835 5027 25869
rect 4975 25823 5027 25835
rect 5145 25964 5197 25997
rect 5145 25930 5155 25964
rect 5189 25930 5197 25964
rect 5145 25869 5197 25930
rect 5145 25835 5155 25869
rect 5189 25835 5197 25869
rect 5145 25823 5197 25835
rect 5435 25869 5487 25997
rect 5435 25835 5443 25869
rect 5477 25835 5487 25869
rect 5435 25823 5487 25835
rect 6433 25869 6485 25997
rect 6433 25835 6443 25869
rect 6477 25835 6485 25869
rect 6433 25823 6485 25835
rect 6539 25869 6591 25997
rect 6539 25835 6547 25869
rect 6581 25835 6591 25869
rect 6539 25823 6591 25835
rect 7537 25869 7589 25997
rect 7537 25835 7547 25869
rect 7581 25835 7589 25869
rect 7537 25823 7589 25835
rect 7643 25869 7695 25997
rect 7643 25835 7651 25869
rect 7685 25835 7695 25869
rect 7643 25823 7695 25835
rect 8641 25869 8693 25997
rect 8641 25835 8651 25869
rect 8685 25835 8693 25869
rect 8641 25823 8693 25835
rect 8747 25869 8799 25997
rect 8747 25835 8755 25869
rect 8789 25835 8799 25869
rect 8747 25823 8799 25835
rect 9745 25869 9797 25997
rect 9745 25835 9755 25869
rect 9789 25835 9797 25869
rect 10035 25971 10087 25997
rect 10035 25937 10043 25971
rect 10077 25937 10087 25971
rect 10035 25869 10087 25937
rect 9745 25823 9797 25835
rect 10035 25835 10043 25869
rect 10077 25835 10087 25869
rect 10035 25823 10087 25835
rect 10481 25971 10533 25997
rect 10481 25937 10491 25971
rect 10525 25937 10533 25971
rect 10481 25869 10533 25937
rect 10481 25835 10491 25869
rect 10525 25835 10533 25869
rect 10481 25823 10533 25835
rect 10587 25869 10639 25997
rect 10587 25835 10595 25869
rect 10629 25835 10639 25869
rect 10587 25823 10639 25835
rect 11585 25869 11637 25997
rect 11585 25835 11595 25869
rect 11629 25835 11637 25869
rect 11585 25823 11637 25835
rect 11691 25869 11743 25997
rect 11691 25835 11699 25869
rect 11733 25835 11743 25869
rect 11691 25823 11743 25835
rect 12689 25869 12741 25997
rect 12689 25835 12699 25869
rect 12733 25835 12741 25869
rect 12689 25823 12741 25835
rect 12795 25869 12847 25997
rect 12795 25835 12803 25869
rect 12837 25835 12847 25869
rect 12795 25823 12847 25835
rect 13793 25869 13845 25997
rect 13793 25835 13803 25869
rect 13837 25835 13845 25869
rect 13793 25823 13845 25835
rect 13899 25869 13951 25997
rect 13899 25835 13907 25869
rect 13941 25835 13951 25869
rect 13899 25823 13951 25835
rect 14897 25869 14949 25997
rect 14897 25835 14907 25869
rect 14941 25835 14949 25869
rect 15187 25971 15239 25997
rect 15187 25937 15195 25971
rect 15229 25937 15239 25971
rect 15187 25869 15239 25937
rect 14897 25823 14949 25835
rect 15187 25835 15195 25869
rect 15229 25835 15239 25869
rect 15187 25823 15239 25835
rect 15449 25971 15501 25997
rect 15449 25937 15459 25971
rect 15493 25937 15501 25971
rect 15449 25869 15501 25937
rect 15449 25835 15459 25869
rect 15493 25835 15501 25869
rect 15449 25823 15501 25835
rect 15555 25869 15607 25997
rect 15555 25835 15563 25869
rect 15597 25835 15607 25869
rect 15555 25823 15607 25835
rect 16553 25869 16605 25997
rect 16553 25835 16563 25869
rect 16597 25835 16605 25869
rect 16553 25823 16605 25835
rect 16659 25869 16711 25997
rect 16659 25835 16667 25869
rect 16701 25835 16711 25869
rect 16659 25823 16711 25835
rect 17657 25869 17709 25997
rect 17657 25835 17667 25869
rect 17701 25835 17709 25869
rect 17657 25823 17709 25835
rect 17763 25869 17815 25997
rect 17763 25835 17771 25869
rect 17805 25835 17815 25869
rect 17763 25823 17815 25835
rect 18761 25869 18813 25997
rect 18761 25835 18771 25869
rect 18805 25835 18813 25869
rect 18761 25823 18813 25835
rect 18867 25869 18919 25997
rect 18867 25835 18875 25869
rect 18909 25835 18919 25869
rect 18867 25823 18919 25835
rect 19865 25869 19917 25997
rect 19865 25835 19875 25869
rect 19909 25835 19917 25869
rect 19865 25823 19917 25835
rect 19971 25964 20023 25997
rect 19971 25930 19979 25964
rect 20013 25930 20023 25964
rect 19971 25869 20023 25930
rect 19971 25835 19979 25869
rect 20013 25835 20023 25869
rect 19971 25823 20023 25835
rect 20141 25964 20193 25997
rect 20141 25930 20151 25964
rect 20185 25930 20193 25964
rect 20141 25869 20193 25930
rect 20141 25835 20151 25869
rect 20185 25835 20193 25869
rect 20141 25823 20193 25835
rect 4975 25717 5027 25729
rect 4975 25683 4983 25717
rect 5017 25683 5027 25717
rect 4975 25622 5027 25683
rect 4975 25588 4983 25622
rect 5017 25588 5027 25622
rect 4975 25555 5027 25588
rect 5145 25717 5197 25729
rect 5145 25683 5155 25717
rect 5189 25683 5197 25717
rect 5145 25622 5197 25683
rect 5145 25588 5155 25622
rect 5189 25588 5197 25622
rect 5145 25555 5197 25588
rect 5435 25717 5487 25729
rect 5435 25683 5443 25717
rect 5477 25683 5487 25717
rect 5435 25615 5487 25683
rect 5435 25581 5443 25615
rect 5477 25581 5487 25615
rect 5435 25555 5487 25581
rect 6065 25717 6117 25729
rect 6065 25683 6075 25717
rect 6109 25683 6117 25717
rect 6065 25615 6117 25683
rect 6065 25581 6075 25615
rect 6109 25581 6117 25615
rect 6065 25555 6117 25581
rect 6171 25717 6223 25729
rect 6171 25683 6179 25717
rect 6213 25683 6223 25717
rect 6171 25555 6223 25683
rect 7169 25717 7221 25729
rect 7169 25683 7179 25717
rect 7213 25683 7221 25717
rect 7459 25717 7511 25729
rect 7169 25555 7221 25683
rect 7459 25683 7467 25717
rect 7501 25683 7511 25717
rect 7459 25615 7511 25683
rect 7459 25581 7467 25615
rect 7501 25581 7511 25615
rect 7459 25555 7511 25581
rect 7905 25717 7957 25729
rect 7905 25683 7915 25717
rect 7949 25683 7957 25717
rect 7905 25615 7957 25683
rect 7905 25581 7915 25615
rect 7949 25581 7957 25615
rect 7905 25555 7957 25581
rect 8011 25717 8063 25729
rect 8011 25683 8019 25717
rect 8053 25683 8063 25717
rect 8011 25555 8063 25683
rect 9009 25717 9061 25729
rect 9009 25683 9019 25717
rect 9053 25683 9061 25717
rect 9009 25555 9061 25683
rect 9115 25717 9167 25729
rect 9115 25683 9123 25717
rect 9157 25683 9167 25717
rect 9115 25555 9167 25683
rect 10113 25717 10165 25729
rect 10113 25683 10123 25717
rect 10157 25683 10165 25717
rect 10113 25555 10165 25683
rect 10219 25717 10271 25729
rect 10219 25683 10227 25717
rect 10261 25683 10271 25717
rect 10219 25555 10271 25683
rect 11217 25717 11269 25729
rect 11217 25683 11227 25717
rect 11261 25683 11269 25717
rect 11217 25555 11269 25683
rect 11323 25717 11375 25729
rect 11323 25683 11331 25717
rect 11365 25683 11375 25717
rect 11323 25555 11375 25683
rect 12321 25717 12373 25729
rect 12321 25683 12331 25717
rect 12365 25683 12373 25717
rect 12611 25717 12663 25729
rect 12321 25555 12373 25683
rect 12611 25683 12619 25717
rect 12653 25683 12663 25717
rect 12611 25615 12663 25683
rect 12611 25581 12619 25615
rect 12653 25581 12663 25615
rect 12611 25555 12663 25581
rect 13057 25717 13109 25729
rect 13057 25683 13067 25717
rect 13101 25683 13109 25717
rect 13057 25615 13109 25683
rect 13057 25581 13067 25615
rect 13101 25581 13109 25615
rect 13057 25555 13109 25581
rect 13163 25717 13215 25729
rect 13163 25683 13171 25717
rect 13205 25683 13215 25717
rect 13163 25555 13215 25683
rect 14161 25717 14213 25729
rect 14161 25683 14171 25717
rect 14205 25683 14213 25717
rect 14161 25555 14213 25683
rect 14267 25717 14319 25729
rect 14267 25683 14275 25717
rect 14309 25683 14319 25717
rect 14267 25555 14319 25683
rect 15265 25717 15317 25729
rect 15265 25683 15275 25717
rect 15309 25683 15317 25717
rect 15265 25555 15317 25683
rect 15371 25717 15423 25729
rect 15371 25683 15379 25717
rect 15413 25683 15423 25717
rect 15371 25555 15423 25683
rect 16369 25717 16421 25729
rect 16369 25683 16379 25717
rect 16413 25683 16421 25717
rect 16369 25555 16421 25683
rect 16475 25717 16527 25729
rect 16475 25683 16483 25717
rect 16517 25683 16527 25717
rect 16475 25555 16527 25683
rect 17473 25717 17525 25729
rect 17473 25683 17483 25717
rect 17517 25683 17525 25717
rect 17763 25717 17815 25729
rect 17473 25555 17525 25683
rect 17763 25683 17771 25717
rect 17805 25683 17815 25717
rect 17763 25555 17815 25683
rect 18761 25717 18813 25729
rect 18761 25683 18771 25717
rect 18805 25683 18813 25717
rect 18761 25555 18813 25683
rect 18867 25717 18919 25729
rect 18867 25683 18875 25717
rect 18909 25683 18919 25717
rect 18867 25555 18919 25683
rect 19865 25717 19917 25729
rect 19865 25683 19875 25717
rect 19909 25683 19917 25717
rect 19865 25555 19917 25683
rect 19971 25717 20023 25729
rect 19971 25683 19979 25717
rect 20013 25683 20023 25717
rect 19971 25622 20023 25683
rect 19971 25588 19979 25622
rect 20013 25588 20023 25622
rect 19971 25555 20023 25588
rect 20141 25717 20193 25729
rect 20141 25683 20151 25717
rect 20185 25683 20193 25717
rect 20141 25622 20193 25683
rect 20141 25588 20151 25622
rect 20185 25588 20193 25622
rect 20141 25555 20193 25588
rect 4975 24876 5027 24909
rect 4975 24842 4983 24876
rect 5017 24842 5027 24876
rect 4975 24781 5027 24842
rect 4975 24747 4983 24781
rect 5017 24747 5027 24781
rect 4975 24735 5027 24747
rect 5145 24876 5197 24909
rect 5145 24842 5155 24876
rect 5189 24842 5197 24876
rect 5145 24781 5197 24842
rect 5145 24747 5155 24781
rect 5189 24747 5197 24781
rect 5145 24735 5197 24747
rect 5435 24781 5487 24909
rect 5435 24747 5443 24781
rect 5477 24747 5487 24781
rect 5435 24735 5487 24747
rect 6433 24781 6485 24909
rect 6433 24747 6443 24781
rect 6477 24747 6485 24781
rect 6433 24735 6485 24747
rect 6539 24781 6591 24909
rect 6539 24747 6547 24781
rect 6581 24747 6591 24781
rect 6539 24735 6591 24747
rect 7537 24781 7589 24909
rect 7537 24747 7547 24781
rect 7581 24747 7589 24781
rect 7537 24735 7589 24747
rect 7643 24781 7695 24909
rect 7643 24747 7651 24781
rect 7685 24747 7695 24781
rect 7643 24735 7695 24747
rect 8641 24781 8693 24909
rect 8641 24747 8651 24781
rect 8685 24747 8693 24781
rect 8641 24735 8693 24747
rect 8747 24781 8799 24909
rect 8747 24747 8755 24781
rect 8789 24747 8799 24781
rect 8747 24735 8799 24747
rect 9745 24781 9797 24909
rect 9745 24747 9755 24781
rect 9789 24747 9797 24781
rect 10035 24883 10087 24909
rect 10035 24849 10043 24883
rect 10077 24849 10087 24883
rect 10035 24781 10087 24849
rect 9745 24735 9797 24747
rect 10035 24747 10043 24781
rect 10077 24747 10087 24781
rect 10035 24735 10087 24747
rect 10481 24883 10533 24909
rect 10481 24849 10491 24883
rect 10525 24849 10533 24883
rect 10481 24781 10533 24849
rect 10481 24747 10491 24781
rect 10525 24747 10533 24781
rect 10481 24735 10533 24747
rect 10587 24781 10639 24909
rect 10587 24747 10595 24781
rect 10629 24747 10639 24781
rect 10587 24735 10639 24747
rect 11585 24781 11637 24909
rect 11585 24747 11595 24781
rect 11629 24747 11637 24781
rect 11585 24735 11637 24747
rect 11691 24781 11743 24909
rect 11691 24747 11699 24781
rect 11733 24747 11743 24781
rect 11691 24735 11743 24747
rect 12689 24781 12741 24909
rect 12689 24747 12699 24781
rect 12733 24747 12741 24781
rect 12689 24735 12741 24747
rect 12795 24781 12847 24909
rect 12795 24747 12803 24781
rect 12837 24747 12847 24781
rect 12795 24735 12847 24747
rect 13793 24781 13845 24909
rect 13793 24747 13803 24781
rect 13837 24747 13845 24781
rect 13793 24735 13845 24747
rect 13899 24781 13951 24909
rect 13899 24747 13907 24781
rect 13941 24747 13951 24781
rect 13899 24735 13951 24747
rect 14897 24781 14949 24909
rect 14897 24747 14907 24781
rect 14941 24747 14949 24781
rect 15187 24883 15239 24909
rect 15187 24849 15195 24883
rect 15229 24849 15239 24883
rect 15187 24781 15239 24849
rect 14897 24735 14949 24747
rect 15187 24747 15195 24781
rect 15229 24747 15239 24781
rect 15187 24735 15239 24747
rect 15449 24883 15501 24909
rect 15449 24849 15459 24883
rect 15493 24849 15501 24883
rect 15449 24781 15501 24849
rect 15449 24747 15459 24781
rect 15493 24747 15501 24781
rect 15449 24735 15501 24747
rect 15555 24781 15607 24909
rect 15555 24747 15563 24781
rect 15597 24747 15607 24781
rect 15555 24735 15607 24747
rect 16553 24781 16605 24909
rect 16553 24747 16563 24781
rect 16597 24747 16605 24781
rect 16553 24735 16605 24747
rect 16659 24781 16711 24909
rect 16659 24747 16667 24781
rect 16701 24747 16711 24781
rect 16659 24735 16711 24747
rect 17657 24781 17709 24909
rect 17657 24747 17667 24781
rect 17701 24747 17709 24781
rect 17657 24735 17709 24747
rect 17763 24781 17815 24909
rect 17763 24747 17771 24781
rect 17805 24747 17815 24781
rect 17763 24735 17815 24747
rect 18761 24781 18813 24909
rect 18761 24747 18771 24781
rect 18805 24747 18813 24781
rect 18761 24735 18813 24747
rect 18867 24781 18919 24909
rect 18867 24747 18875 24781
rect 18909 24747 18919 24781
rect 18867 24735 18919 24747
rect 19865 24781 19917 24909
rect 19865 24747 19875 24781
rect 19909 24747 19917 24781
rect 19865 24735 19917 24747
rect 19971 24876 20023 24909
rect 19971 24842 19979 24876
rect 20013 24842 20023 24876
rect 19971 24781 20023 24842
rect 19971 24747 19979 24781
rect 20013 24747 20023 24781
rect 19971 24735 20023 24747
rect 20141 24876 20193 24909
rect 20141 24842 20151 24876
rect 20185 24842 20193 24876
rect 20141 24781 20193 24842
rect 20141 24747 20151 24781
rect 20185 24747 20193 24781
rect 20141 24735 20193 24747
rect 4975 24629 5027 24641
rect 4975 24595 4983 24629
rect 5017 24595 5027 24629
rect 4975 24534 5027 24595
rect 4975 24500 4983 24534
rect 5017 24500 5027 24534
rect 4975 24467 5027 24500
rect 5145 24629 5197 24641
rect 5145 24595 5155 24629
rect 5189 24595 5197 24629
rect 5145 24534 5197 24595
rect 5145 24500 5155 24534
rect 5189 24500 5197 24534
rect 5145 24467 5197 24500
rect 5435 24629 5487 24641
rect 5435 24595 5443 24629
rect 5477 24595 5487 24629
rect 5435 24527 5487 24595
rect 5435 24493 5443 24527
rect 5477 24493 5487 24527
rect 5435 24467 5487 24493
rect 6065 24629 6117 24641
rect 6065 24595 6075 24629
rect 6109 24595 6117 24629
rect 6065 24527 6117 24595
rect 6065 24493 6075 24527
rect 6109 24493 6117 24527
rect 6065 24467 6117 24493
rect 6171 24629 6223 24641
rect 6171 24595 6179 24629
rect 6213 24595 6223 24629
rect 6171 24467 6223 24595
rect 7169 24629 7221 24641
rect 7169 24595 7179 24629
rect 7213 24595 7221 24629
rect 7459 24629 7511 24641
rect 7169 24467 7221 24595
rect 7459 24595 7467 24629
rect 7501 24595 7511 24629
rect 7459 24527 7511 24595
rect 7459 24493 7467 24527
rect 7501 24493 7511 24527
rect 7459 24467 7511 24493
rect 7905 24629 7957 24641
rect 7905 24595 7915 24629
rect 7949 24595 7957 24629
rect 7905 24527 7957 24595
rect 7905 24493 7915 24527
rect 7949 24493 7957 24527
rect 7905 24467 7957 24493
rect 8011 24629 8063 24641
rect 8011 24595 8019 24629
rect 8053 24595 8063 24629
rect 8011 24467 8063 24595
rect 9009 24629 9061 24641
rect 9009 24595 9019 24629
rect 9053 24595 9061 24629
rect 9009 24467 9061 24595
rect 9115 24629 9167 24641
rect 9115 24595 9123 24629
rect 9157 24595 9167 24629
rect 9115 24467 9167 24595
rect 10113 24629 10165 24641
rect 10113 24595 10123 24629
rect 10157 24595 10165 24629
rect 10113 24467 10165 24595
rect 10219 24629 10271 24641
rect 10219 24595 10227 24629
rect 10261 24595 10271 24629
rect 10219 24467 10271 24595
rect 11217 24629 11269 24641
rect 11217 24595 11227 24629
rect 11261 24595 11269 24629
rect 11217 24467 11269 24595
rect 11323 24629 11375 24641
rect 11323 24595 11331 24629
rect 11365 24595 11375 24629
rect 11323 24467 11375 24595
rect 12321 24629 12373 24641
rect 12321 24595 12331 24629
rect 12365 24595 12373 24629
rect 12611 24629 12663 24641
rect 12321 24467 12373 24595
rect 12611 24595 12619 24629
rect 12653 24595 12663 24629
rect 12611 24527 12663 24595
rect 12611 24493 12619 24527
rect 12653 24493 12663 24527
rect 12611 24467 12663 24493
rect 13057 24629 13109 24641
rect 13057 24595 13067 24629
rect 13101 24595 13109 24629
rect 13057 24527 13109 24595
rect 13057 24493 13067 24527
rect 13101 24493 13109 24527
rect 13057 24467 13109 24493
rect 13163 24629 13215 24641
rect 13163 24595 13171 24629
rect 13205 24595 13215 24629
rect 13163 24467 13215 24595
rect 14161 24629 14213 24641
rect 14161 24595 14171 24629
rect 14205 24595 14213 24629
rect 14161 24467 14213 24595
rect 14267 24629 14319 24641
rect 14267 24595 14275 24629
rect 14309 24595 14319 24629
rect 14267 24467 14319 24595
rect 15265 24629 15317 24641
rect 15265 24595 15275 24629
rect 15309 24595 15317 24629
rect 15265 24467 15317 24595
rect 15371 24629 15423 24641
rect 15371 24595 15379 24629
rect 15413 24595 15423 24629
rect 15371 24467 15423 24595
rect 16369 24629 16421 24641
rect 16369 24595 16379 24629
rect 16413 24595 16421 24629
rect 16369 24467 16421 24595
rect 16475 24629 16527 24641
rect 16475 24595 16483 24629
rect 16517 24595 16527 24629
rect 16475 24467 16527 24595
rect 17473 24629 17525 24641
rect 17473 24595 17483 24629
rect 17517 24595 17525 24629
rect 17763 24629 17815 24641
rect 17473 24467 17525 24595
rect 17763 24595 17771 24629
rect 17805 24595 17815 24629
rect 17763 24467 17815 24595
rect 18761 24629 18813 24641
rect 18761 24595 18771 24629
rect 18805 24595 18813 24629
rect 18761 24467 18813 24595
rect 18867 24629 18919 24641
rect 18867 24595 18875 24629
rect 18909 24595 18919 24629
rect 18867 24467 18919 24595
rect 19865 24629 19917 24641
rect 19865 24595 19875 24629
rect 19909 24595 19917 24629
rect 19865 24467 19917 24595
rect 19971 24629 20023 24641
rect 19971 24595 19979 24629
rect 20013 24595 20023 24629
rect 19971 24534 20023 24595
rect 19971 24500 19979 24534
rect 20013 24500 20023 24534
rect 19971 24467 20023 24500
rect 20141 24629 20193 24641
rect 20141 24595 20151 24629
rect 20185 24595 20193 24629
rect 20141 24534 20193 24595
rect 20141 24500 20151 24534
rect 20185 24500 20193 24534
rect 20141 24467 20193 24500
rect 4975 23788 5027 23821
rect 4975 23754 4983 23788
rect 5017 23754 5027 23788
rect 4975 23693 5027 23754
rect 4975 23659 4983 23693
rect 5017 23659 5027 23693
rect 4975 23647 5027 23659
rect 5145 23788 5197 23821
rect 5145 23754 5155 23788
rect 5189 23754 5197 23788
rect 5145 23693 5197 23754
rect 5145 23659 5155 23693
rect 5189 23659 5197 23693
rect 5145 23647 5197 23659
rect 5435 23693 5487 23821
rect 5435 23659 5443 23693
rect 5477 23659 5487 23693
rect 5435 23647 5487 23659
rect 6433 23693 6485 23821
rect 6433 23659 6443 23693
rect 6477 23659 6485 23693
rect 6433 23647 6485 23659
rect 6539 23693 6591 23821
rect 6539 23659 6547 23693
rect 6581 23659 6591 23693
rect 6539 23647 6591 23659
rect 7537 23693 7589 23821
rect 7537 23659 7547 23693
rect 7581 23659 7589 23693
rect 7537 23647 7589 23659
rect 7643 23693 7695 23821
rect 7643 23659 7651 23693
rect 7685 23659 7695 23693
rect 7643 23647 7695 23659
rect 8641 23693 8693 23821
rect 8641 23659 8651 23693
rect 8685 23659 8693 23693
rect 8641 23647 8693 23659
rect 8747 23693 8799 23821
rect 8747 23659 8755 23693
rect 8789 23659 8799 23693
rect 8747 23647 8799 23659
rect 9745 23693 9797 23821
rect 9745 23659 9755 23693
rect 9789 23659 9797 23693
rect 10035 23795 10087 23821
rect 10035 23761 10043 23795
rect 10077 23761 10087 23795
rect 10035 23693 10087 23761
rect 9745 23647 9797 23659
rect 10035 23659 10043 23693
rect 10077 23659 10087 23693
rect 10035 23647 10087 23659
rect 10481 23795 10533 23821
rect 10481 23761 10491 23795
rect 10525 23761 10533 23795
rect 10481 23693 10533 23761
rect 10481 23659 10491 23693
rect 10525 23659 10533 23693
rect 10481 23647 10533 23659
rect 10587 23693 10639 23821
rect 10587 23659 10595 23693
rect 10629 23659 10639 23693
rect 10587 23647 10639 23659
rect 11585 23693 11637 23821
rect 11585 23659 11595 23693
rect 11629 23659 11637 23693
rect 11585 23647 11637 23659
rect 11691 23693 11743 23821
rect 11691 23659 11699 23693
rect 11733 23659 11743 23693
rect 11691 23647 11743 23659
rect 12689 23693 12741 23821
rect 12689 23659 12699 23693
rect 12733 23659 12741 23693
rect 12689 23647 12741 23659
rect 12795 23693 12847 23821
rect 12795 23659 12803 23693
rect 12837 23659 12847 23693
rect 12795 23647 12847 23659
rect 13793 23693 13845 23821
rect 13793 23659 13803 23693
rect 13837 23659 13845 23693
rect 13793 23647 13845 23659
rect 13899 23693 13951 23821
rect 13899 23659 13907 23693
rect 13941 23659 13951 23693
rect 13899 23647 13951 23659
rect 14897 23693 14949 23821
rect 14897 23659 14907 23693
rect 14941 23659 14949 23693
rect 15187 23795 15239 23821
rect 15187 23761 15195 23795
rect 15229 23761 15239 23795
rect 15187 23693 15239 23761
rect 14897 23647 14949 23659
rect 15187 23659 15195 23693
rect 15229 23659 15239 23693
rect 15187 23647 15239 23659
rect 15449 23795 15501 23821
rect 15449 23761 15459 23795
rect 15493 23761 15501 23795
rect 15449 23693 15501 23761
rect 15449 23659 15459 23693
rect 15493 23659 15501 23693
rect 15449 23647 15501 23659
rect 15555 23693 15607 23821
rect 15555 23659 15563 23693
rect 15597 23659 15607 23693
rect 15555 23647 15607 23659
rect 16553 23693 16605 23821
rect 16553 23659 16563 23693
rect 16597 23659 16605 23693
rect 16553 23647 16605 23659
rect 16659 23693 16711 23821
rect 16659 23659 16667 23693
rect 16701 23659 16711 23693
rect 16659 23647 16711 23659
rect 17657 23693 17709 23821
rect 17657 23659 17667 23693
rect 17701 23659 17709 23693
rect 17657 23647 17709 23659
rect 17763 23693 17815 23821
rect 17763 23659 17771 23693
rect 17805 23659 17815 23693
rect 17763 23647 17815 23659
rect 18761 23693 18813 23821
rect 18761 23659 18771 23693
rect 18805 23659 18813 23693
rect 18761 23647 18813 23659
rect 18867 23693 18919 23821
rect 18867 23659 18875 23693
rect 18909 23659 18919 23693
rect 18867 23647 18919 23659
rect 19865 23693 19917 23821
rect 19865 23659 19875 23693
rect 19909 23659 19917 23693
rect 19865 23647 19917 23659
rect 19971 23788 20023 23821
rect 19971 23754 19979 23788
rect 20013 23754 20023 23788
rect 19971 23693 20023 23754
rect 19971 23659 19979 23693
rect 20013 23659 20023 23693
rect 19971 23647 20023 23659
rect 20141 23788 20193 23821
rect 20141 23754 20151 23788
rect 20185 23754 20193 23788
rect 20141 23693 20193 23754
rect 20141 23659 20151 23693
rect 20185 23659 20193 23693
rect 20141 23647 20193 23659
rect 4975 23541 5027 23553
rect 4975 23507 4983 23541
rect 5017 23507 5027 23541
rect 4975 23446 5027 23507
rect 4975 23412 4983 23446
rect 5017 23412 5027 23446
rect 4975 23379 5027 23412
rect 5145 23541 5197 23553
rect 5145 23507 5155 23541
rect 5189 23507 5197 23541
rect 5145 23446 5197 23507
rect 5145 23412 5155 23446
rect 5189 23412 5197 23446
rect 5145 23379 5197 23412
rect 5435 23541 5487 23553
rect 5435 23507 5443 23541
rect 5477 23507 5487 23541
rect 5435 23439 5487 23507
rect 5435 23405 5443 23439
rect 5477 23405 5487 23439
rect 5435 23379 5487 23405
rect 6065 23541 6117 23553
rect 6065 23507 6075 23541
rect 6109 23507 6117 23541
rect 6065 23439 6117 23507
rect 6065 23405 6075 23439
rect 6109 23405 6117 23439
rect 6065 23379 6117 23405
rect 6171 23541 6223 23553
rect 6171 23507 6179 23541
rect 6213 23507 6223 23541
rect 6171 23379 6223 23507
rect 7169 23541 7221 23553
rect 7169 23507 7179 23541
rect 7213 23507 7221 23541
rect 7459 23541 7511 23553
rect 7169 23379 7221 23507
rect 7459 23507 7467 23541
rect 7501 23507 7511 23541
rect 7459 23439 7511 23507
rect 7459 23405 7467 23439
rect 7501 23405 7511 23439
rect 7459 23379 7511 23405
rect 7905 23541 7957 23553
rect 7905 23507 7915 23541
rect 7949 23507 7957 23541
rect 7905 23439 7957 23507
rect 7905 23405 7915 23439
rect 7949 23405 7957 23439
rect 7905 23379 7957 23405
rect 8011 23541 8063 23553
rect 8011 23507 8019 23541
rect 8053 23507 8063 23541
rect 8011 23379 8063 23507
rect 9009 23541 9061 23553
rect 9009 23507 9019 23541
rect 9053 23507 9061 23541
rect 9009 23379 9061 23507
rect 9115 23541 9167 23553
rect 9115 23507 9123 23541
rect 9157 23507 9167 23541
rect 9115 23379 9167 23507
rect 10113 23541 10165 23553
rect 10113 23507 10123 23541
rect 10157 23507 10165 23541
rect 10113 23379 10165 23507
rect 10219 23541 10271 23553
rect 10219 23507 10227 23541
rect 10261 23507 10271 23541
rect 10219 23379 10271 23507
rect 11217 23541 11269 23553
rect 11217 23507 11227 23541
rect 11261 23507 11269 23541
rect 11217 23379 11269 23507
rect 11323 23541 11375 23553
rect 11323 23507 11331 23541
rect 11365 23507 11375 23541
rect 11323 23379 11375 23507
rect 12321 23541 12373 23553
rect 12321 23507 12331 23541
rect 12365 23507 12373 23541
rect 12611 23541 12663 23553
rect 12321 23379 12373 23507
rect 12611 23507 12619 23541
rect 12653 23507 12663 23541
rect 12611 23439 12663 23507
rect 12611 23405 12619 23439
rect 12653 23405 12663 23439
rect 12611 23379 12663 23405
rect 13057 23541 13109 23553
rect 13057 23507 13067 23541
rect 13101 23507 13109 23541
rect 13057 23439 13109 23507
rect 13057 23405 13067 23439
rect 13101 23405 13109 23439
rect 13057 23379 13109 23405
rect 13163 23541 13215 23553
rect 13163 23507 13171 23541
rect 13205 23507 13215 23541
rect 13163 23379 13215 23507
rect 14161 23541 14213 23553
rect 14161 23507 14171 23541
rect 14205 23507 14213 23541
rect 14161 23379 14213 23507
rect 14267 23541 14319 23553
rect 14267 23507 14275 23541
rect 14309 23507 14319 23541
rect 14267 23379 14319 23507
rect 15265 23541 15317 23553
rect 15265 23507 15275 23541
rect 15309 23507 15317 23541
rect 15265 23379 15317 23507
rect 15371 23541 15423 23553
rect 15371 23507 15379 23541
rect 15413 23507 15423 23541
rect 15371 23379 15423 23507
rect 16369 23541 16421 23553
rect 16369 23507 16379 23541
rect 16413 23507 16421 23541
rect 16369 23379 16421 23507
rect 16475 23541 16527 23553
rect 16475 23507 16483 23541
rect 16517 23507 16527 23541
rect 16475 23379 16527 23507
rect 17473 23541 17525 23553
rect 17473 23507 17483 23541
rect 17517 23507 17525 23541
rect 17763 23541 17815 23553
rect 17473 23379 17525 23507
rect 17763 23507 17771 23541
rect 17805 23507 17815 23541
rect 17763 23379 17815 23507
rect 18761 23541 18813 23553
rect 18761 23507 18771 23541
rect 18805 23507 18813 23541
rect 18761 23379 18813 23507
rect 18867 23541 18919 23553
rect 18867 23507 18875 23541
rect 18909 23507 18919 23541
rect 18867 23379 18919 23507
rect 19865 23541 19917 23553
rect 19865 23507 19875 23541
rect 19909 23507 19917 23541
rect 19865 23379 19917 23507
rect 19971 23541 20023 23553
rect 19971 23507 19979 23541
rect 20013 23507 20023 23541
rect 19971 23446 20023 23507
rect 19971 23412 19979 23446
rect 20013 23412 20023 23446
rect 19971 23379 20023 23412
rect 20141 23541 20193 23553
rect 20141 23507 20151 23541
rect 20185 23507 20193 23541
rect 20141 23446 20193 23507
rect 20141 23412 20151 23446
rect 20185 23412 20193 23446
rect 20141 23379 20193 23412
rect 4975 22700 5027 22733
rect 4975 22666 4983 22700
rect 5017 22666 5027 22700
rect 4975 22605 5027 22666
rect 4975 22571 4983 22605
rect 5017 22571 5027 22605
rect 4975 22559 5027 22571
rect 5145 22700 5197 22733
rect 5145 22666 5155 22700
rect 5189 22666 5197 22700
rect 5145 22605 5197 22666
rect 5145 22571 5155 22605
rect 5189 22571 5197 22605
rect 5145 22559 5197 22571
rect 5435 22605 5487 22733
rect 5435 22571 5443 22605
rect 5477 22571 5487 22605
rect 5435 22559 5487 22571
rect 6433 22605 6485 22733
rect 6433 22571 6443 22605
rect 6477 22571 6485 22605
rect 6433 22559 6485 22571
rect 6539 22605 6591 22733
rect 6539 22571 6547 22605
rect 6581 22571 6591 22605
rect 6539 22559 6591 22571
rect 7537 22605 7589 22733
rect 7537 22571 7547 22605
rect 7581 22571 7589 22605
rect 7537 22559 7589 22571
rect 7643 22605 7695 22733
rect 7643 22571 7651 22605
rect 7685 22571 7695 22605
rect 7643 22559 7695 22571
rect 8641 22605 8693 22733
rect 8641 22571 8651 22605
rect 8685 22571 8693 22605
rect 8641 22559 8693 22571
rect 8747 22605 8799 22733
rect 8747 22571 8755 22605
rect 8789 22571 8799 22605
rect 8747 22559 8799 22571
rect 9745 22605 9797 22733
rect 9745 22571 9755 22605
rect 9789 22571 9797 22605
rect 10035 22707 10087 22733
rect 10035 22673 10043 22707
rect 10077 22673 10087 22707
rect 10035 22605 10087 22673
rect 9745 22559 9797 22571
rect 10035 22571 10043 22605
rect 10077 22571 10087 22605
rect 10035 22559 10087 22571
rect 10481 22707 10533 22733
rect 10481 22673 10491 22707
rect 10525 22673 10533 22707
rect 10481 22605 10533 22673
rect 10481 22571 10491 22605
rect 10525 22571 10533 22605
rect 10481 22559 10533 22571
rect 10587 22605 10639 22733
rect 10587 22571 10595 22605
rect 10629 22571 10639 22605
rect 10587 22559 10639 22571
rect 11585 22605 11637 22733
rect 11585 22571 11595 22605
rect 11629 22571 11637 22605
rect 11585 22559 11637 22571
rect 11691 22605 11743 22733
rect 11691 22571 11699 22605
rect 11733 22571 11743 22605
rect 11691 22559 11743 22571
rect 12689 22605 12741 22733
rect 12689 22571 12699 22605
rect 12733 22571 12741 22605
rect 12689 22559 12741 22571
rect 12795 22605 12847 22733
rect 12795 22571 12803 22605
rect 12837 22571 12847 22605
rect 12795 22559 12847 22571
rect 13793 22605 13845 22733
rect 13793 22571 13803 22605
rect 13837 22571 13845 22605
rect 13793 22559 13845 22571
rect 13899 22605 13951 22733
rect 13899 22571 13907 22605
rect 13941 22571 13951 22605
rect 13899 22559 13951 22571
rect 14897 22605 14949 22733
rect 14897 22571 14907 22605
rect 14941 22571 14949 22605
rect 15187 22707 15239 22733
rect 15187 22673 15195 22707
rect 15229 22673 15239 22707
rect 15187 22605 15239 22673
rect 14897 22559 14949 22571
rect 15187 22571 15195 22605
rect 15229 22571 15239 22605
rect 15187 22559 15239 22571
rect 15449 22707 15501 22733
rect 15449 22673 15459 22707
rect 15493 22673 15501 22707
rect 15449 22605 15501 22673
rect 15449 22571 15459 22605
rect 15493 22571 15501 22605
rect 15449 22559 15501 22571
rect 15555 22605 15607 22733
rect 15555 22571 15563 22605
rect 15597 22571 15607 22605
rect 15555 22559 15607 22571
rect 16553 22605 16605 22733
rect 16553 22571 16563 22605
rect 16597 22571 16605 22605
rect 16553 22559 16605 22571
rect 16659 22605 16711 22733
rect 16659 22571 16667 22605
rect 16701 22571 16711 22605
rect 16659 22559 16711 22571
rect 17657 22605 17709 22733
rect 17657 22571 17667 22605
rect 17701 22571 17709 22605
rect 17657 22559 17709 22571
rect 17763 22605 17815 22733
rect 17763 22571 17771 22605
rect 17805 22571 17815 22605
rect 17763 22559 17815 22571
rect 18761 22605 18813 22733
rect 18761 22571 18771 22605
rect 18805 22571 18813 22605
rect 18761 22559 18813 22571
rect 18867 22605 18919 22733
rect 18867 22571 18875 22605
rect 18909 22571 18919 22605
rect 18867 22559 18919 22571
rect 19865 22605 19917 22733
rect 19865 22571 19875 22605
rect 19909 22571 19917 22605
rect 19865 22559 19917 22571
rect 19971 22700 20023 22733
rect 19971 22666 19979 22700
rect 20013 22666 20023 22700
rect 19971 22605 20023 22666
rect 19971 22571 19979 22605
rect 20013 22571 20023 22605
rect 19971 22559 20023 22571
rect 20141 22700 20193 22733
rect 20141 22666 20151 22700
rect 20185 22666 20193 22700
rect 20141 22605 20193 22666
rect 20141 22571 20151 22605
rect 20185 22571 20193 22605
rect 20141 22559 20193 22571
rect 4975 22453 5027 22465
rect 4975 22419 4983 22453
rect 5017 22419 5027 22453
rect 4975 22358 5027 22419
rect 4975 22324 4983 22358
rect 5017 22324 5027 22358
rect 4975 22291 5027 22324
rect 5145 22453 5197 22465
rect 5145 22419 5155 22453
rect 5189 22419 5197 22453
rect 5145 22358 5197 22419
rect 5145 22324 5155 22358
rect 5189 22324 5197 22358
rect 5145 22291 5197 22324
rect 5435 22453 5487 22465
rect 5435 22419 5443 22453
rect 5477 22419 5487 22453
rect 5435 22351 5487 22419
rect 5435 22317 5443 22351
rect 5477 22317 5487 22351
rect 5435 22291 5487 22317
rect 6065 22453 6117 22465
rect 6065 22419 6075 22453
rect 6109 22419 6117 22453
rect 6065 22351 6117 22419
rect 6065 22317 6075 22351
rect 6109 22317 6117 22351
rect 6065 22291 6117 22317
rect 6171 22453 6223 22465
rect 6171 22419 6179 22453
rect 6213 22419 6223 22453
rect 6171 22291 6223 22419
rect 7169 22453 7221 22465
rect 7169 22419 7179 22453
rect 7213 22419 7221 22453
rect 7459 22453 7511 22465
rect 7169 22291 7221 22419
rect 7459 22419 7467 22453
rect 7501 22419 7511 22453
rect 7459 22351 7511 22419
rect 7459 22317 7467 22351
rect 7501 22317 7511 22351
rect 7459 22291 7511 22317
rect 7905 22453 7957 22465
rect 7905 22419 7915 22453
rect 7949 22419 7957 22453
rect 7905 22351 7957 22419
rect 7905 22317 7915 22351
rect 7949 22317 7957 22351
rect 7905 22291 7957 22317
rect 8011 22453 8063 22465
rect 8011 22419 8019 22453
rect 8053 22419 8063 22453
rect 8011 22291 8063 22419
rect 9009 22453 9061 22465
rect 9009 22419 9019 22453
rect 9053 22419 9061 22453
rect 9009 22291 9061 22419
rect 9115 22453 9167 22465
rect 9115 22419 9123 22453
rect 9157 22419 9167 22453
rect 9115 22291 9167 22419
rect 10113 22453 10165 22465
rect 10113 22419 10123 22453
rect 10157 22419 10165 22453
rect 10113 22291 10165 22419
rect 10219 22453 10271 22465
rect 10219 22419 10227 22453
rect 10261 22419 10271 22453
rect 10219 22291 10271 22419
rect 11217 22453 11269 22465
rect 11217 22419 11227 22453
rect 11261 22419 11269 22453
rect 11217 22291 11269 22419
rect 11323 22453 11375 22465
rect 11323 22419 11331 22453
rect 11365 22419 11375 22453
rect 11323 22291 11375 22419
rect 12321 22453 12373 22465
rect 12321 22419 12331 22453
rect 12365 22419 12373 22453
rect 12611 22453 12663 22465
rect 12321 22291 12373 22419
rect 12611 22419 12619 22453
rect 12653 22419 12663 22453
rect 12611 22351 12663 22419
rect 12611 22317 12619 22351
rect 12653 22317 12663 22351
rect 12611 22291 12663 22317
rect 13057 22453 13109 22465
rect 13057 22419 13067 22453
rect 13101 22419 13109 22453
rect 13057 22351 13109 22419
rect 13057 22317 13067 22351
rect 13101 22317 13109 22351
rect 13057 22291 13109 22317
rect 13163 22453 13215 22465
rect 13163 22419 13171 22453
rect 13205 22419 13215 22453
rect 13163 22291 13215 22419
rect 14161 22453 14213 22465
rect 14161 22419 14171 22453
rect 14205 22419 14213 22453
rect 14161 22291 14213 22419
rect 14267 22453 14319 22465
rect 14267 22419 14275 22453
rect 14309 22419 14319 22453
rect 14267 22291 14319 22419
rect 15265 22453 15317 22465
rect 15265 22419 15275 22453
rect 15309 22419 15317 22453
rect 15265 22291 15317 22419
rect 15371 22453 15423 22465
rect 15371 22419 15379 22453
rect 15413 22419 15423 22453
rect 15371 22291 15423 22419
rect 16369 22453 16421 22465
rect 16369 22419 16379 22453
rect 16413 22419 16421 22453
rect 16369 22291 16421 22419
rect 16475 22453 16527 22465
rect 16475 22419 16483 22453
rect 16517 22419 16527 22453
rect 16475 22291 16527 22419
rect 17473 22453 17525 22465
rect 17473 22419 17483 22453
rect 17517 22419 17525 22453
rect 17763 22453 17815 22465
rect 17473 22291 17525 22419
rect 17763 22419 17771 22453
rect 17805 22419 17815 22453
rect 17763 22291 17815 22419
rect 18761 22453 18813 22465
rect 18761 22419 18771 22453
rect 18805 22419 18813 22453
rect 18761 22291 18813 22419
rect 18867 22453 18919 22465
rect 18867 22419 18875 22453
rect 18909 22419 18919 22453
rect 18867 22291 18919 22419
rect 19865 22453 19917 22465
rect 19865 22419 19875 22453
rect 19909 22419 19917 22453
rect 19865 22291 19917 22419
rect 19971 22453 20023 22465
rect 19971 22419 19979 22453
rect 20013 22419 20023 22453
rect 19971 22358 20023 22419
rect 19971 22324 19979 22358
rect 20013 22324 20023 22358
rect 19971 22291 20023 22324
rect 20141 22453 20193 22465
rect 20141 22419 20151 22453
rect 20185 22419 20193 22453
rect 20141 22358 20193 22419
rect 20141 22324 20151 22358
rect 20185 22324 20193 22358
rect 20141 22291 20193 22324
rect 4975 21612 5027 21645
rect 4975 21578 4983 21612
rect 5017 21578 5027 21612
rect 4975 21517 5027 21578
rect 4975 21483 4983 21517
rect 5017 21483 5027 21517
rect 4975 21471 5027 21483
rect 5145 21612 5197 21645
rect 5145 21578 5155 21612
rect 5189 21578 5197 21612
rect 5145 21517 5197 21578
rect 5145 21483 5155 21517
rect 5189 21483 5197 21517
rect 5145 21471 5197 21483
rect 5435 21517 5487 21645
rect 5435 21483 5443 21517
rect 5477 21483 5487 21517
rect 5435 21471 5487 21483
rect 6433 21517 6485 21645
rect 6433 21483 6443 21517
rect 6477 21483 6485 21517
rect 6433 21471 6485 21483
rect 6539 21517 6591 21645
rect 6539 21483 6547 21517
rect 6581 21483 6591 21517
rect 6539 21471 6591 21483
rect 7537 21517 7589 21645
rect 7537 21483 7547 21517
rect 7581 21483 7589 21517
rect 7537 21471 7589 21483
rect 7643 21517 7695 21645
rect 7643 21483 7651 21517
rect 7685 21483 7695 21517
rect 7643 21471 7695 21483
rect 8641 21517 8693 21645
rect 8641 21483 8651 21517
rect 8685 21483 8693 21517
rect 8641 21471 8693 21483
rect 8747 21517 8799 21645
rect 8747 21483 8755 21517
rect 8789 21483 8799 21517
rect 8747 21471 8799 21483
rect 9745 21517 9797 21645
rect 9745 21483 9755 21517
rect 9789 21483 9797 21517
rect 10035 21619 10087 21645
rect 10035 21585 10043 21619
rect 10077 21585 10087 21619
rect 10035 21517 10087 21585
rect 9745 21471 9797 21483
rect 10035 21483 10043 21517
rect 10077 21483 10087 21517
rect 10035 21471 10087 21483
rect 10481 21619 10533 21645
rect 10481 21585 10491 21619
rect 10525 21585 10533 21619
rect 10481 21517 10533 21585
rect 10481 21483 10491 21517
rect 10525 21483 10533 21517
rect 10481 21471 10533 21483
rect 10587 21517 10639 21645
rect 10587 21483 10595 21517
rect 10629 21483 10639 21517
rect 10587 21471 10639 21483
rect 11585 21517 11637 21645
rect 11585 21483 11595 21517
rect 11629 21483 11637 21517
rect 11585 21471 11637 21483
rect 11691 21517 11743 21645
rect 11691 21483 11699 21517
rect 11733 21483 11743 21517
rect 11691 21471 11743 21483
rect 12689 21517 12741 21645
rect 12689 21483 12699 21517
rect 12733 21483 12741 21517
rect 12689 21471 12741 21483
rect 12795 21517 12847 21645
rect 12795 21483 12803 21517
rect 12837 21483 12847 21517
rect 12795 21471 12847 21483
rect 13793 21517 13845 21645
rect 13793 21483 13803 21517
rect 13837 21483 13845 21517
rect 13793 21471 13845 21483
rect 13899 21517 13951 21645
rect 13899 21483 13907 21517
rect 13941 21483 13951 21517
rect 13899 21471 13951 21483
rect 14897 21517 14949 21645
rect 14897 21483 14907 21517
rect 14941 21483 14949 21517
rect 15187 21619 15239 21645
rect 15187 21585 15195 21619
rect 15229 21585 15239 21619
rect 15187 21517 15239 21585
rect 14897 21471 14949 21483
rect 15187 21483 15195 21517
rect 15229 21483 15239 21517
rect 15187 21471 15239 21483
rect 15449 21619 15501 21645
rect 15449 21585 15459 21619
rect 15493 21585 15501 21619
rect 15449 21517 15501 21585
rect 15449 21483 15459 21517
rect 15493 21483 15501 21517
rect 15449 21471 15501 21483
rect 15555 21517 15607 21645
rect 15555 21483 15563 21517
rect 15597 21483 15607 21517
rect 15555 21471 15607 21483
rect 16553 21517 16605 21645
rect 16553 21483 16563 21517
rect 16597 21483 16605 21517
rect 16553 21471 16605 21483
rect 16659 21517 16711 21645
rect 16659 21483 16667 21517
rect 16701 21483 16711 21517
rect 16659 21471 16711 21483
rect 17657 21517 17709 21645
rect 17657 21483 17667 21517
rect 17701 21483 17709 21517
rect 17657 21471 17709 21483
rect 17763 21517 17815 21645
rect 17763 21483 17771 21517
rect 17805 21483 17815 21517
rect 17763 21471 17815 21483
rect 18761 21517 18813 21645
rect 18761 21483 18771 21517
rect 18805 21483 18813 21517
rect 18761 21471 18813 21483
rect 18867 21517 18919 21645
rect 18867 21483 18875 21517
rect 18909 21483 18919 21517
rect 18867 21471 18919 21483
rect 19865 21517 19917 21645
rect 19865 21483 19875 21517
rect 19909 21483 19917 21517
rect 19865 21471 19917 21483
rect 19971 21612 20023 21645
rect 19971 21578 19979 21612
rect 20013 21578 20023 21612
rect 19971 21517 20023 21578
rect 19971 21483 19979 21517
rect 20013 21483 20023 21517
rect 19971 21471 20023 21483
rect 20141 21612 20193 21645
rect 20141 21578 20151 21612
rect 20185 21578 20193 21612
rect 20141 21517 20193 21578
rect 20141 21483 20151 21517
rect 20185 21483 20193 21517
rect 20141 21471 20193 21483
rect 4975 21365 5027 21377
rect 4975 21331 4983 21365
rect 5017 21331 5027 21365
rect 4975 21270 5027 21331
rect 4975 21236 4983 21270
rect 5017 21236 5027 21270
rect 4975 21203 5027 21236
rect 5145 21365 5197 21377
rect 5145 21331 5155 21365
rect 5189 21331 5197 21365
rect 5145 21270 5197 21331
rect 5145 21236 5155 21270
rect 5189 21236 5197 21270
rect 5145 21203 5197 21236
rect 5435 21365 5487 21377
rect 5435 21331 5443 21365
rect 5477 21331 5487 21365
rect 5435 21263 5487 21331
rect 5435 21229 5443 21263
rect 5477 21229 5487 21263
rect 5435 21203 5487 21229
rect 6065 21365 6117 21377
rect 6065 21331 6075 21365
rect 6109 21331 6117 21365
rect 6065 21263 6117 21331
rect 6065 21229 6075 21263
rect 6109 21229 6117 21263
rect 6065 21203 6117 21229
rect 6171 21365 6223 21377
rect 6171 21331 6179 21365
rect 6213 21331 6223 21365
rect 6171 21203 6223 21331
rect 7169 21365 7221 21377
rect 7169 21331 7179 21365
rect 7213 21331 7221 21365
rect 7459 21365 7511 21377
rect 7169 21203 7221 21331
rect 7459 21331 7467 21365
rect 7501 21331 7511 21365
rect 7459 21263 7511 21331
rect 7459 21229 7467 21263
rect 7501 21229 7511 21263
rect 7459 21203 7511 21229
rect 7905 21365 7957 21377
rect 7905 21331 7915 21365
rect 7949 21331 7957 21365
rect 7905 21263 7957 21331
rect 7905 21229 7915 21263
rect 7949 21229 7957 21263
rect 7905 21203 7957 21229
rect 8011 21365 8063 21377
rect 8011 21331 8019 21365
rect 8053 21331 8063 21365
rect 8011 21203 8063 21331
rect 9009 21365 9061 21377
rect 9009 21331 9019 21365
rect 9053 21331 9061 21365
rect 9009 21203 9061 21331
rect 9115 21365 9167 21377
rect 9115 21331 9123 21365
rect 9157 21331 9167 21365
rect 9115 21203 9167 21331
rect 10113 21365 10165 21377
rect 10113 21331 10123 21365
rect 10157 21331 10165 21365
rect 10113 21203 10165 21331
rect 10219 21365 10271 21377
rect 10219 21331 10227 21365
rect 10261 21331 10271 21365
rect 10219 21203 10271 21331
rect 11217 21365 11269 21377
rect 11217 21331 11227 21365
rect 11261 21331 11269 21365
rect 11217 21203 11269 21331
rect 11323 21365 11375 21377
rect 11323 21331 11331 21365
rect 11365 21331 11375 21365
rect 11323 21203 11375 21331
rect 12321 21365 12373 21377
rect 12321 21331 12331 21365
rect 12365 21331 12373 21365
rect 12611 21365 12663 21377
rect 12321 21203 12373 21331
rect 12611 21331 12619 21365
rect 12653 21331 12663 21365
rect 12611 21263 12663 21331
rect 12611 21229 12619 21263
rect 12653 21229 12663 21263
rect 12611 21203 12663 21229
rect 13057 21365 13109 21377
rect 13057 21331 13067 21365
rect 13101 21331 13109 21365
rect 13057 21263 13109 21331
rect 13057 21229 13067 21263
rect 13101 21229 13109 21263
rect 13057 21203 13109 21229
rect 13163 21365 13215 21377
rect 13163 21331 13171 21365
rect 13205 21331 13215 21365
rect 13163 21203 13215 21331
rect 14161 21365 14213 21377
rect 14161 21331 14171 21365
rect 14205 21331 14213 21365
rect 14161 21203 14213 21331
rect 14267 21365 14319 21377
rect 14267 21331 14275 21365
rect 14309 21331 14319 21365
rect 14267 21203 14319 21331
rect 15265 21365 15317 21377
rect 15265 21331 15275 21365
rect 15309 21331 15317 21365
rect 15265 21203 15317 21331
rect 15371 21365 15423 21377
rect 15371 21331 15379 21365
rect 15413 21331 15423 21365
rect 15371 21203 15423 21331
rect 16369 21365 16421 21377
rect 16369 21331 16379 21365
rect 16413 21331 16421 21365
rect 16369 21203 16421 21331
rect 16475 21365 16527 21377
rect 16475 21331 16483 21365
rect 16517 21331 16527 21365
rect 16475 21203 16527 21331
rect 17473 21365 17525 21377
rect 17473 21331 17483 21365
rect 17517 21331 17525 21365
rect 17763 21365 17815 21377
rect 17473 21203 17525 21331
rect 17763 21331 17771 21365
rect 17805 21331 17815 21365
rect 17763 21203 17815 21331
rect 18761 21365 18813 21377
rect 18761 21331 18771 21365
rect 18805 21331 18813 21365
rect 18761 21203 18813 21331
rect 18867 21365 18919 21377
rect 18867 21331 18875 21365
rect 18909 21331 18919 21365
rect 18867 21203 18919 21331
rect 19865 21365 19917 21377
rect 19865 21331 19875 21365
rect 19909 21331 19917 21365
rect 19865 21203 19917 21331
rect 19971 21365 20023 21377
rect 19971 21331 19979 21365
rect 20013 21331 20023 21365
rect 19971 21270 20023 21331
rect 19971 21236 19979 21270
rect 20013 21236 20023 21270
rect 19971 21203 20023 21236
rect 20141 21365 20193 21377
rect 20141 21331 20151 21365
rect 20185 21331 20193 21365
rect 20141 21270 20193 21331
rect 20141 21236 20151 21270
rect 20185 21236 20193 21270
rect 20141 21203 20193 21236
rect 4975 20524 5027 20557
rect 4975 20490 4983 20524
rect 5017 20490 5027 20524
rect 4975 20429 5027 20490
rect 4975 20395 4983 20429
rect 5017 20395 5027 20429
rect 4975 20383 5027 20395
rect 5145 20524 5197 20557
rect 5145 20490 5155 20524
rect 5189 20490 5197 20524
rect 5145 20429 5197 20490
rect 5145 20395 5155 20429
rect 5189 20395 5197 20429
rect 5145 20383 5197 20395
rect 5435 20429 5487 20557
rect 5435 20395 5443 20429
rect 5477 20395 5487 20429
rect 5435 20383 5487 20395
rect 6433 20429 6485 20557
rect 6433 20395 6443 20429
rect 6477 20395 6485 20429
rect 6433 20383 6485 20395
rect 6539 20429 6591 20557
rect 6539 20395 6547 20429
rect 6581 20395 6591 20429
rect 6539 20383 6591 20395
rect 7537 20429 7589 20557
rect 7537 20395 7547 20429
rect 7581 20395 7589 20429
rect 7537 20383 7589 20395
rect 7643 20429 7695 20557
rect 7643 20395 7651 20429
rect 7685 20395 7695 20429
rect 7643 20383 7695 20395
rect 8641 20429 8693 20557
rect 8641 20395 8651 20429
rect 8685 20395 8693 20429
rect 8641 20383 8693 20395
rect 8747 20429 8799 20557
rect 8747 20395 8755 20429
rect 8789 20395 8799 20429
rect 8747 20383 8799 20395
rect 9745 20429 9797 20557
rect 9745 20395 9755 20429
rect 9789 20395 9797 20429
rect 10035 20531 10087 20557
rect 10035 20497 10043 20531
rect 10077 20497 10087 20531
rect 10035 20429 10087 20497
rect 9745 20383 9797 20395
rect 10035 20395 10043 20429
rect 10077 20395 10087 20429
rect 10035 20383 10087 20395
rect 10481 20531 10533 20557
rect 10481 20497 10491 20531
rect 10525 20497 10533 20531
rect 10481 20429 10533 20497
rect 10481 20395 10491 20429
rect 10525 20395 10533 20429
rect 10481 20383 10533 20395
rect 10587 20429 10639 20557
rect 10587 20395 10595 20429
rect 10629 20395 10639 20429
rect 10587 20383 10639 20395
rect 11585 20429 11637 20557
rect 11585 20395 11595 20429
rect 11629 20395 11637 20429
rect 11585 20383 11637 20395
rect 11691 20429 11743 20557
rect 11691 20395 11699 20429
rect 11733 20395 11743 20429
rect 11691 20383 11743 20395
rect 12689 20429 12741 20557
rect 12689 20395 12699 20429
rect 12733 20395 12741 20429
rect 12689 20383 12741 20395
rect 12795 20429 12847 20557
rect 12795 20395 12803 20429
rect 12837 20395 12847 20429
rect 12795 20383 12847 20395
rect 13793 20429 13845 20557
rect 13793 20395 13803 20429
rect 13837 20395 13845 20429
rect 13793 20383 13845 20395
rect 13899 20429 13951 20557
rect 13899 20395 13907 20429
rect 13941 20395 13951 20429
rect 13899 20383 13951 20395
rect 14897 20429 14949 20557
rect 14897 20395 14907 20429
rect 14941 20395 14949 20429
rect 15187 20531 15239 20557
rect 15187 20497 15195 20531
rect 15229 20497 15239 20531
rect 15187 20429 15239 20497
rect 14897 20383 14949 20395
rect 15187 20395 15195 20429
rect 15229 20395 15239 20429
rect 15187 20383 15239 20395
rect 15449 20531 15501 20557
rect 15449 20497 15459 20531
rect 15493 20497 15501 20531
rect 15449 20429 15501 20497
rect 15449 20395 15459 20429
rect 15493 20395 15501 20429
rect 15449 20383 15501 20395
rect 15555 20429 15607 20557
rect 15555 20395 15563 20429
rect 15597 20395 15607 20429
rect 15555 20383 15607 20395
rect 16553 20429 16605 20557
rect 16553 20395 16563 20429
rect 16597 20395 16605 20429
rect 16553 20383 16605 20395
rect 16659 20429 16711 20557
rect 16659 20395 16667 20429
rect 16701 20395 16711 20429
rect 16659 20383 16711 20395
rect 17657 20429 17709 20557
rect 17657 20395 17667 20429
rect 17701 20395 17709 20429
rect 17657 20383 17709 20395
rect 17763 20429 17815 20557
rect 17763 20395 17771 20429
rect 17805 20395 17815 20429
rect 17763 20383 17815 20395
rect 18761 20429 18813 20557
rect 18761 20395 18771 20429
rect 18805 20395 18813 20429
rect 18761 20383 18813 20395
rect 18867 20429 18919 20557
rect 18867 20395 18875 20429
rect 18909 20395 18919 20429
rect 18867 20383 18919 20395
rect 19865 20429 19917 20557
rect 19865 20395 19875 20429
rect 19909 20395 19917 20429
rect 19865 20383 19917 20395
rect 19971 20524 20023 20557
rect 19971 20490 19979 20524
rect 20013 20490 20023 20524
rect 19971 20429 20023 20490
rect 19971 20395 19979 20429
rect 20013 20395 20023 20429
rect 19971 20383 20023 20395
rect 20141 20524 20193 20557
rect 20141 20490 20151 20524
rect 20185 20490 20193 20524
rect 20141 20429 20193 20490
rect 20141 20395 20151 20429
rect 20185 20395 20193 20429
rect 20141 20383 20193 20395
rect 4975 20277 5027 20289
rect 4975 20243 4983 20277
rect 5017 20243 5027 20277
rect 4975 20182 5027 20243
rect 4975 20148 4983 20182
rect 5017 20148 5027 20182
rect 4975 20115 5027 20148
rect 5145 20277 5197 20289
rect 5145 20243 5155 20277
rect 5189 20243 5197 20277
rect 5145 20182 5197 20243
rect 5145 20148 5155 20182
rect 5189 20148 5197 20182
rect 5145 20115 5197 20148
rect 5435 20277 5487 20289
rect 5435 20243 5443 20277
rect 5477 20243 5487 20277
rect 5435 20175 5487 20243
rect 5435 20141 5443 20175
rect 5477 20141 5487 20175
rect 5435 20115 5487 20141
rect 6065 20277 6117 20289
rect 6065 20243 6075 20277
rect 6109 20243 6117 20277
rect 6065 20175 6117 20243
rect 6065 20141 6075 20175
rect 6109 20141 6117 20175
rect 6065 20115 6117 20141
rect 6171 20277 6223 20289
rect 6171 20243 6179 20277
rect 6213 20243 6223 20277
rect 6171 20115 6223 20243
rect 7169 20277 7221 20289
rect 7169 20243 7179 20277
rect 7213 20243 7221 20277
rect 7459 20277 7511 20289
rect 7169 20115 7221 20243
rect 7459 20243 7467 20277
rect 7501 20243 7511 20277
rect 7459 20175 7511 20243
rect 7459 20141 7467 20175
rect 7501 20141 7511 20175
rect 7459 20115 7511 20141
rect 7905 20277 7957 20289
rect 7905 20243 7915 20277
rect 7949 20243 7957 20277
rect 7905 20175 7957 20243
rect 7905 20141 7915 20175
rect 7949 20141 7957 20175
rect 7905 20115 7957 20141
rect 8011 20277 8063 20289
rect 8011 20243 8019 20277
rect 8053 20243 8063 20277
rect 8011 20115 8063 20243
rect 9009 20277 9061 20289
rect 9009 20243 9019 20277
rect 9053 20243 9061 20277
rect 9009 20115 9061 20243
rect 9115 20277 9167 20289
rect 9115 20243 9123 20277
rect 9157 20243 9167 20277
rect 9115 20115 9167 20243
rect 10113 20277 10165 20289
rect 10113 20243 10123 20277
rect 10157 20243 10165 20277
rect 10113 20115 10165 20243
rect 10219 20277 10271 20289
rect 10219 20243 10227 20277
rect 10261 20243 10271 20277
rect 10219 20115 10271 20243
rect 11217 20277 11269 20289
rect 11217 20243 11227 20277
rect 11261 20243 11269 20277
rect 11217 20115 11269 20243
rect 11323 20277 11375 20289
rect 11323 20243 11331 20277
rect 11365 20243 11375 20277
rect 11323 20115 11375 20243
rect 12321 20277 12373 20289
rect 12321 20243 12331 20277
rect 12365 20243 12373 20277
rect 12611 20277 12663 20289
rect 12321 20115 12373 20243
rect 12611 20243 12619 20277
rect 12653 20243 12663 20277
rect 12611 20175 12663 20243
rect 12611 20141 12619 20175
rect 12653 20141 12663 20175
rect 12611 20115 12663 20141
rect 13057 20277 13109 20289
rect 13057 20243 13067 20277
rect 13101 20243 13109 20277
rect 13057 20175 13109 20243
rect 13057 20141 13067 20175
rect 13101 20141 13109 20175
rect 13057 20115 13109 20141
rect 13163 20277 13215 20289
rect 13163 20243 13171 20277
rect 13205 20243 13215 20277
rect 13163 20115 13215 20243
rect 14161 20277 14213 20289
rect 14161 20243 14171 20277
rect 14205 20243 14213 20277
rect 14161 20115 14213 20243
rect 14267 20277 14319 20289
rect 14267 20243 14275 20277
rect 14309 20243 14319 20277
rect 14267 20115 14319 20243
rect 15265 20277 15317 20289
rect 15265 20243 15275 20277
rect 15309 20243 15317 20277
rect 15265 20115 15317 20243
rect 15371 20277 15423 20289
rect 15371 20243 15379 20277
rect 15413 20243 15423 20277
rect 15371 20115 15423 20243
rect 16369 20277 16421 20289
rect 16369 20243 16379 20277
rect 16413 20243 16421 20277
rect 16369 20115 16421 20243
rect 16475 20277 16527 20289
rect 16475 20243 16483 20277
rect 16517 20243 16527 20277
rect 16475 20115 16527 20243
rect 17473 20277 17525 20289
rect 17473 20243 17483 20277
rect 17517 20243 17525 20277
rect 17763 20277 17815 20289
rect 17473 20115 17525 20243
rect 17763 20243 17771 20277
rect 17805 20243 17815 20277
rect 17763 20115 17815 20243
rect 18761 20277 18813 20289
rect 18761 20243 18771 20277
rect 18805 20243 18813 20277
rect 18761 20115 18813 20243
rect 18867 20277 18919 20289
rect 18867 20243 18875 20277
rect 18909 20243 18919 20277
rect 18867 20115 18919 20243
rect 19865 20277 19917 20289
rect 19865 20243 19875 20277
rect 19909 20243 19917 20277
rect 19865 20115 19917 20243
rect 19971 20277 20023 20289
rect 19971 20243 19979 20277
rect 20013 20243 20023 20277
rect 19971 20182 20023 20243
rect 19971 20148 19979 20182
rect 20013 20148 20023 20182
rect 19971 20115 20023 20148
rect 20141 20277 20193 20289
rect 20141 20243 20151 20277
rect 20185 20243 20193 20277
rect 20141 20182 20193 20243
rect 20141 20148 20151 20182
rect 20185 20148 20193 20182
rect 20141 20115 20193 20148
rect 4975 19436 5027 19469
rect 4975 19402 4983 19436
rect 5017 19402 5027 19436
rect 4975 19341 5027 19402
rect 4975 19307 4983 19341
rect 5017 19307 5027 19341
rect 4975 19295 5027 19307
rect 5145 19436 5197 19469
rect 5145 19402 5155 19436
rect 5189 19402 5197 19436
rect 5145 19341 5197 19402
rect 5145 19307 5155 19341
rect 5189 19307 5197 19341
rect 5145 19295 5197 19307
rect 5435 19341 5487 19469
rect 5435 19307 5443 19341
rect 5477 19307 5487 19341
rect 5435 19295 5487 19307
rect 6433 19341 6485 19469
rect 6433 19307 6443 19341
rect 6477 19307 6485 19341
rect 6433 19295 6485 19307
rect 6539 19341 6591 19469
rect 6539 19307 6547 19341
rect 6581 19307 6591 19341
rect 6539 19295 6591 19307
rect 7537 19341 7589 19469
rect 7537 19307 7547 19341
rect 7581 19307 7589 19341
rect 7537 19295 7589 19307
rect 7643 19341 7695 19469
rect 7643 19307 7651 19341
rect 7685 19307 7695 19341
rect 7643 19295 7695 19307
rect 8641 19341 8693 19469
rect 8641 19307 8651 19341
rect 8685 19307 8693 19341
rect 8641 19295 8693 19307
rect 8747 19341 8799 19469
rect 8747 19307 8755 19341
rect 8789 19307 8799 19341
rect 8747 19295 8799 19307
rect 9745 19341 9797 19469
rect 9745 19307 9755 19341
rect 9789 19307 9797 19341
rect 10035 19443 10087 19469
rect 10035 19409 10043 19443
rect 10077 19409 10087 19443
rect 10035 19341 10087 19409
rect 9745 19295 9797 19307
rect 10035 19307 10043 19341
rect 10077 19307 10087 19341
rect 10035 19295 10087 19307
rect 10481 19443 10533 19469
rect 10481 19409 10491 19443
rect 10525 19409 10533 19443
rect 10481 19341 10533 19409
rect 10481 19307 10491 19341
rect 10525 19307 10533 19341
rect 10481 19295 10533 19307
rect 10587 19341 10639 19469
rect 10587 19307 10595 19341
rect 10629 19307 10639 19341
rect 10587 19295 10639 19307
rect 11585 19341 11637 19469
rect 11585 19307 11595 19341
rect 11629 19307 11637 19341
rect 11585 19295 11637 19307
rect 11691 19341 11743 19469
rect 11691 19307 11699 19341
rect 11733 19307 11743 19341
rect 11691 19295 11743 19307
rect 12689 19341 12741 19469
rect 12689 19307 12699 19341
rect 12733 19307 12741 19341
rect 12689 19295 12741 19307
rect 12795 19341 12847 19469
rect 12795 19307 12803 19341
rect 12837 19307 12847 19341
rect 12795 19295 12847 19307
rect 13793 19341 13845 19469
rect 13793 19307 13803 19341
rect 13837 19307 13845 19341
rect 13793 19295 13845 19307
rect 13899 19341 13951 19469
rect 13899 19307 13907 19341
rect 13941 19307 13951 19341
rect 13899 19295 13951 19307
rect 14897 19341 14949 19469
rect 14897 19307 14907 19341
rect 14941 19307 14949 19341
rect 15187 19443 15239 19469
rect 15187 19409 15195 19443
rect 15229 19409 15239 19443
rect 15187 19341 15239 19409
rect 14897 19295 14949 19307
rect 15187 19307 15195 19341
rect 15229 19307 15239 19341
rect 15187 19295 15239 19307
rect 15449 19443 15501 19469
rect 15449 19409 15459 19443
rect 15493 19409 15501 19443
rect 15449 19341 15501 19409
rect 15449 19307 15459 19341
rect 15493 19307 15501 19341
rect 15449 19295 15501 19307
rect 15555 19341 15607 19469
rect 15555 19307 15563 19341
rect 15597 19307 15607 19341
rect 15555 19295 15607 19307
rect 16553 19341 16605 19469
rect 16553 19307 16563 19341
rect 16597 19307 16605 19341
rect 16553 19295 16605 19307
rect 16659 19341 16711 19469
rect 16659 19307 16667 19341
rect 16701 19307 16711 19341
rect 16659 19295 16711 19307
rect 17657 19341 17709 19469
rect 17657 19307 17667 19341
rect 17701 19307 17709 19341
rect 17657 19295 17709 19307
rect 17763 19341 17815 19469
rect 17763 19307 17771 19341
rect 17805 19307 17815 19341
rect 17763 19295 17815 19307
rect 18761 19341 18813 19469
rect 18761 19307 18771 19341
rect 18805 19307 18813 19341
rect 18761 19295 18813 19307
rect 18867 19341 18919 19469
rect 18867 19307 18875 19341
rect 18909 19307 18919 19341
rect 18867 19295 18919 19307
rect 19865 19341 19917 19469
rect 19865 19307 19875 19341
rect 19909 19307 19917 19341
rect 19865 19295 19917 19307
rect 19971 19436 20023 19469
rect 19971 19402 19979 19436
rect 20013 19402 20023 19436
rect 19971 19341 20023 19402
rect 19971 19307 19979 19341
rect 20013 19307 20023 19341
rect 19971 19295 20023 19307
rect 20141 19436 20193 19469
rect 20141 19402 20151 19436
rect 20185 19402 20193 19436
rect 20141 19341 20193 19402
rect 20141 19307 20151 19341
rect 20185 19307 20193 19341
rect 20141 19295 20193 19307
rect 4975 19189 5027 19201
rect 4975 19155 4983 19189
rect 5017 19155 5027 19189
rect 4975 19094 5027 19155
rect 4975 19060 4983 19094
rect 5017 19060 5027 19094
rect 4975 19027 5027 19060
rect 5145 19189 5197 19201
rect 5145 19155 5155 19189
rect 5189 19155 5197 19189
rect 5145 19094 5197 19155
rect 5145 19060 5155 19094
rect 5189 19060 5197 19094
rect 5145 19027 5197 19060
rect 5435 19189 5487 19201
rect 5435 19155 5443 19189
rect 5477 19155 5487 19189
rect 5435 19087 5487 19155
rect 5435 19053 5443 19087
rect 5477 19053 5487 19087
rect 5435 19027 5487 19053
rect 6065 19189 6117 19201
rect 6065 19155 6075 19189
rect 6109 19155 6117 19189
rect 6065 19087 6117 19155
rect 6065 19053 6075 19087
rect 6109 19053 6117 19087
rect 6065 19027 6117 19053
rect 6171 19189 6223 19201
rect 6171 19155 6179 19189
rect 6213 19155 6223 19189
rect 6171 19027 6223 19155
rect 7169 19189 7221 19201
rect 7169 19155 7179 19189
rect 7213 19155 7221 19189
rect 7459 19189 7511 19201
rect 7169 19027 7221 19155
rect 7459 19155 7467 19189
rect 7501 19155 7511 19189
rect 7459 19087 7511 19155
rect 7459 19053 7467 19087
rect 7501 19053 7511 19087
rect 7459 19027 7511 19053
rect 7905 19189 7957 19201
rect 7905 19155 7915 19189
rect 7949 19155 7957 19189
rect 7905 19087 7957 19155
rect 7905 19053 7915 19087
rect 7949 19053 7957 19087
rect 7905 19027 7957 19053
rect 8011 19189 8063 19201
rect 8011 19155 8019 19189
rect 8053 19155 8063 19189
rect 8011 19027 8063 19155
rect 9009 19189 9061 19201
rect 9009 19155 9019 19189
rect 9053 19155 9061 19189
rect 9009 19027 9061 19155
rect 9115 19189 9167 19201
rect 9115 19155 9123 19189
rect 9157 19155 9167 19189
rect 9115 19027 9167 19155
rect 10113 19189 10165 19201
rect 10113 19155 10123 19189
rect 10157 19155 10165 19189
rect 10113 19027 10165 19155
rect 10219 19189 10271 19201
rect 10219 19155 10227 19189
rect 10261 19155 10271 19189
rect 10219 19027 10271 19155
rect 11217 19189 11269 19201
rect 11217 19155 11227 19189
rect 11261 19155 11269 19189
rect 11217 19027 11269 19155
rect 11323 19189 11375 19201
rect 11323 19155 11331 19189
rect 11365 19155 11375 19189
rect 11323 19027 11375 19155
rect 12321 19189 12373 19201
rect 12321 19155 12331 19189
rect 12365 19155 12373 19189
rect 12611 19189 12663 19201
rect 12321 19027 12373 19155
rect 12611 19155 12619 19189
rect 12653 19155 12663 19189
rect 12611 19087 12663 19155
rect 12611 19053 12619 19087
rect 12653 19053 12663 19087
rect 12611 19027 12663 19053
rect 13057 19189 13109 19201
rect 13057 19155 13067 19189
rect 13101 19155 13109 19189
rect 13057 19087 13109 19155
rect 13057 19053 13067 19087
rect 13101 19053 13109 19087
rect 13057 19027 13109 19053
rect 13163 19189 13215 19201
rect 13163 19155 13171 19189
rect 13205 19155 13215 19189
rect 13163 19027 13215 19155
rect 14161 19189 14213 19201
rect 14161 19155 14171 19189
rect 14205 19155 14213 19189
rect 14161 19027 14213 19155
rect 14267 19189 14319 19201
rect 14267 19155 14275 19189
rect 14309 19155 14319 19189
rect 14267 19027 14319 19155
rect 15265 19189 15317 19201
rect 15265 19155 15275 19189
rect 15309 19155 15317 19189
rect 15265 19027 15317 19155
rect 15371 19189 15423 19201
rect 15371 19155 15379 19189
rect 15413 19155 15423 19189
rect 15371 19027 15423 19155
rect 16369 19189 16421 19201
rect 16369 19155 16379 19189
rect 16413 19155 16421 19189
rect 16369 19027 16421 19155
rect 16475 19189 16527 19201
rect 16475 19155 16483 19189
rect 16517 19155 16527 19189
rect 16475 19027 16527 19155
rect 17473 19189 17525 19201
rect 17473 19155 17483 19189
rect 17517 19155 17525 19189
rect 17763 19189 17815 19201
rect 17473 19027 17525 19155
rect 17763 19155 17771 19189
rect 17805 19155 17815 19189
rect 17763 19027 17815 19155
rect 18761 19189 18813 19201
rect 18761 19155 18771 19189
rect 18805 19155 18813 19189
rect 18761 19027 18813 19155
rect 18867 19189 18919 19201
rect 18867 19155 18875 19189
rect 18909 19155 18919 19189
rect 18867 19027 18919 19155
rect 19865 19189 19917 19201
rect 19865 19155 19875 19189
rect 19909 19155 19917 19189
rect 19865 19027 19917 19155
rect 19971 19189 20023 19201
rect 19971 19155 19979 19189
rect 20013 19155 20023 19189
rect 19971 19094 20023 19155
rect 19971 19060 19979 19094
rect 20013 19060 20023 19094
rect 19971 19027 20023 19060
rect 20141 19189 20193 19201
rect 20141 19155 20151 19189
rect 20185 19155 20193 19189
rect 20141 19094 20193 19155
rect 20141 19060 20151 19094
rect 20185 19060 20193 19094
rect 20141 19027 20193 19060
rect 4975 18348 5027 18381
rect 4975 18314 4983 18348
rect 5017 18314 5027 18348
rect 4975 18253 5027 18314
rect 4975 18219 4983 18253
rect 5017 18219 5027 18253
rect 4975 18207 5027 18219
rect 5145 18348 5197 18381
rect 5145 18314 5155 18348
rect 5189 18314 5197 18348
rect 5145 18253 5197 18314
rect 5145 18219 5155 18253
rect 5189 18219 5197 18253
rect 5145 18207 5197 18219
rect 5435 18253 5487 18381
rect 5435 18219 5443 18253
rect 5477 18219 5487 18253
rect 5435 18207 5487 18219
rect 6433 18253 6485 18381
rect 6433 18219 6443 18253
rect 6477 18219 6485 18253
rect 6433 18207 6485 18219
rect 6539 18253 6591 18381
rect 6539 18219 6547 18253
rect 6581 18219 6591 18253
rect 6539 18207 6591 18219
rect 7537 18253 7589 18381
rect 7537 18219 7547 18253
rect 7581 18219 7589 18253
rect 7537 18207 7589 18219
rect 7643 18253 7695 18381
rect 7643 18219 7651 18253
rect 7685 18219 7695 18253
rect 7643 18207 7695 18219
rect 8641 18253 8693 18381
rect 8641 18219 8651 18253
rect 8685 18219 8693 18253
rect 8641 18207 8693 18219
rect 8747 18253 8799 18381
rect 8747 18219 8755 18253
rect 8789 18219 8799 18253
rect 8747 18207 8799 18219
rect 9745 18253 9797 18381
rect 9745 18219 9755 18253
rect 9789 18219 9797 18253
rect 10035 18355 10087 18381
rect 10035 18321 10043 18355
rect 10077 18321 10087 18355
rect 10035 18253 10087 18321
rect 9745 18207 9797 18219
rect 10035 18219 10043 18253
rect 10077 18219 10087 18253
rect 10035 18207 10087 18219
rect 10481 18355 10533 18381
rect 10481 18321 10491 18355
rect 10525 18321 10533 18355
rect 10481 18253 10533 18321
rect 10481 18219 10491 18253
rect 10525 18219 10533 18253
rect 10481 18207 10533 18219
rect 10587 18253 10639 18381
rect 10587 18219 10595 18253
rect 10629 18219 10639 18253
rect 10587 18207 10639 18219
rect 11585 18253 11637 18381
rect 11585 18219 11595 18253
rect 11629 18219 11637 18253
rect 11585 18207 11637 18219
rect 11691 18253 11743 18381
rect 11691 18219 11699 18253
rect 11733 18219 11743 18253
rect 11691 18207 11743 18219
rect 12689 18253 12741 18381
rect 12689 18219 12699 18253
rect 12733 18219 12741 18253
rect 12689 18207 12741 18219
rect 12795 18253 12847 18381
rect 12795 18219 12803 18253
rect 12837 18219 12847 18253
rect 12795 18207 12847 18219
rect 13793 18253 13845 18381
rect 13793 18219 13803 18253
rect 13837 18219 13845 18253
rect 13793 18207 13845 18219
rect 13899 18253 13951 18381
rect 13899 18219 13907 18253
rect 13941 18219 13951 18253
rect 13899 18207 13951 18219
rect 14897 18253 14949 18381
rect 14897 18219 14907 18253
rect 14941 18219 14949 18253
rect 15187 18355 15239 18381
rect 15187 18321 15195 18355
rect 15229 18321 15239 18355
rect 15187 18253 15239 18321
rect 14897 18207 14949 18219
rect 15187 18219 15195 18253
rect 15229 18219 15239 18253
rect 15187 18207 15239 18219
rect 15449 18355 15501 18381
rect 15449 18321 15459 18355
rect 15493 18321 15501 18355
rect 15449 18253 15501 18321
rect 15449 18219 15459 18253
rect 15493 18219 15501 18253
rect 15449 18207 15501 18219
rect 15555 18253 15607 18381
rect 15555 18219 15563 18253
rect 15597 18219 15607 18253
rect 15555 18207 15607 18219
rect 16553 18253 16605 18381
rect 16553 18219 16563 18253
rect 16597 18219 16605 18253
rect 16553 18207 16605 18219
rect 16659 18253 16711 18381
rect 16659 18219 16667 18253
rect 16701 18219 16711 18253
rect 16659 18207 16711 18219
rect 17657 18253 17709 18381
rect 17657 18219 17667 18253
rect 17701 18219 17709 18253
rect 17657 18207 17709 18219
rect 17763 18253 17815 18381
rect 17763 18219 17771 18253
rect 17805 18219 17815 18253
rect 17763 18207 17815 18219
rect 18761 18253 18813 18381
rect 18761 18219 18771 18253
rect 18805 18219 18813 18253
rect 18761 18207 18813 18219
rect 18867 18253 18919 18381
rect 18867 18219 18875 18253
rect 18909 18219 18919 18253
rect 18867 18207 18919 18219
rect 19865 18253 19917 18381
rect 19865 18219 19875 18253
rect 19909 18219 19917 18253
rect 19865 18207 19917 18219
rect 19971 18348 20023 18381
rect 19971 18314 19979 18348
rect 20013 18314 20023 18348
rect 19971 18253 20023 18314
rect 19971 18219 19979 18253
rect 20013 18219 20023 18253
rect 19971 18207 20023 18219
rect 20141 18348 20193 18381
rect 20141 18314 20151 18348
rect 20185 18314 20193 18348
rect 20141 18253 20193 18314
rect 20141 18219 20151 18253
rect 20185 18219 20193 18253
rect 20141 18207 20193 18219
rect 4975 18101 5027 18113
rect 4975 18067 4983 18101
rect 5017 18067 5027 18101
rect 4975 18006 5027 18067
rect 4975 17972 4983 18006
rect 5017 17972 5027 18006
rect 4975 17939 5027 17972
rect 5145 18101 5197 18113
rect 5145 18067 5155 18101
rect 5189 18067 5197 18101
rect 5145 18006 5197 18067
rect 5145 17972 5155 18006
rect 5189 17972 5197 18006
rect 5145 17939 5197 17972
rect 5435 18101 5487 18113
rect 5435 18067 5443 18101
rect 5477 18067 5487 18101
rect 5435 17999 5487 18067
rect 5435 17965 5443 17999
rect 5477 17965 5487 17999
rect 5435 17939 5487 17965
rect 6065 18101 6117 18113
rect 6065 18067 6075 18101
rect 6109 18067 6117 18101
rect 6065 17999 6117 18067
rect 6065 17965 6075 17999
rect 6109 17965 6117 17999
rect 6065 17939 6117 17965
rect 6171 18101 6223 18113
rect 6171 18067 6179 18101
rect 6213 18067 6223 18101
rect 6171 17939 6223 18067
rect 7169 18101 7221 18113
rect 7169 18067 7179 18101
rect 7213 18067 7221 18101
rect 7459 18101 7511 18113
rect 7169 17939 7221 18067
rect 7459 18067 7467 18101
rect 7501 18067 7511 18101
rect 7459 17999 7511 18067
rect 7459 17965 7467 17999
rect 7501 17965 7511 17999
rect 7459 17939 7511 17965
rect 7905 18101 7957 18113
rect 7905 18067 7915 18101
rect 7949 18067 7957 18101
rect 7905 17999 7957 18067
rect 7905 17965 7915 17999
rect 7949 17965 7957 17999
rect 7905 17939 7957 17965
rect 8011 18101 8063 18113
rect 8011 18067 8019 18101
rect 8053 18067 8063 18101
rect 8011 17939 8063 18067
rect 9009 18101 9061 18113
rect 9009 18067 9019 18101
rect 9053 18067 9061 18101
rect 9009 17939 9061 18067
rect 9115 18101 9167 18113
rect 9115 18067 9123 18101
rect 9157 18067 9167 18101
rect 9115 17939 9167 18067
rect 10113 18101 10165 18113
rect 10113 18067 10123 18101
rect 10157 18067 10165 18101
rect 10113 17939 10165 18067
rect 10219 18101 10271 18113
rect 10219 18067 10227 18101
rect 10261 18067 10271 18101
rect 10219 17939 10271 18067
rect 11217 18101 11269 18113
rect 11217 18067 11227 18101
rect 11261 18067 11269 18101
rect 11217 17939 11269 18067
rect 11323 18101 11375 18113
rect 11323 18067 11331 18101
rect 11365 18067 11375 18101
rect 11323 17939 11375 18067
rect 12321 18101 12373 18113
rect 12321 18067 12331 18101
rect 12365 18067 12373 18101
rect 12611 18101 12663 18113
rect 12321 17939 12373 18067
rect 12611 18067 12619 18101
rect 12653 18067 12663 18101
rect 12611 17999 12663 18067
rect 12611 17965 12619 17999
rect 12653 17965 12663 17999
rect 12611 17939 12663 17965
rect 13057 18101 13109 18113
rect 13057 18067 13067 18101
rect 13101 18067 13109 18101
rect 13057 17999 13109 18067
rect 13057 17965 13067 17999
rect 13101 17965 13109 17999
rect 13057 17939 13109 17965
rect 13163 18101 13215 18113
rect 13163 18067 13171 18101
rect 13205 18067 13215 18101
rect 13163 17939 13215 18067
rect 14161 18101 14213 18113
rect 14161 18067 14171 18101
rect 14205 18067 14213 18101
rect 14161 17939 14213 18067
rect 14267 18101 14319 18113
rect 14267 18067 14275 18101
rect 14309 18067 14319 18101
rect 14267 17939 14319 18067
rect 15265 18101 15317 18113
rect 15265 18067 15275 18101
rect 15309 18067 15317 18101
rect 15265 17939 15317 18067
rect 15371 18101 15423 18113
rect 15371 18067 15379 18101
rect 15413 18067 15423 18101
rect 15371 17939 15423 18067
rect 16369 18101 16421 18113
rect 16369 18067 16379 18101
rect 16413 18067 16421 18101
rect 16369 17939 16421 18067
rect 16475 18101 16527 18113
rect 16475 18067 16483 18101
rect 16517 18067 16527 18101
rect 16475 17939 16527 18067
rect 17473 18101 17525 18113
rect 17473 18067 17483 18101
rect 17517 18067 17525 18101
rect 17763 18101 17815 18113
rect 17473 17939 17525 18067
rect 17763 18067 17771 18101
rect 17805 18067 17815 18101
rect 17763 17939 17815 18067
rect 18761 18101 18813 18113
rect 18761 18067 18771 18101
rect 18805 18067 18813 18101
rect 18761 17939 18813 18067
rect 18867 18101 18919 18113
rect 18867 18067 18875 18101
rect 18909 18067 18919 18101
rect 18867 17939 18919 18067
rect 19865 18101 19917 18113
rect 19865 18067 19875 18101
rect 19909 18067 19917 18101
rect 19865 17939 19917 18067
rect 19971 18101 20023 18113
rect 19971 18067 19979 18101
rect 20013 18067 20023 18101
rect 19971 18006 20023 18067
rect 19971 17972 19979 18006
rect 20013 17972 20023 18006
rect 19971 17939 20023 17972
rect 20141 18101 20193 18113
rect 20141 18067 20151 18101
rect 20185 18067 20193 18101
rect 20141 18006 20193 18067
rect 20141 17972 20151 18006
rect 20185 17972 20193 18006
rect 20141 17939 20193 17972
rect 4975 17260 5027 17293
rect 4975 17226 4983 17260
rect 5017 17226 5027 17260
rect 4975 17165 5027 17226
rect 4975 17131 4983 17165
rect 5017 17131 5027 17165
rect 4975 17119 5027 17131
rect 5145 17260 5197 17293
rect 5145 17226 5155 17260
rect 5189 17226 5197 17260
rect 5145 17165 5197 17226
rect 5145 17131 5155 17165
rect 5189 17131 5197 17165
rect 5145 17119 5197 17131
rect 5435 17165 5487 17293
rect 5435 17131 5443 17165
rect 5477 17131 5487 17165
rect 5435 17119 5487 17131
rect 6433 17165 6485 17293
rect 6433 17131 6443 17165
rect 6477 17131 6485 17165
rect 6433 17119 6485 17131
rect 6539 17165 6591 17293
rect 6539 17131 6547 17165
rect 6581 17131 6591 17165
rect 6539 17119 6591 17131
rect 7537 17165 7589 17293
rect 7537 17131 7547 17165
rect 7581 17131 7589 17165
rect 7537 17119 7589 17131
rect 7643 17165 7695 17293
rect 7643 17131 7651 17165
rect 7685 17131 7695 17165
rect 7643 17119 7695 17131
rect 8641 17165 8693 17293
rect 8641 17131 8651 17165
rect 8685 17131 8693 17165
rect 8641 17119 8693 17131
rect 8747 17165 8799 17293
rect 8747 17131 8755 17165
rect 8789 17131 8799 17165
rect 8747 17119 8799 17131
rect 9745 17165 9797 17293
rect 9745 17131 9755 17165
rect 9789 17131 9797 17165
rect 10035 17267 10087 17293
rect 10035 17233 10043 17267
rect 10077 17233 10087 17267
rect 10035 17165 10087 17233
rect 9745 17119 9797 17131
rect 10035 17131 10043 17165
rect 10077 17131 10087 17165
rect 10035 17119 10087 17131
rect 10481 17267 10533 17293
rect 10481 17233 10491 17267
rect 10525 17233 10533 17267
rect 10481 17165 10533 17233
rect 10481 17131 10491 17165
rect 10525 17131 10533 17165
rect 10481 17119 10533 17131
rect 10587 17165 10639 17293
rect 10587 17131 10595 17165
rect 10629 17131 10639 17165
rect 10587 17119 10639 17131
rect 11585 17165 11637 17293
rect 11585 17131 11595 17165
rect 11629 17131 11637 17165
rect 11585 17119 11637 17131
rect 11691 17165 11743 17293
rect 11691 17131 11699 17165
rect 11733 17131 11743 17165
rect 11691 17119 11743 17131
rect 12689 17165 12741 17293
rect 12689 17131 12699 17165
rect 12733 17131 12741 17165
rect 12689 17119 12741 17131
rect 12795 17165 12847 17293
rect 12795 17131 12803 17165
rect 12837 17131 12847 17165
rect 12795 17119 12847 17131
rect 13793 17165 13845 17293
rect 13793 17131 13803 17165
rect 13837 17131 13845 17165
rect 13793 17119 13845 17131
rect 13899 17165 13951 17293
rect 13899 17131 13907 17165
rect 13941 17131 13951 17165
rect 13899 17119 13951 17131
rect 14897 17165 14949 17293
rect 14897 17131 14907 17165
rect 14941 17131 14949 17165
rect 15187 17267 15239 17293
rect 15187 17233 15195 17267
rect 15229 17233 15239 17267
rect 15187 17165 15239 17233
rect 14897 17119 14949 17131
rect 15187 17131 15195 17165
rect 15229 17131 15239 17165
rect 15187 17119 15239 17131
rect 15449 17267 15501 17293
rect 15449 17233 15459 17267
rect 15493 17233 15501 17267
rect 15449 17165 15501 17233
rect 15449 17131 15459 17165
rect 15493 17131 15501 17165
rect 15449 17119 15501 17131
rect 15555 17165 15607 17293
rect 15555 17131 15563 17165
rect 15597 17131 15607 17165
rect 15555 17119 15607 17131
rect 16553 17165 16605 17293
rect 16553 17131 16563 17165
rect 16597 17131 16605 17165
rect 16553 17119 16605 17131
rect 16659 17165 16711 17293
rect 16659 17131 16667 17165
rect 16701 17131 16711 17165
rect 16659 17119 16711 17131
rect 17657 17165 17709 17293
rect 17657 17131 17667 17165
rect 17701 17131 17709 17165
rect 17657 17119 17709 17131
rect 17763 17165 17815 17293
rect 17763 17131 17771 17165
rect 17805 17131 17815 17165
rect 17763 17119 17815 17131
rect 18761 17165 18813 17293
rect 18761 17131 18771 17165
rect 18805 17131 18813 17165
rect 18761 17119 18813 17131
rect 18867 17165 18919 17293
rect 18867 17131 18875 17165
rect 18909 17131 18919 17165
rect 18867 17119 18919 17131
rect 19865 17165 19917 17293
rect 19865 17131 19875 17165
rect 19909 17131 19917 17165
rect 19865 17119 19917 17131
rect 19971 17260 20023 17293
rect 19971 17226 19979 17260
rect 20013 17226 20023 17260
rect 19971 17165 20023 17226
rect 19971 17131 19979 17165
rect 20013 17131 20023 17165
rect 19971 17119 20023 17131
rect 20141 17260 20193 17293
rect 20141 17226 20151 17260
rect 20185 17226 20193 17260
rect 20141 17165 20193 17226
rect 20141 17131 20151 17165
rect 20185 17131 20193 17165
rect 20141 17119 20193 17131
rect 4975 17013 5027 17025
rect 4975 16979 4983 17013
rect 5017 16979 5027 17013
rect 4975 16918 5027 16979
rect 4975 16884 4983 16918
rect 5017 16884 5027 16918
rect 4975 16851 5027 16884
rect 5145 17013 5197 17025
rect 5145 16979 5155 17013
rect 5189 16979 5197 17013
rect 5145 16918 5197 16979
rect 5145 16884 5155 16918
rect 5189 16884 5197 16918
rect 5145 16851 5197 16884
rect 5435 17013 5487 17025
rect 5435 16979 5443 17013
rect 5477 16979 5487 17013
rect 5435 16911 5487 16979
rect 5435 16877 5443 16911
rect 5477 16877 5487 16911
rect 5435 16851 5487 16877
rect 6065 17013 6117 17025
rect 6065 16979 6075 17013
rect 6109 16979 6117 17013
rect 6065 16911 6117 16979
rect 6065 16877 6075 16911
rect 6109 16877 6117 16911
rect 6065 16851 6117 16877
rect 6171 17013 6223 17025
rect 6171 16979 6179 17013
rect 6213 16979 6223 17013
rect 6171 16851 6223 16979
rect 7169 17013 7221 17025
rect 7169 16979 7179 17013
rect 7213 16979 7221 17013
rect 7459 17013 7511 17025
rect 7169 16851 7221 16979
rect 7459 16979 7467 17013
rect 7501 16979 7511 17013
rect 7459 16911 7511 16979
rect 7459 16877 7467 16911
rect 7501 16877 7511 16911
rect 7459 16851 7511 16877
rect 7905 17013 7957 17025
rect 7905 16979 7915 17013
rect 7949 16979 7957 17013
rect 7905 16911 7957 16979
rect 7905 16877 7915 16911
rect 7949 16877 7957 16911
rect 7905 16851 7957 16877
rect 8011 17013 8063 17025
rect 8011 16979 8019 17013
rect 8053 16979 8063 17013
rect 8011 16851 8063 16979
rect 9009 17013 9061 17025
rect 9009 16979 9019 17013
rect 9053 16979 9061 17013
rect 9009 16851 9061 16979
rect 9115 17013 9167 17025
rect 9115 16979 9123 17013
rect 9157 16979 9167 17013
rect 9115 16851 9167 16979
rect 10113 17013 10165 17025
rect 10113 16979 10123 17013
rect 10157 16979 10165 17013
rect 10113 16851 10165 16979
rect 10219 17013 10271 17025
rect 10219 16979 10227 17013
rect 10261 16979 10271 17013
rect 10219 16851 10271 16979
rect 11217 17013 11269 17025
rect 11217 16979 11227 17013
rect 11261 16979 11269 17013
rect 11217 16851 11269 16979
rect 11323 17013 11375 17025
rect 11323 16979 11331 17013
rect 11365 16979 11375 17013
rect 11323 16851 11375 16979
rect 12321 17013 12373 17025
rect 12321 16979 12331 17013
rect 12365 16979 12373 17013
rect 12611 17013 12663 17025
rect 12321 16851 12373 16979
rect 12611 16979 12619 17013
rect 12653 16979 12663 17013
rect 12611 16911 12663 16979
rect 12611 16877 12619 16911
rect 12653 16877 12663 16911
rect 12611 16851 12663 16877
rect 13057 17013 13109 17025
rect 13057 16979 13067 17013
rect 13101 16979 13109 17013
rect 13057 16911 13109 16979
rect 13057 16877 13067 16911
rect 13101 16877 13109 16911
rect 13057 16851 13109 16877
rect 13163 17013 13215 17025
rect 13163 16979 13171 17013
rect 13205 16979 13215 17013
rect 13163 16851 13215 16979
rect 14161 17013 14213 17025
rect 14161 16979 14171 17013
rect 14205 16979 14213 17013
rect 14161 16851 14213 16979
rect 14267 17013 14319 17025
rect 14267 16979 14275 17013
rect 14309 16979 14319 17013
rect 14267 16851 14319 16979
rect 15265 17013 15317 17025
rect 15265 16979 15275 17013
rect 15309 16979 15317 17013
rect 15265 16851 15317 16979
rect 15371 17013 15423 17025
rect 15371 16979 15379 17013
rect 15413 16979 15423 17013
rect 15371 16851 15423 16979
rect 16369 17013 16421 17025
rect 16369 16979 16379 17013
rect 16413 16979 16421 17013
rect 16369 16851 16421 16979
rect 16475 17013 16527 17025
rect 16475 16979 16483 17013
rect 16517 16979 16527 17013
rect 16475 16851 16527 16979
rect 17473 17013 17525 17025
rect 17473 16979 17483 17013
rect 17517 16979 17525 17013
rect 17763 17013 17815 17025
rect 17473 16851 17525 16979
rect 17763 16979 17771 17013
rect 17805 16979 17815 17013
rect 17763 16851 17815 16979
rect 18761 17013 18813 17025
rect 18761 16979 18771 17013
rect 18805 16979 18813 17013
rect 18761 16851 18813 16979
rect 18867 17013 18919 17025
rect 18867 16979 18875 17013
rect 18909 16979 18919 17013
rect 18867 16851 18919 16979
rect 19865 17013 19917 17025
rect 19865 16979 19875 17013
rect 19909 16979 19917 17013
rect 19865 16851 19917 16979
rect 19971 17013 20023 17025
rect 19971 16979 19979 17013
rect 20013 16979 20023 17013
rect 19971 16918 20023 16979
rect 19971 16884 19979 16918
rect 20013 16884 20023 16918
rect 19971 16851 20023 16884
rect 20141 17013 20193 17025
rect 20141 16979 20151 17013
rect 20185 16979 20193 17013
rect 20141 16918 20193 16979
rect 20141 16884 20151 16918
rect 20185 16884 20193 16918
rect 20141 16851 20193 16884
rect 4975 16172 5027 16205
rect 4975 16138 4983 16172
rect 5017 16138 5027 16172
rect 4975 16077 5027 16138
rect 4975 16043 4983 16077
rect 5017 16043 5027 16077
rect 4975 16031 5027 16043
rect 5145 16172 5197 16205
rect 5145 16138 5155 16172
rect 5189 16138 5197 16172
rect 5145 16077 5197 16138
rect 5145 16043 5155 16077
rect 5189 16043 5197 16077
rect 5145 16031 5197 16043
rect 5435 16077 5487 16205
rect 5435 16043 5443 16077
rect 5477 16043 5487 16077
rect 5435 16031 5487 16043
rect 6433 16077 6485 16205
rect 6433 16043 6443 16077
rect 6477 16043 6485 16077
rect 6433 16031 6485 16043
rect 6539 16077 6591 16205
rect 6539 16043 6547 16077
rect 6581 16043 6591 16077
rect 6539 16031 6591 16043
rect 7537 16077 7589 16205
rect 7537 16043 7547 16077
rect 7581 16043 7589 16077
rect 7537 16031 7589 16043
rect 7643 16077 7695 16205
rect 7643 16043 7651 16077
rect 7685 16043 7695 16077
rect 7643 16031 7695 16043
rect 8641 16077 8693 16205
rect 8641 16043 8651 16077
rect 8685 16043 8693 16077
rect 8641 16031 8693 16043
rect 8747 16077 8799 16205
rect 8747 16043 8755 16077
rect 8789 16043 8799 16077
rect 8747 16031 8799 16043
rect 9745 16077 9797 16205
rect 9745 16043 9755 16077
rect 9789 16043 9797 16077
rect 10035 16179 10087 16205
rect 10035 16145 10043 16179
rect 10077 16145 10087 16179
rect 10035 16077 10087 16145
rect 9745 16031 9797 16043
rect 10035 16043 10043 16077
rect 10077 16043 10087 16077
rect 10035 16031 10087 16043
rect 10481 16179 10533 16205
rect 10481 16145 10491 16179
rect 10525 16145 10533 16179
rect 10481 16077 10533 16145
rect 10481 16043 10491 16077
rect 10525 16043 10533 16077
rect 10481 16031 10533 16043
rect 10587 16077 10639 16205
rect 10587 16043 10595 16077
rect 10629 16043 10639 16077
rect 10587 16031 10639 16043
rect 11585 16077 11637 16205
rect 11585 16043 11595 16077
rect 11629 16043 11637 16077
rect 11585 16031 11637 16043
rect 11691 16077 11743 16205
rect 11691 16043 11699 16077
rect 11733 16043 11743 16077
rect 11691 16031 11743 16043
rect 12689 16077 12741 16205
rect 12689 16043 12699 16077
rect 12733 16043 12741 16077
rect 12689 16031 12741 16043
rect 12795 16077 12847 16205
rect 12795 16043 12803 16077
rect 12837 16043 12847 16077
rect 12795 16031 12847 16043
rect 13793 16077 13845 16205
rect 13793 16043 13803 16077
rect 13837 16043 13845 16077
rect 13793 16031 13845 16043
rect 13899 16077 13951 16205
rect 13899 16043 13907 16077
rect 13941 16043 13951 16077
rect 13899 16031 13951 16043
rect 14897 16077 14949 16205
rect 14897 16043 14907 16077
rect 14941 16043 14949 16077
rect 15187 16179 15239 16205
rect 15187 16145 15195 16179
rect 15229 16145 15239 16179
rect 15187 16077 15239 16145
rect 14897 16031 14949 16043
rect 15187 16043 15195 16077
rect 15229 16043 15239 16077
rect 15187 16031 15239 16043
rect 15449 16179 15501 16205
rect 15449 16145 15459 16179
rect 15493 16145 15501 16179
rect 15449 16077 15501 16145
rect 15449 16043 15459 16077
rect 15493 16043 15501 16077
rect 15449 16031 15501 16043
rect 15555 16077 15607 16205
rect 15555 16043 15563 16077
rect 15597 16043 15607 16077
rect 15555 16031 15607 16043
rect 16553 16077 16605 16205
rect 16553 16043 16563 16077
rect 16597 16043 16605 16077
rect 16553 16031 16605 16043
rect 16659 16077 16711 16205
rect 16659 16043 16667 16077
rect 16701 16043 16711 16077
rect 16659 16031 16711 16043
rect 17657 16077 17709 16205
rect 17657 16043 17667 16077
rect 17701 16043 17709 16077
rect 17657 16031 17709 16043
rect 17763 16077 17815 16205
rect 17763 16043 17771 16077
rect 17805 16043 17815 16077
rect 17763 16031 17815 16043
rect 18761 16077 18813 16205
rect 18761 16043 18771 16077
rect 18805 16043 18813 16077
rect 18761 16031 18813 16043
rect 18867 16077 18919 16205
rect 18867 16043 18875 16077
rect 18909 16043 18919 16077
rect 18867 16031 18919 16043
rect 19865 16077 19917 16205
rect 19865 16043 19875 16077
rect 19909 16043 19917 16077
rect 19865 16031 19917 16043
rect 19971 16172 20023 16205
rect 19971 16138 19979 16172
rect 20013 16138 20023 16172
rect 19971 16077 20023 16138
rect 19971 16043 19979 16077
rect 20013 16043 20023 16077
rect 19971 16031 20023 16043
rect 20141 16172 20193 16205
rect 20141 16138 20151 16172
rect 20185 16138 20193 16172
rect 20141 16077 20193 16138
rect 20141 16043 20151 16077
rect 20185 16043 20193 16077
rect 20141 16031 20193 16043
rect 4975 15925 5027 15937
rect 4975 15891 4983 15925
rect 5017 15891 5027 15925
rect 4975 15830 5027 15891
rect 4975 15796 4983 15830
rect 5017 15796 5027 15830
rect 4975 15763 5027 15796
rect 5145 15925 5197 15937
rect 5145 15891 5155 15925
rect 5189 15891 5197 15925
rect 5145 15830 5197 15891
rect 5145 15796 5155 15830
rect 5189 15796 5197 15830
rect 5145 15763 5197 15796
rect 5435 15925 5487 15937
rect 5435 15891 5443 15925
rect 5477 15891 5487 15925
rect 5435 15823 5487 15891
rect 5435 15789 5443 15823
rect 5477 15789 5487 15823
rect 5435 15763 5487 15789
rect 6065 15925 6117 15937
rect 6065 15891 6075 15925
rect 6109 15891 6117 15925
rect 6065 15823 6117 15891
rect 6065 15789 6075 15823
rect 6109 15789 6117 15823
rect 6065 15763 6117 15789
rect 6171 15925 6223 15937
rect 6171 15891 6179 15925
rect 6213 15891 6223 15925
rect 6171 15763 6223 15891
rect 7169 15925 7221 15937
rect 7169 15891 7179 15925
rect 7213 15891 7221 15925
rect 7459 15925 7511 15937
rect 7169 15763 7221 15891
rect 7459 15891 7467 15925
rect 7501 15891 7511 15925
rect 7459 15823 7511 15891
rect 7459 15789 7467 15823
rect 7501 15789 7511 15823
rect 7459 15763 7511 15789
rect 7905 15925 7957 15937
rect 7905 15891 7915 15925
rect 7949 15891 7957 15925
rect 7905 15823 7957 15891
rect 7905 15789 7915 15823
rect 7949 15789 7957 15823
rect 7905 15763 7957 15789
rect 8011 15925 8063 15937
rect 8011 15891 8019 15925
rect 8053 15891 8063 15925
rect 8011 15763 8063 15891
rect 9009 15925 9061 15937
rect 9009 15891 9019 15925
rect 9053 15891 9061 15925
rect 9009 15763 9061 15891
rect 9115 15925 9167 15937
rect 9115 15891 9123 15925
rect 9157 15891 9167 15925
rect 9115 15763 9167 15891
rect 10113 15925 10165 15937
rect 10113 15891 10123 15925
rect 10157 15891 10165 15925
rect 10113 15763 10165 15891
rect 10219 15925 10271 15937
rect 10219 15891 10227 15925
rect 10261 15891 10271 15925
rect 10219 15763 10271 15891
rect 11217 15925 11269 15937
rect 11217 15891 11227 15925
rect 11261 15891 11269 15925
rect 11217 15763 11269 15891
rect 11323 15925 11375 15937
rect 11323 15891 11331 15925
rect 11365 15891 11375 15925
rect 11323 15763 11375 15891
rect 12321 15925 12373 15937
rect 12321 15891 12331 15925
rect 12365 15891 12373 15925
rect 12611 15925 12663 15937
rect 12321 15763 12373 15891
rect 12611 15891 12619 15925
rect 12653 15891 12663 15925
rect 12611 15823 12663 15891
rect 12611 15789 12619 15823
rect 12653 15789 12663 15823
rect 12611 15763 12663 15789
rect 13057 15925 13109 15937
rect 13057 15891 13067 15925
rect 13101 15891 13109 15925
rect 13057 15823 13109 15891
rect 13057 15789 13067 15823
rect 13101 15789 13109 15823
rect 13057 15763 13109 15789
rect 13163 15925 13215 15937
rect 13163 15891 13171 15925
rect 13205 15891 13215 15925
rect 13163 15763 13215 15891
rect 14161 15925 14213 15937
rect 14161 15891 14171 15925
rect 14205 15891 14213 15925
rect 14161 15763 14213 15891
rect 14267 15925 14319 15937
rect 14267 15891 14275 15925
rect 14309 15891 14319 15925
rect 14267 15763 14319 15891
rect 15265 15925 15317 15937
rect 15265 15891 15275 15925
rect 15309 15891 15317 15925
rect 15265 15763 15317 15891
rect 15371 15925 15423 15937
rect 15371 15891 15379 15925
rect 15413 15891 15423 15925
rect 15371 15763 15423 15891
rect 16369 15925 16421 15937
rect 16369 15891 16379 15925
rect 16413 15891 16421 15925
rect 16369 15763 16421 15891
rect 16475 15925 16527 15937
rect 16475 15891 16483 15925
rect 16517 15891 16527 15925
rect 16475 15763 16527 15891
rect 17473 15925 17525 15937
rect 17473 15891 17483 15925
rect 17517 15891 17525 15925
rect 17763 15925 17815 15937
rect 17473 15763 17525 15891
rect 17763 15891 17771 15925
rect 17805 15891 17815 15925
rect 17763 15763 17815 15891
rect 18761 15925 18813 15937
rect 18761 15891 18771 15925
rect 18805 15891 18813 15925
rect 18761 15763 18813 15891
rect 18867 15925 18919 15937
rect 18867 15891 18875 15925
rect 18909 15891 18919 15925
rect 18867 15763 18919 15891
rect 19865 15925 19917 15937
rect 19865 15891 19875 15925
rect 19909 15891 19917 15925
rect 19865 15763 19917 15891
rect 19971 15925 20023 15937
rect 19971 15891 19979 15925
rect 20013 15891 20023 15925
rect 19971 15830 20023 15891
rect 19971 15796 19979 15830
rect 20013 15796 20023 15830
rect 19971 15763 20023 15796
rect 20141 15925 20193 15937
rect 20141 15891 20151 15925
rect 20185 15891 20193 15925
rect 20141 15830 20193 15891
rect 20141 15796 20151 15830
rect 20185 15796 20193 15830
rect 20141 15763 20193 15796
rect 4975 15084 5027 15117
rect 4975 15050 4983 15084
rect 5017 15050 5027 15084
rect 4975 14989 5027 15050
rect 4975 14955 4983 14989
rect 5017 14955 5027 14989
rect 4975 14943 5027 14955
rect 5145 15084 5197 15117
rect 5145 15050 5155 15084
rect 5189 15050 5197 15084
rect 5145 14989 5197 15050
rect 5145 14955 5155 14989
rect 5189 14955 5197 14989
rect 5145 14943 5197 14955
rect 5435 14989 5487 15117
rect 5435 14955 5443 14989
rect 5477 14955 5487 14989
rect 5435 14943 5487 14955
rect 6433 14989 6485 15117
rect 6433 14955 6443 14989
rect 6477 14955 6485 14989
rect 6433 14943 6485 14955
rect 6539 14989 6591 15117
rect 6539 14955 6547 14989
rect 6581 14955 6591 14989
rect 6539 14943 6591 14955
rect 7537 14989 7589 15117
rect 7537 14955 7547 14989
rect 7581 14955 7589 14989
rect 7537 14943 7589 14955
rect 7643 14989 7695 15117
rect 7643 14955 7651 14989
rect 7685 14955 7695 14989
rect 7643 14943 7695 14955
rect 8641 14989 8693 15117
rect 8641 14955 8651 14989
rect 8685 14955 8693 14989
rect 8641 14943 8693 14955
rect 8747 14989 8799 15117
rect 8747 14955 8755 14989
rect 8789 14955 8799 14989
rect 8747 14943 8799 14955
rect 9745 14989 9797 15117
rect 9745 14955 9755 14989
rect 9789 14955 9797 14989
rect 10035 15091 10087 15117
rect 10035 15057 10043 15091
rect 10077 15057 10087 15091
rect 10035 14989 10087 15057
rect 9745 14943 9797 14955
rect 10035 14955 10043 14989
rect 10077 14955 10087 14989
rect 10035 14943 10087 14955
rect 10481 15091 10533 15117
rect 10481 15057 10491 15091
rect 10525 15057 10533 15091
rect 10481 14989 10533 15057
rect 10481 14955 10491 14989
rect 10525 14955 10533 14989
rect 10481 14943 10533 14955
rect 10587 14989 10639 15117
rect 10587 14955 10595 14989
rect 10629 14955 10639 14989
rect 10587 14943 10639 14955
rect 11585 14989 11637 15117
rect 11585 14955 11595 14989
rect 11629 14955 11637 14989
rect 11585 14943 11637 14955
rect 11691 14989 11743 15117
rect 11691 14955 11699 14989
rect 11733 14955 11743 14989
rect 11691 14943 11743 14955
rect 12689 14989 12741 15117
rect 13326 15027 13376 15143
rect 12689 14955 12699 14989
rect 12733 14955 12741 14989
rect 12689 14943 12741 14955
rect 12817 15015 12869 15027
rect 12817 14981 12825 15015
rect 12859 14981 12869 15015
rect 12817 14943 12869 14981
rect 12899 14989 12953 15027
rect 12899 14955 12909 14989
rect 12943 14955 12953 14989
rect 12899 14943 12953 14955
rect 13053 15015 13105 15027
rect 13053 14981 13063 15015
rect 13097 14981 13105 15015
rect 13053 14943 13105 14981
rect 13159 15015 13211 15027
rect 13159 14981 13167 15015
rect 13201 14981 13211 15015
rect 13159 14943 13211 14981
rect 13311 14989 13376 15027
rect 13311 14955 13326 14989
rect 13360 14955 13376 14989
rect 13311 14943 13376 14955
rect 13406 15015 13458 15143
rect 13406 14981 13416 15015
rect 13450 14981 13458 15015
rect 13406 14943 13458 14981
rect 13531 15091 13583 15117
rect 13531 15057 13539 15091
rect 13573 15057 13583 15091
rect 13531 14989 13583 15057
rect 13531 14955 13539 14989
rect 13573 14955 13583 14989
rect 13531 14943 13583 14955
rect 13793 15091 13845 15117
rect 13793 15057 13803 15091
rect 13837 15057 13845 15091
rect 13793 14989 13845 15057
rect 13793 14955 13803 14989
rect 13837 14955 13845 14989
rect 13793 14943 13845 14955
rect 13899 14989 13951 15117
rect 13899 14955 13907 14989
rect 13941 14955 13951 14989
rect 13899 14943 13951 14955
rect 14897 14989 14949 15117
rect 14897 14955 14907 14989
rect 14941 14955 14949 14989
rect 15095 15084 15147 15117
rect 15095 15050 15103 15084
rect 15137 15050 15147 15084
rect 15095 14989 15147 15050
rect 14897 14943 14949 14955
rect 15095 14955 15103 14989
rect 15137 14955 15147 14989
rect 15095 14943 15147 14955
rect 15265 15084 15317 15117
rect 15265 15050 15275 15084
rect 15309 15050 15317 15084
rect 15265 14989 15317 15050
rect 15902 15027 15952 15143
rect 15265 14955 15275 14989
rect 15309 14955 15317 14989
rect 15265 14943 15317 14955
rect 15393 15015 15445 15027
rect 15393 14981 15401 15015
rect 15435 14981 15445 15015
rect 15393 14943 15445 14981
rect 15475 14989 15529 15027
rect 15475 14955 15485 14989
rect 15519 14955 15529 14989
rect 15475 14943 15529 14955
rect 15629 15015 15681 15027
rect 15629 14981 15639 15015
rect 15673 14981 15681 15015
rect 15629 14943 15681 14981
rect 15735 15015 15787 15027
rect 15735 14981 15743 15015
rect 15777 14981 15787 15015
rect 15735 14943 15787 14981
rect 15887 14989 15952 15027
rect 15887 14955 15902 14989
rect 15936 14955 15952 14989
rect 15887 14943 15952 14955
rect 15982 15015 16034 15143
rect 15982 14981 15992 15015
rect 16026 14981 16034 15015
rect 15982 14943 16034 14981
rect 16107 15091 16159 15117
rect 16107 15057 16115 15091
rect 16149 15057 16159 15091
rect 16107 14989 16159 15057
rect 16107 14955 16115 14989
rect 16149 14955 16159 14989
rect 16107 14943 16159 14955
rect 16553 15091 16605 15117
rect 16553 15057 16563 15091
rect 16597 15057 16605 15091
rect 16553 14989 16605 15057
rect 16553 14955 16563 14989
rect 16597 14955 16605 14989
rect 16553 14943 16605 14955
rect 16659 14989 16711 15117
rect 16659 14955 16667 14989
rect 16701 14955 16711 14989
rect 16659 14943 16711 14955
rect 17657 14989 17709 15117
rect 17657 14955 17667 14989
rect 17701 14955 17709 14989
rect 17657 14943 17709 14955
rect 17763 14989 17815 15117
rect 17763 14955 17771 14989
rect 17805 14955 17815 14989
rect 17763 14943 17815 14955
rect 18761 14989 18813 15117
rect 18761 14955 18771 14989
rect 18805 14955 18813 14989
rect 18761 14943 18813 14955
rect 18867 14989 18919 15117
rect 18867 14955 18875 14989
rect 18909 14955 18919 14989
rect 18867 14943 18919 14955
rect 19865 14989 19917 15117
rect 19865 14955 19875 14989
rect 19909 14955 19917 14989
rect 19865 14943 19917 14955
rect 19971 15084 20023 15117
rect 19971 15050 19979 15084
rect 20013 15050 20023 15084
rect 19971 14989 20023 15050
rect 19971 14955 19979 14989
rect 20013 14955 20023 14989
rect 19971 14943 20023 14955
rect 20141 15084 20193 15117
rect 20141 15050 20151 15084
rect 20185 15050 20193 15084
rect 20141 14989 20193 15050
rect 20141 14955 20151 14989
rect 20185 14955 20193 14989
rect 20141 14943 20193 14955
rect 4975 14837 5027 14849
rect 4975 14803 4983 14837
rect 5017 14803 5027 14837
rect 4975 14742 5027 14803
rect 4975 14708 4983 14742
rect 5017 14708 5027 14742
rect 4975 14675 5027 14708
rect 5145 14837 5197 14849
rect 5145 14803 5155 14837
rect 5189 14803 5197 14837
rect 5145 14742 5197 14803
rect 5145 14708 5155 14742
rect 5189 14708 5197 14742
rect 5145 14675 5197 14708
rect 5435 14837 5487 14849
rect 5435 14803 5443 14837
rect 5477 14803 5487 14837
rect 5435 14735 5487 14803
rect 5435 14701 5443 14735
rect 5477 14701 5487 14735
rect 5435 14675 5487 14701
rect 6065 14837 6117 14849
rect 6065 14803 6075 14837
rect 6109 14803 6117 14837
rect 6065 14735 6117 14803
rect 6065 14701 6075 14735
rect 6109 14701 6117 14735
rect 6065 14675 6117 14701
rect 6171 14837 6223 14849
rect 6171 14803 6179 14837
rect 6213 14803 6223 14837
rect 6171 14675 6223 14803
rect 7169 14837 7221 14849
rect 7169 14803 7179 14837
rect 7213 14803 7221 14837
rect 7367 14837 7419 14849
rect 7169 14675 7221 14803
rect 7367 14803 7375 14837
rect 7409 14803 7419 14837
rect 7367 14675 7419 14803
rect 8365 14837 8417 14849
rect 8365 14803 8375 14837
rect 8409 14803 8417 14837
rect 8365 14675 8417 14803
rect 8471 14837 8523 14849
rect 8471 14803 8479 14837
rect 8513 14803 8523 14837
rect 8471 14675 8523 14803
rect 9469 14837 9521 14849
rect 9469 14803 9479 14837
rect 9513 14803 9521 14837
rect 9469 14675 9521 14803
rect 9575 14837 9627 14849
rect 9575 14803 9583 14837
rect 9617 14803 9627 14837
rect 9575 14675 9627 14803
rect 10573 14837 10625 14849
rect 10573 14803 10583 14837
rect 10617 14803 10625 14837
rect 11319 14837 11371 14849
rect 11319 14810 11327 14837
rect 10573 14675 10625 14803
rect 10721 14777 10777 14810
rect 10721 14743 10733 14777
rect 10767 14743 10777 14777
rect 10721 14726 10777 14743
rect 10807 14777 10873 14810
rect 10807 14743 10819 14777
rect 10853 14743 10873 14777
rect 10807 14726 10873 14743
rect 10903 14726 10945 14810
rect 10975 14777 11159 14810
rect 10975 14743 11016 14777
rect 11050 14743 11091 14777
rect 11125 14743 11159 14777
rect 10975 14726 11159 14743
rect 11189 14726 11262 14810
rect 11292 14803 11327 14810
rect 11361 14803 11371 14837
rect 11292 14769 11371 14803
rect 11292 14735 11327 14769
rect 11361 14735 11371 14769
rect 11292 14726 11371 14735
rect 11319 14701 11371 14726
rect 11319 14667 11327 14701
rect 11361 14667 11371 14701
rect 11319 14649 11371 14667
rect 11401 14837 11453 14849
rect 11401 14803 11411 14837
rect 11445 14803 11453 14837
rect 11401 14769 11453 14803
rect 11401 14735 11411 14769
rect 11445 14735 11453 14769
rect 11401 14701 11453 14735
rect 11401 14667 11411 14701
rect 11445 14667 11453 14701
rect 11691 14837 11743 14849
rect 11691 14803 11699 14837
rect 11733 14803 11743 14837
rect 11691 14735 11743 14803
rect 11691 14701 11699 14735
rect 11733 14701 11743 14735
rect 11691 14675 11743 14701
rect 12321 14837 12373 14849
rect 12321 14803 12331 14837
rect 12365 14803 12373 14837
rect 13343 14837 13395 14849
rect 12321 14735 12373 14803
rect 12321 14701 12331 14735
rect 12365 14701 12373 14735
rect 12321 14675 12373 14701
rect 13343 14810 13351 14837
rect 12745 14777 12801 14810
rect 12745 14743 12757 14777
rect 12791 14743 12801 14777
rect 12745 14726 12801 14743
rect 12831 14777 12897 14810
rect 12831 14743 12843 14777
rect 12877 14743 12897 14777
rect 12831 14726 12897 14743
rect 12927 14726 12969 14810
rect 12999 14777 13183 14810
rect 12999 14743 13040 14777
rect 13074 14743 13115 14777
rect 13149 14743 13183 14777
rect 12999 14726 13183 14743
rect 13213 14726 13286 14810
rect 13316 14803 13351 14810
rect 13385 14803 13395 14837
rect 13316 14769 13395 14803
rect 13316 14735 13351 14769
rect 13385 14735 13395 14769
rect 13316 14726 13395 14735
rect 11401 14649 11453 14667
rect 13343 14701 13395 14726
rect 13343 14667 13351 14701
rect 13385 14667 13395 14701
rect 13343 14649 13395 14667
rect 13425 14837 13477 14849
rect 13425 14803 13435 14837
rect 13469 14803 13477 14837
rect 13425 14769 13477 14803
rect 13425 14735 13435 14769
rect 13469 14735 13477 14769
rect 13425 14701 13477 14735
rect 13425 14667 13435 14701
rect 13469 14667 13477 14701
rect 13531 14837 13583 14849
rect 13531 14803 13539 14837
rect 13573 14803 13583 14837
rect 13531 14735 13583 14803
rect 13531 14701 13539 14735
rect 13573 14701 13583 14735
rect 13531 14675 13583 14701
rect 14161 14837 14213 14849
rect 14161 14803 14171 14837
rect 14205 14803 14213 14837
rect 14161 14735 14213 14803
rect 14161 14701 14171 14735
rect 14205 14701 14213 14735
rect 14161 14675 14213 14701
rect 14267 14829 14319 14849
rect 14267 14795 14275 14829
rect 14309 14795 14319 14829
rect 14267 14761 14319 14795
rect 14267 14727 14275 14761
rect 14309 14727 14319 14761
rect 14267 14691 14319 14727
rect 14349 14829 14407 14849
rect 14349 14795 14361 14829
rect 14395 14795 14407 14829
rect 14349 14761 14407 14795
rect 14349 14727 14361 14761
rect 14395 14727 14407 14761
rect 14349 14691 14407 14727
rect 14437 14829 14489 14849
rect 14437 14795 14447 14829
rect 14481 14795 14489 14829
rect 14437 14748 14489 14795
rect 14437 14714 14447 14748
rect 14481 14714 14489 14748
rect 14437 14691 14489 14714
rect 14543 14801 14595 14849
rect 14543 14767 14551 14801
rect 14585 14767 14595 14801
rect 14543 14733 14595 14767
rect 14543 14699 14551 14733
rect 14585 14699 14595 14733
rect 13425 14649 13477 14667
rect 14543 14649 14595 14699
rect 14625 14837 14691 14849
rect 14625 14803 14635 14837
rect 14669 14803 14691 14837
rect 14625 14769 14691 14803
rect 14625 14735 14635 14769
rect 14669 14735 14691 14769
rect 14756 14837 14810 14849
rect 14756 14803 14764 14837
rect 14798 14803 14810 14837
rect 14756 14765 14810 14803
rect 14840 14811 14894 14849
rect 14840 14777 14850 14811
rect 14884 14777 14894 14811
rect 14840 14765 14894 14777
rect 14924 14837 15002 14849
rect 14924 14803 14934 14837
rect 14968 14803 15002 14837
rect 14924 14765 15002 14803
rect 15032 14765 15086 14849
rect 15116 14836 15172 14849
rect 15116 14802 15126 14836
rect 15160 14802 15172 14836
rect 15116 14765 15172 14802
rect 15202 14829 15271 14849
rect 15202 14795 15223 14829
rect 15257 14795 15271 14829
rect 15202 14765 15271 14795
rect 14625 14721 14691 14735
rect 14625 14649 14675 14721
rect 15217 14681 15271 14765
rect 15301 14837 15353 14849
rect 15301 14803 15311 14837
rect 15345 14803 15353 14837
rect 15301 14681 15353 14803
rect 15416 14811 15468 14849
rect 15416 14777 15424 14811
rect 15458 14777 15468 14811
rect 15416 14765 15468 14777
rect 15498 14827 15565 14849
rect 15498 14793 15508 14827
rect 15542 14793 15565 14827
rect 15498 14765 15565 14793
rect 15595 14811 15705 14849
rect 15595 14777 15605 14811
rect 15639 14777 15705 14811
rect 15595 14765 15705 14777
rect 15735 14835 15804 14849
rect 15735 14801 15759 14835
rect 15793 14801 15804 14835
rect 15735 14765 15804 14801
rect 15834 14829 15896 14849
rect 15834 14795 15852 14829
rect 15886 14795 15896 14829
rect 15834 14765 15896 14795
rect 15926 14837 15978 14849
rect 15926 14803 15936 14837
rect 15970 14803 15978 14837
rect 15926 14765 15978 14803
rect 16111 14829 16163 14843
rect 16111 14795 16119 14829
rect 16153 14795 16163 14829
rect 16111 14761 16163 14795
rect 16111 14727 16119 14761
rect 16153 14727 16163 14761
rect 16111 14715 16163 14727
rect 16193 14813 16247 14843
rect 16193 14779 16203 14813
rect 16237 14779 16247 14813
rect 16193 14715 16247 14779
rect 16277 14829 16329 14843
rect 16277 14795 16287 14829
rect 16321 14795 16329 14829
rect 16277 14761 16329 14795
rect 16277 14727 16287 14761
rect 16321 14727 16329 14761
rect 16277 14715 16329 14727
rect 16475 14837 16527 14849
rect 16475 14803 16483 14837
rect 16517 14803 16527 14837
rect 16475 14675 16527 14803
rect 17473 14837 17525 14849
rect 17473 14803 17483 14837
rect 17517 14803 17525 14837
rect 17763 14837 17815 14849
rect 17473 14675 17525 14803
rect 17763 14803 17771 14837
rect 17805 14803 17815 14837
rect 17763 14675 17815 14803
rect 18761 14837 18813 14849
rect 18761 14803 18771 14837
rect 18805 14803 18813 14837
rect 18761 14675 18813 14803
rect 18867 14837 18919 14849
rect 18867 14803 18875 14837
rect 18909 14803 18919 14837
rect 18867 14675 18919 14803
rect 19865 14837 19917 14849
rect 19865 14803 19875 14837
rect 19909 14803 19917 14837
rect 19865 14675 19917 14803
rect 19971 14837 20023 14849
rect 19971 14803 19979 14837
rect 20013 14803 20023 14837
rect 19971 14742 20023 14803
rect 19971 14708 19979 14742
rect 20013 14708 20023 14742
rect 19971 14675 20023 14708
rect 20141 14837 20193 14849
rect 20141 14803 20151 14837
rect 20185 14803 20193 14837
rect 20141 14742 20193 14803
rect 20141 14708 20151 14742
rect 20185 14708 20193 14742
rect 20141 14675 20193 14708
rect 4975 13996 5027 14029
rect 4975 13962 4983 13996
rect 5017 13962 5027 13996
rect 4975 13901 5027 13962
rect 4975 13867 4983 13901
rect 5017 13867 5027 13901
rect 4975 13855 5027 13867
rect 5145 13996 5197 14029
rect 5145 13962 5155 13996
rect 5189 13962 5197 13996
rect 5145 13901 5197 13962
rect 5145 13867 5155 13901
rect 5189 13867 5197 13901
rect 5145 13855 5197 13867
rect 5435 13901 5487 14029
rect 5435 13867 5443 13901
rect 5477 13867 5487 13901
rect 5435 13855 5487 13867
rect 6433 13901 6485 14029
rect 6433 13867 6443 13901
rect 6477 13867 6485 13901
rect 6433 13855 6485 13867
rect 6539 13901 6591 14029
rect 6539 13867 6547 13901
rect 6581 13867 6591 13901
rect 6539 13855 6591 13867
rect 7537 13901 7589 14029
rect 7537 13867 7547 13901
rect 7581 13867 7589 13901
rect 7537 13855 7589 13867
rect 7643 13901 7695 14029
rect 7643 13867 7651 13901
rect 7685 13867 7695 13901
rect 7643 13855 7695 13867
rect 8641 13901 8693 14029
rect 8641 13867 8651 13901
rect 8685 13867 8693 13901
rect 8641 13855 8693 13867
rect 8747 13901 8799 14029
rect 8747 13867 8755 13901
rect 8789 13867 8799 13901
rect 8747 13855 8799 13867
rect 9745 13901 9797 14029
rect 9745 13867 9755 13901
rect 9789 13867 9797 13901
rect 10127 14005 10179 14055
rect 10127 13971 10135 14005
rect 10169 13971 10179 14005
rect 10127 13937 10179 13971
rect 10127 13903 10135 13937
rect 10169 13903 10179 13937
rect 9745 13855 9797 13867
rect 10127 13855 10179 13903
rect 10209 13983 10259 14055
rect 10209 13969 10275 13983
rect 10209 13935 10219 13969
rect 10253 13935 10275 13969
rect 10801 13939 10855 14023
rect 10209 13901 10275 13935
rect 10209 13867 10219 13901
rect 10253 13867 10275 13901
rect 10209 13855 10275 13867
rect 10340 13901 10394 13939
rect 10340 13867 10348 13901
rect 10382 13867 10394 13901
rect 10340 13855 10394 13867
rect 10424 13927 10478 13939
rect 10424 13893 10434 13927
rect 10468 13893 10478 13927
rect 10424 13855 10478 13893
rect 10508 13901 10586 13939
rect 10508 13867 10518 13901
rect 10552 13867 10586 13901
rect 10508 13855 10586 13867
rect 10616 13855 10670 13939
rect 10700 13902 10756 13939
rect 10700 13868 10710 13902
rect 10744 13868 10756 13902
rect 10700 13855 10756 13868
rect 10786 13909 10855 13939
rect 10786 13875 10807 13909
rect 10841 13875 10855 13909
rect 10786 13855 10855 13875
rect 10885 13901 10937 14023
rect 11967 13990 12019 14013
rect 11695 13977 11747 13989
rect 11695 13943 11703 13977
rect 11737 13943 11747 13977
rect 10885 13867 10895 13901
rect 10929 13867 10937 13901
rect 10885 13855 10937 13867
rect 11000 13927 11052 13939
rect 11000 13893 11008 13927
rect 11042 13893 11052 13927
rect 11000 13855 11052 13893
rect 11082 13911 11149 13939
rect 11082 13877 11092 13911
rect 11126 13877 11149 13911
rect 11082 13855 11149 13877
rect 11179 13927 11289 13939
rect 11179 13893 11189 13927
rect 11223 13893 11289 13927
rect 11179 13855 11289 13893
rect 11319 13903 11388 13939
rect 11319 13869 11343 13903
rect 11377 13869 11388 13903
rect 11319 13855 11388 13869
rect 11418 13909 11480 13939
rect 11418 13875 11436 13909
rect 11470 13875 11480 13909
rect 11418 13855 11480 13875
rect 11510 13901 11562 13939
rect 11510 13867 11520 13901
rect 11554 13867 11562 13901
rect 11510 13855 11562 13867
rect 11695 13909 11747 13943
rect 11695 13875 11703 13909
rect 11737 13875 11747 13909
rect 11695 13861 11747 13875
rect 11777 13925 11831 13989
rect 11777 13891 11787 13925
rect 11821 13891 11831 13925
rect 11777 13861 11831 13891
rect 11861 13977 11913 13989
rect 11861 13943 11871 13977
rect 11905 13943 11913 13977
rect 11861 13909 11913 13943
rect 11861 13875 11871 13909
rect 11905 13875 11913 13909
rect 11861 13861 11913 13875
rect 11967 13956 11975 13990
rect 12009 13956 12019 13990
rect 11967 13909 12019 13956
rect 11967 13875 11975 13909
rect 12009 13875 12019 13909
rect 11967 13855 12019 13875
rect 12049 13977 12107 14013
rect 12049 13943 12061 13977
rect 12095 13943 12107 13977
rect 12049 13909 12107 13943
rect 12049 13875 12061 13909
rect 12095 13875 12107 13909
rect 12049 13855 12107 13875
rect 12137 13977 12189 14013
rect 12137 13943 12147 13977
rect 12181 13943 12189 13977
rect 12137 13909 12189 13943
rect 12137 13875 12147 13909
rect 12181 13875 12189 13909
rect 12137 13855 12189 13875
rect 12260 13925 12313 14055
rect 12260 13891 12268 13925
rect 12302 13891 12313 13925
rect 12260 13855 12313 13891
rect 12343 14031 12399 14055
rect 12343 13997 12354 14031
rect 12388 13997 12399 14031
rect 12343 13945 12399 13997
rect 12343 13911 12354 13945
rect 12388 13911 12399 13945
rect 12343 13855 12399 13911
rect 12429 13925 12485 14055
rect 12429 13891 12440 13925
rect 12474 13891 12485 13925
rect 12429 13855 12485 13891
rect 12515 14031 12571 14055
rect 12515 13997 12526 14031
rect 12560 13997 12571 14031
rect 12515 13945 12571 13997
rect 12515 13911 12526 13945
rect 12560 13911 12571 13945
rect 12515 13855 12571 13911
rect 12601 13925 12657 14055
rect 12601 13891 12612 13925
rect 12646 13891 12657 13925
rect 12601 13855 12657 13891
rect 12687 14031 12743 14055
rect 12687 13997 12698 14031
rect 12732 13997 12743 14031
rect 12687 13945 12743 13997
rect 12687 13911 12698 13945
rect 12732 13911 12743 13945
rect 12687 13855 12743 13911
rect 12773 13925 12829 14055
rect 12773 13891 12784 13925
rect 12818 13891 12829 13925
rect 12773 13855 12829 13891
rect 12859 14031 12915 14055
rect 12859 13997 12870 14031
rect 12904 13997 12915 14031
rect 12859 13945 12915 13997
rect 12859 13911 12870 13945
rect 12904 13911 12915 13945
rect 12859 13855 12915 13911
rect 12945 13925 13000 14055
rect 12945 13891 12955 13925
rect 12989 13891 13000 13925
rect 12945 13855 13000 13891
rect 13030 14031 13086 14055
rect 13030 13997 13041 14031
rect 13075 13997 13086 14031
rect 13030 13945 13086 13997
rect 13030 13911 13041 13945
rect 13075 13911 13086 13945
rect 13030 13855 13086 13911
rect 13116 13925 13172 14055
rect 13116 13891 13127 13925
rect 13161 13891 13172 13925
rect 13116 13855 13172 13891
rect 13202 14031 13258 14055
rect 13202 13997 13213 14031
rect 13247 13997 13258 14031
rect 13202 13945 13258 13997
rect 13202 13911 13213 13945
rect 13247 13911 13258 13945
rect 13202 13855 13258 13911
rect 13288 13925 13344 14055
rect 13288 13891 13299 13925
rect 13333 13891 13344 13925
rect 13288 13855 13344 13891
rect 13374 14031 13430 14055
rect 13374 13997 13385 14031
rect 13419 13997 13430 14031
rect 13374 13945 13430 13997
rect 13374 13911 13385 13945
rect 13419 13911 13430 13945
rect 13374 13855 13430 13911
rect 13460 13925 13516 14055
rect 13460 13891 13471 13925
rect 13505 13891 13516 13925
rect 13460 13855 13516 13891
rect 13546 14031 13602 14055
rect 13546 13997 13557 14031
rect 13591 13997 13602 14031
rect 13546 13945 13602 13997
rect 13546 13911 13557 13945
rect 13591 13911 13602 13945
rect 13546 13855 13602 13911
rect 13632 13969 13688 14055
rect 13632 13935 13643 13969
rect 13677 13935 13688 13969
rect 13632 13901 13688 13935
rect 13632 13867 13643 13901
rect 13677 13867 13688 13901
rect 13632 13855 13688 13867
rect 13718 13985 13774 14055
rect 13718 13951 13729 13985
rect 13763 13951 13774 13985
rect 13718 13917 13774 13951
rect 13718 13883 13729 13917
rect 13763 13883 13774 13917
rect 13718 13855 13774 13883
rect 13804 13969 13860 14055
rect 13804 13935 13815 13969
rect 13849 13935 13860 13969
rect 13804 13901 13860 13935
rect 13804 13867 13815 13901
rect 13849 13867 13860 13901
rect 13804 13855 13860 13867
rect 13890 13977 13946 14055
rect 13890 13943 13901 13977
rect 13935 13943 13946 13977
rect 13890 13909 13946 13943
rect 13890 13875 13901 13909
rect 13935 13875 13946 13909
rect 13890 13855 13946 13875
rect 13976 13969 14029 14055
rect 13976 13935 13987 13969
rect 14021 13935 14029 13969
rect 14798 13939 14848 14055
rect 13976 13901 14029 13935
rect 13976 13867 13987 13901
rect 14021 13867 14029 13901
rect 13976 13855 14029 13867
rect 14289 13927 14341 13939
rect 14289 13893 14297 13927
rect 14331 13893 14341 13927
rect 14289 13855 14341 13893
rect 14371 13901 14425 13939
rect 14371 13867 14381 13901
rect 14415 13867 14425 13901
rect 14371 13855 14425 13867
rect 14525 13927 14577 13939
rect 14525 13893 14535 13927
rect 14569 13893 14577 13927
rect 14525 13855 14577 13893
rect 14631 13927 14683 13939
rect 14631 13893 14639 13927
rect 14673 13893 14683 13927
rect 14631 13855 14683 13893
rect 14783 13901 14848 13939
rect 14783 13867 14798 13901
rect 14832 13867 14848 13901
rect 14783 13855 14848 13867
rect 14878 13927 14930 14055
rect 14878 13893 14888 13927
rect 14922 13893 14930 13927
rect 14878 13855 14930 13893
rect 15187 14037 15239 14055
rect 15187 14003 15195 14037
rect 15229 14003 15239 14037
rect 15187 13969 15239 14003
rect 15187 13935 15195 13969
rect 15229 13935 15239 13969
rect 15187 13901 15239 13935
rect 15187 13867 15195 13901
rect 15229 13867 15239 13901
rect 15187 13855 15239 13867
rect 15269 14037 15321 14055
rect 15269 14003 15279 14037
rect 15313 14003 15321 14037
rect 15269 13978 15321 14003
rect 16015 13990 16067 14013
rect 15269 13969 15348 13978
rect 15269 13935 15279 13969
rect 15313 13935 15348 13969
rect 15269 13901 15348 13935
rect 15269 13867 15279 13901
rect 15313 13894 15348 13901
rect 15378 13894 15451 13978
rect 15481 13961 15665 13978
rect 15481 13927 15515 13961
rect 15549 13927 15590 13961
rect 15624 13927 15665 13961
rect 15481 13894 15665 13927
rect 15695 13894 15737 13978
rect 15767 13961 15833 13978
rect 15767 13927 15787 13961
rect 15821 13927 15833 13961
rect 15767 13894 15833 13927
rect 15863 13961 15919 13978
rect 15863 13927 15873 13961
rect 15907 13927 15919 13961
rect 15863 13894 15919 13927
rect 16015 13956 16023 13990
rect 16057 13956 16067 13990
rect 16015 13909 16067 13956
rect 15313 13867 15321 13894
rect 16015 13875 16023 13909
rect 16057 13875 16067 13909
rect 15269 13855 15321 13867
rect 16015 13855 16067 13875
rect 16097 13977 16155 14013
rect 16097 13943 16109 13977
rect 16143 13943 16155 13977
rect 16097 13909 16155 13943
rect 16097 13875 16109 13909
rect 16143 13875 16155 13909
rect 16097 13855 16155 13875
rect 16185 13977 16237 14013
rect 16185 13943 16195 13977
rect 16229 13943 16237 13977
rect 16185 13909 16237 13943
rect 16185 13875 16195 13909
rect 16229 13875 16237 13909
rect 16185 13855 16237 13875
rect 16291 13990 16343 14013
rect 16291 13956 16299 13990
rect 16333 13956 16343 13990
rect 16291 13909 16343 13956
rect 16291 13875 16299 13909
rect 16333 13875 16343 13909
rect 16291 13855 16343 13875
rect 16373 13977 16431 14013
rect 16373 13943 16385 13977
rect 16419 13943 16431 13977
rect 16373 13909 16431 13943
rect 16373 13875 16385 13909
rect 16419 13875 16431 13909
rect 16373 13855 16431 13875
rect 16461 13977 16513 14013
rect 16461 13943 16471 13977
rect 16505 13943 16513 13977
rect 16461 13909 16513 13943
rect 16461 13875 16471 13909
rect 16505 13875 16513 13909
rect 16461 13855 16513 13875
rect 16659 13901 16711 14029
rect 16659 13867 16667 13901
rect 16701 13867 16711 13901
rect 16659 13855 16711 13867
rect 17657 13901 17709 14029
rect 17657 13867 17667 13901
rect 17701 13867 17709 13901
rect 17657 13855 17709 13867
rect 17763 13901 17815 14029
rect 17763 13867 17771 13901
rect 17805 13867 17815 13901
rect 17763 13855 17815 13867
rect 18761 13901 18813 14029
rect 18761 13867 18771 13901
rect 18805 13867 18813 13901
rect 18761 13855 18813 13867
rect 18867 13901 18919 14029
rect 18867 13867 18875 13901
rect 18909 13867 18919 13901
rect 18867 13855 18919 13867
rect 19865 13901 19917 14029
rect 19865 13867 19875 13901
rect 19909 13867 19917 13901
rect 19865 13855 19917 13867
rect 19971 13996 20023 14029
rect 19971 13962 19979 13996
rect 20013 13962 20023 13996
rect 19971 13901 20023 13962
rect 19971 13867 19979 13901
rect 20013 13867 20023 13901
rect 19971 13855 20023 13867
rect 20141 13996 20193 14029
rect 20141 13962 20151 13996
rect 20185 13962 20193 13996
rect 20141 13901 20193 13962
rect 20141 13867 20151 13901
rect 20185 13867 20193 13901
rect 20141 13855 20193 13867
rect 4975 13749 5027 13761
rect 4975 13715 4983 13749
rect 5017 13715 5027 13749
rect 4975 13654 5027 13715
rect 4975 13620 4983 13654
rect 5017 13620 5027 13654
rect 4975 13587 5027 13620
rect 5145 13749 5197 13761
rect 5145 13715 5155 13749
rect 5189 13715 5197 13749
rect 5145 13654 5197 13715
rect 5145 13620 5155 13654
rect 5189 13620 5197 13654
rect 5145 13587 5197 13620
rect 5435 13749 5487 13761
rect 5435 13715 5443 13749
rect 5477 13715 5487 13749
rect 5435 13647 5487 13715
rect 5435 13613 5443 13647
rect 5477 13613 5487 13647
rect 5435 13587 5487 13613
rect 6065 13749 6117 13761
rect 6065 13715 6075 13749
rect 6109 13715 6117 13749
rect 6065 13647 6117 13715
rect 6065 13613 6075 13647
rect 6109 13613 6117 13647
rect 6065 13587 6117 13613
rect 6171 13749 6223 13761
rect 6171 13715 6179 13749
rect 6213 13715 6223 13749
rect 6171 13587 6223 13715
rect 7169 13749 7221 13761
rect 7169 13715 7179 13749
rect 7213 13715 7221 13749
rect 7459 13749 7511 13761
rect 7169 13587 7221 13715
rect 7459 13715 7467 13749
rect 7501 13715 7511 13749
rect 7459 13587 7511 13715
rect 8457 13749 8509 13761
rect 8457 13715 8467 13749
rect 8501 13715 8509 13749
rect 8457 13587 8509 13715
rect 8563 13749 8615 13761
rect 8563 13715 8571 13749
rect 8605 13715 8615 13749
rect 8563 13587 8615 13715
rect 9561 13749 9613 13761
rect 9561 13715 9571 13749
rect 9605 13715 9613 13749
rect 9561 13587 9613 13715
rect 9667 13741 9719 13761
rect 9667 13707 9675 13741
rect 9709 13707 9719 13741
rect 9667 13673 9719 13707
rect 9667 13639 9675 13673
rect 9709 13639 9719 13673
rect 9667 13603 9719 13639
rect 9749 13741 9807 13761
rect 9749 13707 9761 13741
rect 9795 13707 9807 13741
rect 9749 13673 9807 13707
rect 9749 13639 9761 13673
rect 9795 13639 9807 13673
rect 9749 13603 9807 13639
rect 9837 13741 9889 13761
rect 9837 13707 9847 13741
rect 9881 13707 9889 13741
rect 9837 13660 9889 13707
rect 9837 13626 9847 13660
rect 9881 13626 9889 13660
rect 9837 13603 9889 13626
rect 9960 13725 10013 13761
rect 9960 13691 9968 13725
rect 10002 13691 10013 13725
rect 9960 13561 10013 13691
rect 10043 13705 10099 13761
rect 10043 13671 10054 13705
rect 10088 13671 10099 13705
rect 10043 13619 10099 13671
rect 10043 13585 10054 13619
rect 10088 13585 10099 13619
rect 10043 13561 10099 13585
rect 10129 13725 10185 13761
rect 10129 13691 10140 13725
rect 10174 13691 10185 13725
rect 10129 13561 10185 13691
rect 10215 13705 10271 13761
rect 10215 13671 10226 13705
rect 10260 13671 10271 13705
rect 10215 13619 10271 13671
rect 10215 13585 10226 13619
rect 10260 13585 10271 13619
rect 10215 13561 10271 13585
rect 10301 13725 10357 13761
rect 10301 13691 10312 13725
rect 10346 13691 10357 13725
rect 10301 13561 10357 13691
rect 10387 13705 10443 13761
rect 10387 13671 10398 13705
rect 10432 13671 10443 13705
rect 10387 13619 10443 13671
rect 10387 13585 10398 13619
rect 10432 13585 10443 13619
rect 10387 13561 10443 13585
rect 10473 13725 10529 13761
rect 10473 13691 10484 13725
rect 10518 13691 10529 13725
rect 10473 13561 10529 13691
rect 10559 13705 10615 13761
rect 10559 13671 10570 13705
rect 10604 13671 10615 13705
rect 10559 13619 10615 13671
rect 10559 13585 10570 13619
rect 10604 13585 10615 13619
rect 10559 13561 10615 13585
rect 10645 13725 10700 13761
rect 10645 13691 10655 13725
rect 10689 13691 10700 13725
rect 10645 13561 10700 13691
rect 10730 13705 10786 13761
rect 10730 13671 10741 13705
rect 10775 13671 10786 13705
rect 10730 13619 10786 13671
rect 10730 13585 10741 13619
rect 10775 13585 10786 13619
rect 10730 13561 10786 13585
rect 10816 13725 10872 13761
rect 10816 13691 10827 13725
rect 10861 13691 10872 13725
rect 10816 13561 10872 13691
rect 10902 13705 10958 13761
rect 10902 13671 10913 13705
rect 10947 13671 10958 13705
rect 10902 13619 10958 13671
rect 10902 13585 10913 13619
rect 10947 13585 10958 13619
rect 10902 13561 10958 13585
rect 10988 13725 11044 13761
rect 10988 13691 10999 13725
rect 11033 13691 11044 13725
rect 10988 13561 11044 13691
rect 11074 13705 11130 13761
rect 11074 13671 11085 13705
rect 11119 13671 11130 13705
rect 11074 13619 11130 13671
rect 11074 13585 11085 13619
rect 11119 13585 11130 13619
rect 11074 13561 11130 13585
rect 11160 13725 11216 13761
rect 11160 13691 11171 13725
rect 11205 13691 11216 13725
rect 11160 13561 11216 13691
rect 11246 13705 11302 13761
rect 11246 13671 11257 13705
rect 11291 13671 11302 13705
rect 11246 13619 11302 13671
rect 11246 13585 11257 13619
rect 11291 13585 11302 13619
rect 11246 13561 11302 13585
rect 11332 13749 11388 13761
rect 11332 13715 11343 13749
rect 11377 13715 11388 13749
rect 11332 13681 11388 13715
rect 11332 13647 11343 13681
rect 11377 13647 11388 13681
rect 11332 13561 11388 13647
rect 11418 13733 11474 13761
rect 11418 13699 11429 13733
rect 11463 13699 11474 13733
rect 11418 13665 11474 13699
rect 11418 13631 11429 13665
rect 11463 13631 11474 13665
rect 11418 13561 11474 13631
rect 11504 13749 11560 13761
rect 11504 13715 11515 13749
rect 11549 13715 11560 13749
rect 11504 13681 11560 13715
rect 11504 13647 11515 13681
rect 11549 13647 11560 13681
rect 11504 13561 11560 13647
rect 11590 13741 11646 13761
rect 11590 13707 11601 13741
rect 11635 13707 11646 13741
rect 11590 13673 11646 13707
rect 11590 13639 11601 13673
rect 11635 13639 11646 13673
rect 11590 13561 11646 13639
rect 11676 13749 11729 13761
rect 11676 13715 11687 13749
rect 11721 13715 11729 13749
rect 11676 13681 11729 13715
rect 11676 13647 11687 13681
rect 11721 13647 11729 13681
rect 11676 13561 11729 13647
rect 11875 13749 11927 13761
rect 11875 13715 11883 13749
rect 11917 13715 11927 13749
rect 11875 13647 11927 13715
rect 11875 13613 11883 13647
rect 11917 13613 11927 13647
rect 11875 13587 11927 13613
rect 12321 13749 12373 13761
rect 12321 13715 12331 13749
rect 12365 13715 12373 13749
rect 12321 13647 12373 13715
rect 12321 13613 12331 13647
rect 12365 13613 12373 13647
rect 12321 13587 12373 13613
rect 12519 13741 12571 13761
rect 12519 13707 12527 13741
rect 12561 13707 12571 13741
rect 12519 13660 12571 13707
rect 12519 13626 12527 13660
rect 12561 13626 12571 13660
rect 12519 13603 12571 13626
rect 12601 13741 12659 13761
rect 12601 13707 12613 13741
rect 12647 13707 12659 13741
rect 12601 13673 12659 13707
rect 12601 13639 12613 13673
rect 12647 13639 12659 13673
rect 12601 13603 12659 13639
rect 12689 13741 12741 13761
rect 12689 13707 12699 13741
rect 12733 13707 12741 13741
rect 12689 13673 12741 13707
rect 12689 13639 12699 13673
rect 12733 13639 12741 13673
rect 12689 13603 12741 13639
rect 12887 13713 12939 13761
rect 12887 13679 12895 13713
rect 12929 13679 12939 13713
rect 12887 13645 12939 13679
rect 12887 13611 12895 13645
rect 12929 13611 12939 13645
rect 12887 13561 12939 13611
rect 12969 13749 13035 13761
rect 12969 13715 12979 13749
rect 13013 13715 13035 13749
rect 12969 13681 13035 13715
rect 12969 13647 12979 13681
rect 13013 13647 13035 13681
rect 13100 13749 13154 13761
rect 13100 13715 13108 13749
rect 13142 13715 13154 13749
rect 13100 13677 13154 13715
rect 13184 13723 13238 13761
rect 13184 13689 13194 13723
rect 13228 13689 13238 13723
rect 13184 13677 13238 13689
rect 13268 13749 13346 13761
rect 13268 13715 13278 13749
rect 13312 13715 13346 13749
rect 13268 13677 13346 13715
rect 13376 13677 13430 13761
rect 13460 13748 13516 13761
rect 13460 13714 13470 13748
rect 13504 13714 13516 13748
rect 13460 13677 13516 13714
rect 13546 13741 13615 13761
rect 13546 13707 13567 13741
rect 13601 13707 13615 13741
rect 13546 13677 13615 13707
rect 12969 13633 13035 13647
rect 12969 13561 13019 13633
rect 13561 13593 13615 13677
rect 13645 13749 13697 13761
rect 13645 13715 13655 13749
rect 13689 13715 13697 13749
rect 13645 13593 13697 13715
rect 13760 13723 13812 13761
rect 13760 13689 13768 13723
rect 13802 13689 13812 13723
rect 13760 13677 13812 13689
rect 13842 13739 13909 13761
rect 13842 13705 13852 13739
rect 13886 13705 13909 13739
rect 13842 13677 13909 13705
rect 13939 13723 14049 13761
rect 13939 13689 13949 13723
rect 13983 13689 14049 13723
rect 13939 13677 14049 13689
rect 14079 13747 14148 13761
rect 14079 13713 14103 13747
rect 14137 13713 14148 13747
rect 14079 13677 14148 13713
rect 14178 13741 14240 13761
rect 14178 13707 14196 13741
rect 14230 13707 14240 13741
rect 14178 13677 14240 13707
rect 14270 13749 14322 13761
rect 14270 13715 14280 13749
rect 14314 13715 14322 13749
rect 14270 13677 14322 13715
rect 14455 13741 14507 13755
rect 14455 13707 14463 13741
rect 14497 13707 14507 13741
rect 14455 13673 14507 13707
rect 14455 13639 14463 13673
rect 14497 13639 14507 13673
rect 14455 13627 14507 13639
rect 14537 13725 14591 13755
rect 14537 13691 14547 13725
rect 14581 13691 14591 13725
rect 14537 13627 14591 13691
rect 14621 13741 14673 13755
rect 14621 13707 14631 13741
rect 14665 13707 14673 13741
rect 14621 13673 14673 13707
rect 14621 13639 14631 13673
rect 14665 13639 14673 13673
rect 14621 13627 14673 13639
rect 14727 13749 14780 13761
rect 14727 13715 14735 13749
rect 14769 13715 14780 13749
rect 14727 13681 14780 13715
rect 14727 13647 14735 13681
rect 14769 13647 14780 13681
rect 14727 13561 14780 13647
rect 14810 13741 14866 13761
rect 14810 13707 14821 13741
rect 14855 13707 14866 13741
rect 14810 13673 14866 13707
rect 14810 13639 14821 13673
rect 14855 13639 14866 13673
rect 14810 13561 14866 13639
rect 14896 13749 14952 13761
rect 14896 13715 14907 13749
rect 14941 13715 14952 13749
rect 14896 13681 14952 13715
rect 14896 13647 14907 13681
rect 14941 13647 14952 13681
rect 14896 13561 14952 13647
rect 14982 13733 15038 13761
rect 14982 13699 14993 13733
rect 15027 13699 15038 13733
rect 14982 13665 15038 13699
rect 14982 13631 14993 13665
rect 15027 13631 15038 13665
rect 14982 13561 15038 13631
rect 15068 13749 15124 13761
rect 15068 13715 15079 13749
rect 15113 13715 15124 13749
rect 15068 13681 15124 13715
rect 15068 13647 15079 13681
rect 15113 13647 15124 13681
rect 15068 13561 15124 13647
rect 15154 13705 15210 13761
rect 15154 13671 15165 13705
rect 15199 13671 15210 13705
rect 15154 13619 15210 13671
rect 15154 13585 15165 13619
rect 15199 13585 15210 13619
rect 15154 13561 15210 13585
rect 15240 13725 15296 13761
rect 15240 13691 15251 13725
rect 15285 13691 15296 13725
rect 15240 13561 15296 13691
rect 15326 13705 15382 13761
rect 15326 13671 15337 13705
rect 15371 13671 15382 13705
rect 15326 13619 15382 13671
rect 15326 13585 15337 13619
rect 15371 13585 15382 13619
rect 15326 13561 15382 13585
rect 15412 13725 15468 13761
rect 15412 13691 15423 13725
rect 15457 13691 15468 13725
rect 15412 13561 15468 13691
rect 15498 13705 15554 13761
rect 15498 13671 15509 13705
rect 15543 13671 15554 13705
rect 15498 13619 15554 13671
rect 15498 13585 15509 13619
rect 15543 13585 15554 13619
rect 15498 13561 15554 13585
rect 15584 13725 15640 13761
rect 15584 13691 15595 13725
rect 15629 13691 15640 13725
rect 15584 13561 15640 13691
rect 15670 13705 15726 13761
rect 15670 13671 15681 13705
rect 15715 13671 15726 13705
rect 15670 13619 15726 13671
rect 15670 13585 15681 13619
rect 15715 13585 15726 13619
rect 15670 13561 15726 13585
rect 15756 13725 15811 13761
rect 15756 13691 15767 13725
rect 15801 13691 15811 13725
rect 15756 13561 15811 13691
rect 15841 13705 15897 13761
rect 15841 13671 15852 13705
rect 15886 13671 15897 13705
rect 15841 13619 15897 13671
rect 15841 13585 15852 13619
rect 15886 13585 15897 13619
rect 15841 13561 15897 13585
rect 15927 13725 15983 13761
rect 15927 13691 15938 13725
rect 15972 13691 15983 13725
rect 15927 13561 15983 13691
rect 16013 13705 16069 13761
rect 16013 13671 16024 13705
rect 16058 13671 16069 13705
rect 16013 13619 16069 13671
rect 16013 13585 16024 13619
rect 16058 13585 16069 13619
rect 16013 13561 16069 13585
rect 16099 13725 16155 13761
rect 16099 13691 16110 13725
rect 16144 13691 16155 13725
rect 16099 13561 16155 13691
rect 16185 13705 16241 13761
rect 16185 13671 16196 13705
rect 16230 13671 16241 13705
rect 16185 13619 16241 13671
rect 16185 13585 16196 13619
rect 16230 13585 16241 13619
rect 16185 13561 16241 13585
rect 16271 13725 16327 13761
rect 16271 13691 16282 13725
rect 16316 13691 16327 13725
rect 16271 13561 16327 13691
rect 16357 13705 16413 13761
rect 16357 13671 16368 13705
rect 16402 13671 16413 13705
rect 16357 13619 16413 13671
rect 16357 13585 16368 13619
rect 16402 13585 16413 13619
rect 16357 13561 16413 13585
rect 16443 13725 16496 13761
rect 16443 13691 16454 13725
rect 16488 13691 16496 13725
rect 16443 13561 16496 13691
rect 16567 13749 16619 13761
rect 16567 13715 16575 13749
rect 16609 13715 16619 13749
rect 16567 13681 16619 13715
rect 16567 13647 16575 13681
rect 16609 13647 16619 13681
rect 16567 13613 16619 13647
rect 16567 13579 16575 13613
rect 16609 13579 16619 13613
rect 16567 13561 16619 13579
rect 16649 13749 16701 13761
rect 16649 13715 16659 13749
rect 16693 13722 16701 13749
rect 17763 13749 17815 13761
rect 16693 13715 16728 13722
rect 16649 13681 16728 13715
rect 16649 13647 16659 13681
rect 16693 13647 16728 13681
rect 16649 13638 16728 13647
rect 16758 13638 16831 13722
rect 16861 13689 17045 13722
rect 16861 13655 16895 13689
rect 16929 13655 16970 13689
rect 17004 13655 17045 13689
rect 16861 13638 17045 13655
rect 17075 13638 17117 13722
rect 17147 13689 17213 13722
rect 17147 13655 17167 13689
rect 17201 13655 17213 13689
rect 17147 13638 17213 13655
rect 17243 13689 17299 13722
rect 17243 13655 17253 13689
rect 17287 13655 17299 13689
rect 17243 13638 17299 13655
rect 16649 13613 16701 13638
rect 16649 13579 16659 13613
rect 16693 13579 16701 13613
rect 16649 13561 16701 13579
rect 17763 13715 17771 13749
rect 17805 13715 17815 13749
rect 17763 13587 17815 13715
rect 18761 13749 18813 13761
rect 18761 13715 18771 13749
rect 18805 13715 18813 13749
rect 18761 13587 18813 13715
rect 18867 13749 18919 13761
rect 18867 13715 18875 13749
rect 18909 13715 18919 13749
rect 18867 13587 18919 13715
rect 19865 13749 19917 13761
rect 19865 13715 19875 13749
rect 19909 13715 19917 13749
rect 19865 13587 19917 13715
rect 19971 13749 20023 13761
rect 19971 13715 19979 13749
rect 20013 13715 20023 13749
rect 19971 13654 20023 13715
rect 19971 13620 19979 13654
rect 20013 13620 20023 13654
rect 19971 13587 20023 13620
rect 20141 13749 20193 13761
rect 20141 13715 20151 13749
rect 20185 13715 20193 13749
rect 20141 13654 20193 13715
rect 20141 13620 20151 13654
rect 20185 13620 20193 13654
rect 20141 13587 20193 13620
rect 4975 12908 5027 12941
rect 4975 12874 4983 12908
rect 5017 12874 5027 12908
rect 4975 12813 5027 12874
rect 4975 12779 4983 12813
rect 5017 12779 5027 12813
rect 4975 12767 5027 12779
rect 5145 12908 5197 12941
rect 5145 12874 5155 12908
rect 5189 12874 5197 12908
rect 5145 12813 5197 12874
rect 5145 12779 5155 12813
rect 5189 12779 5197 12813
rect 5145 12767 5197 12779
rect 5251 12915 5303 12941
rect 5251 12881 5259 12915
rect 5293 12881 5303 12915
rect 5251 12813 5303 12881
rect 5251 12779 5259 12813
rect 5293 12779 5303 12813
rect 5251 12767 5303 12779
rect 5697 12915 5749 12941
rect 5697 12881 5707 12915
rect 5741 12881 5749 12915
rect 5697 12813 5749 12881
rect 5697 12779 5707 12813
rect 5741 12779 5749 12813
rect 5697 12767 5749 12779
rect 5803 12813 5855 12941
rect 5803 12779 5811 12813
rect 5845 12779 5855 12813
rect 5803 12767 5855 12779
rect 6801 12813 6853 12941
rect 6801 12779 6811 12813
rect 6845 12779 6853 12813
rect 6801 12767 6853 12779
rect 6907 12813 6959 12941
rect 6907 12779 6915 12813
rect 6949 12779 6959 12813
rect 6907 12767 6959 12779
rect 7905 12813 7957 12941
rect 7905 12779 7915 12813
rect 7949 12779 7957 12813
rect 7905 12767 7957 12779
rect 8011 12813 8063 12941
rect 8011 12779 8019 12813
rect 8053 12779 8063 12813
rect 8011 12767 8063 12779
rect 9009 12813 9061 12941
rect 9646 12851 9696 12967
rect 9009 12779 9019 12813
rect 9053 12779 9061 12813
rect 9009 12767 9061 12779
rect 9137 12839 9189 12851
rect 9137 12805 9145 12839
rect 9179 12805 9189 12839
rect 9137 12767 9189 12805
rect 9219 12813 9273 12851
rect 9219 12779 9229 12813
rect 9263 12779 9273 12813
rect 9219 12767 9273 12779
rect 9373 12839 9425 12851
rect 9373 12805 9383 12839
rect 9417 12805 9425 12839
rect 9373 12767 9425 12805
rect 9479 12839 9531 12851
rect 9479 12805 9487 12839
rect 9521 12805 9531 12839
rect 9479 12767 9531 12805
rect 9631 12813 9696 12851
rect 9631 12779 9646 12813
rect 9680 12779 9696 12813
rect 9631 12767 9696 12779
rect 9726 12839 9778 12967
rect 9726 12805 9736 12839
rect 9770 12805 9778 12839
rect 9726 12767 9778 12805
rect 10035 12915 10087 12941
rect 10035 12881 10043 12915
rect 10077 12881 10087 12915
rect 10035 12813 10087 12881
rect 10035 12779 10043 12813
rect 10077 12779 10087 12813
rect 10035 12767 10087 12779
rect 10297 12915 10349 12941
rect 10297 12881 10307 12915
rect 10341 12881 10349 12915
rect 10297 12813 10349 12881
rect 10297 12779 10307 12813
rect 10341 12779 10349 12813
rect 10297 12767 10349 12779
rect 10403 12917 10455 12967
rect 10403 12883 10411 12917
rect 10445 12883 10455 12917
rect 10403 12849 10455 12883
rect 10403 12815 10411 12849
rect 10445 12815 10455 12849
rect 10403 12767 10455 12815
rect 10485 12895 10535 12967
rect 10485 12881 10551 12895
rect 10485 12847 10495 12881
rect 10529 12847 10551 12881
rect 11077 12851 11131 12935
rect 10485 12813 10551 12847
rect 10485 12779 10495 12813
rect 10529 12779 10551 12813
rect 10485 12767 10551 12779
rect 10616 12813 10670 12851
rect 10616 12779 10624 12813
rect 10658 12779 10670 12813
rect 10616 12767 10670 12779
rect 10700 12839 10754 12851
rect 10700 12805 10710 12839
rect 10744 12805 10754 12839
rect 10700 12767 10754 12805
rect 10784 12813 10862 12851
rect 10784 12779 10794 12813
rect 10828 12779 10862 12813
rect 10784 12767 10862 12779
rect 10892 12767 10946 12851
rect 10976 12814 11032 12851
rect 10976 12780 10986 12814
rect 11020 12780 11032 12814
rect 10976 12767 11032 12780
rect 11062 12821 11131 12851
rect 11062 12787 11083 12821
rect 11117 12787 11131 12821
rect 11062 12767 11131 12787
rect 11161 12813 11213 12935
rect 11971 12889 12023 12901
rect 11971 12855 11979 12889
rect 12013 12855 12023 12889
rect 11161 12779 11171 12813
rect 11205 12779 11213 12813
rect 11161 12767 11213 12779
rect 11276 12839 11328 12851
rect 11276 12805 11284 12839
rect 11318 12805 11328 12839
rect 11276 12767 11328 12805
rect 11358 12823 11425 12851
rect 11358 12789 11368 12823
rect 11402 12789 11425 12823
rect 11358 12767 11425 12789
rect 11455 12839 11565 12851
rect 11455 12805 11465 12839
rect 11499 12805 11565 12839
rect 11455 12767 11565 12805
rect 11595 12815 11664 12851
rect 11595 12781 11619 12815
rect 11653 12781 11664 12815
rect 11595 12767 11664 12781
rect 11694 12821 11756 12851
rect 11694 12787 11712 12821
rect 11746 12787 11756 12821
rect 11694 12767 11756 12787
rect 11786 12813 11838 12851
rect 11786 12779 11796 12813
rect 11830 12779 11838 12813
rect 11786 12767 11838 12779
rect 11971 12821 12023 12855
rect 11971 12787 11979 12821
rect 12013 12787 12023 12821
rect 11971 12773 12023 12787
rect 12053 12837 12107 12901
rect 12053 12803 12063 12837
rect 12097 12803 12107 12837
rect 12053 12773 12107 12803
rect 12137 12889 12189 12901
rect 12137 12855 12147 12889
rect 12181 12855 12189 12889
rect 12137 12821 12189 12855
rect 12137 12787 12147 12821
rect 12181 12787 12189 12821
rect 12137 12773 12189 12787
rect 12243 12889 12295 12901
rect 12243 12855 12251 12889
rect 12285 12855 12295 12889
rect 12243 12821 12295 12855
rect 12243 12787 12251 12821
rect 12285 12787 12295 12821
rect 12243 12773 12295 12787
rect 12325 12837 12379 12901
rect 12325 12803 12335 12837
rect 12369 12803 12379 12837
rect 12325 12773 12379 12803
rect 12409 12889 12461 12901
rect 12409 12855 12419 12889
rect 12453 12855 12461 12889
rect 12409 12821 12461 12855
rect 12409 12787 12419 12821
rect 12453 12787 12461 12821
rect 12409 12773 12461 12787
rect 12594 12813 12646 12851
rect 12594 12779 12602 12813
rect 12636 12779 12646 12813
rect 12594 12767 12646 12779
rect 12676 12821 12738 12851
rect 12676 12787 12686 12821
rect 12720 12787 12738 12821
rect 12676 12767 12738 12787
rect 12768 12815 12837 12851
rect 12768 12781 12779 12815
rect 12813 12781 12837 12815
rect 12768 12767 12837 12781
rect 12867 12839 12977 12851
rect 12867 12805 12933 12839
rect 12967 12805 12977 12839
rect 12867 12767 12977 12805
rect 13007 12823 13074 12851
rect 13007 12789 13030 12823
rect 13064 12789 13074 12823
rect 13007 12767 13074 12789
rect 13104 12839 13156 12851
rect 13104 12805 13114 12839
rect 13148 12805 13156 12839
rect 13104 12767 13156 12805
rect 13219 12813 13271 12935
rect 13219 12779 13227 12813
rect 13261 12779 13271 12813
rect 13219 12767 13271 12779
rect 13301 12851 13355 12935
rect 13897 12895 13947 12967
rect 13881 12881 13947 12895
rect 13301 12821 13370 12851
rect 13301 12787 13315 12821
rect 13349 12787 13370 12821
rect 13301 12767 13370 12787
rect 13400 12814 13456 12851
rect 13400 12780 13412 12814
rect 13446 12780 13456 12814
rect 13400 12767 13456 12780
rect 13486 12767 13540 12851
rect 13570 12813 13648 12851
rect 13570 12779 13604 12813
rect 13638 12779 13648 12813
rect 13570 12767 13648 12779
rect 13678 12839 13732 12851
rect 13678 12805 13688 12839
rect 13722 12805 13732 12839
rect 13678 12767 13732 12805
rect 13762 12813 13816 12851
rect 13762 12779 13774 12813
rect 13808 12779 13816 12813
rect 13762 12767 13816 12779
rect 13881 12847 13903 12881
rect 13937 12847 13947 12881
rect 13881 12813 13947 12847
rect 13881 12779 13903 12813
rect 13937 12779 13947 12813
rect 13881 12767 13947 12779
rect 13977 12917 14029 12967
rect 13977 12883 13987 12917
rect 14021 12883 14029 12917
rect 13977 12849 14029 12883
rect 13977 12815 13987 12849
rect 14021 12815 14029 12849
rect 13977 12767 14029 12815
rect 14083 12949 14135 12967
rect 14083 12915 14091 12949
rect 14125 12915 14135 12949
rect 14083 12881 14135 12915
rect 14083 12847 14091 12881
rect 14125 12847 14135 12881
rect 14083 12813 14135 12847
rect 14083 12779 14091 12813
rect 14125 12779 14135 12813
rect 14083 12767 14135 12779
rect 14165 12949 14217 12967
rect 14165 12915 14175 12949
rect 14209 12915 14217 12949
rect 14165 12890 14217 12915
rect 14165 12881 14244 12890
rect 14165 12847 14175 12881
rect 14209 12847 14244 12881
rect 14165 12813 14244 12847
rect 14165 12779 14175 12813
rect 14209 12806 14244 12813
rect 14274 12806 14347 12890
rect 14377 12873 14561 12890
rect 14377 12839 14411 12873
rect 14445 12839 14486 12873
rect 14520 12839 14561 12873
rect 14377 12806 14561 12839
rect 14591 12806 14633 12890
rect 14663 12873 14729 12890
rect 14663 12839 14683 12873
rect 14717 12839 14729 12873
rect 14663 12806 14729 12839
rect 14759 12873 14815 12890
rect 14759 12839 14769 12873
rect 14803 12839 14815 12873
rect 14759 12806 14815 12839
rect 14209 12779 14217 12806
rect 15095 12917 15147 12967
rect 15095 12883 15103 12917
rect 15137 12883 15147 12917
rect 15095 12849 15147 12883
rect 15095 12815 15103 12849
rect 15137 12815 15147 12849
rect 14165 12767 14217 12779
rect 15095 12767 15147 12815
rect 15177 12895 15227 12967
rect 15177 12881 15243 12895
rect 15177 12847 15187 12881
rect 15221 12847 15243 12881
rect 15769 12851 15823 12935
rect 15177 12813 15243 12847
rect 15177 12779 15187 12813
rect 15221 12779 15243 12813
rect 15177 12767 15243 12779
rect 15308 12813 15362 12851
rect 15308 12779 15316 12813
rect 15350 12779 15362 12813
rect 15308 12767 15362 12779
rect 15392 12839 15446 12851
rect 15392 12805 15402 12839
rect 15436 12805 15446 12839
rect 15392 12767 15446 12805
rect 15476 12813 15554 12851
rect 15476 12779 15486 12813
rect 15520 12779 15554 12813
rect 15476 12767 15554 12779
rect 15584 12767 15638 12851
rect 15668 12814 15724 12851
rect 15668 12780 15678 12814
rect 15712 12780 15724 12814
rect 15668 12767 15724 12780
rect 15754 12821 15823 12851
rect 15754 12787 15775 12821
rect 15809 12787 15823 12821
rect 15754 12767 15823 12787
rect 15853 12813 15905 12935
rect 16663 12889 16715 12901
rect 16663 12855 16671 12889
rect 16705 12855 16715 12889
rect 15853 12779 15863 12813
rect 15897 12779 15905 12813
rect 15853 12767 15905 12779
rect 15968 12839 16020 12851
rect 15968 12805 15976 12839
rect 16010 12805 16020 12839
rect 15968 12767 16020 12805
rect 16050 12823 16117 12851
rect 16050 12789 16060 12823
rect 16094 12789 16117 12823
rect 16050 12767 16117 12789
rect 16147 12839 16257 12851
rect 16147 12805 16157 12839
rect 16191 12805 16257 12839
rect 16147 12767 16257 12805
rect 16287 12815 16356 12851
rect 16287 12781 16311 12815
rect 16345 12781 16356 12815
rect 16287 12767 16356 12781
rect 16386 12821 16448 12851
rect 16386 12787 16404 12821
rect 16438 12787 16448 12821
rect 16386 12767 16448 12787
rect 16478 12813 16530 12851
rect 16478 12779 16488 12813
rect 16522 12779 16530 12813
rect 16478 12767 16530 12779
rect 16663 12821 16715 12855
rect 16663 12787 16671 12821
rect 16705 12787 16715 12821
rect 16663 12773 16715 12787
rect 16745 12837 16799 12901
rect 16745 12803 16755 12837
rect 16789 12803 16799 12837
rect 16745 12773 16799 12803
rect 16829 12889 16881 12901
rect 16829 12855 16839 12889
rect 16873 12855 16881 12889
rect 16829 12821 16881 12855
rect 16829 12787 16839 12821
rect 16873 12787 16881 12821
rect 16829 12773 16881 12787
rect 16954 12839 17006 12967
rect 16954 12805 16962 12839
rect 16996 12805 17006 12839
rect 16954 12767 17006 12805
rect 17036 12851 17086 12967
rect 17036 12813 17101 12851
rect 17036 12779 17052 12813
rect 17086 12779 17101 12813
rect 17036 12767 17101 12779
rect 17201 12839 17253 12851
rect 17201 12805 17211 12839
rect 17245 12805 17253 12839
rect 17201 12767 17253 12805
rect 17307 12839 17359 12851
rect 17307 12805 17315 12839
rect 17349 12805 17359 12839
rect 17307 12767 17359 12805
rect 17459 12813 17513 12851
rect 17459 12779 17469 12813
rect 17503 12779 17513 12813
rect 17459 12767 17513 12779
rect 17543 12839 17595 12851
rect 17543 12805 17553 12839
rect 17587 12805 17595 12839
rect 17543 12767 17595 12805
rect 17763 12813 17815 12941
rect 17763 12779 17771 12813
rect 17805 12779 17815 12813
rect 17763 12767 17815 12779
rect 18761 12813 18813 12941
rect 18761 12779 18771 12813
rect 18805 12779 18813 12813
rect 18761 12767 18813 12779
rect 18867 12813 18919 12941
rect 18867 12779 18875 12813
rect 18909 12779 18919 12813
rect 18867 12767 18919 12779
rect 19865 12813 19917 12941
rect 19865 12779 19875 12813
rect 19909 12779 19917 12813
rect 19865 12767 19917 12779
rect 19971 12908 20023 12941
rect 19971 12874 19979 12908
rect 20013 12874 20023 12908
rect 19971 12813 20023 12874
rect 19971 12779 19979 12813
rect 20013 12779 20023 12813
rect 19971 12767 20023 12779
rect 20141 12908 20193 12941
rect 20141 12874 20151 12908
rect 20185 12874 20193 12908
rect 20141 12813 20193 12874
rect 20141 12779 20151 12813
rect 20185 12779 20193 12813
rect 20141 12767 20193 12779
rect 4975 12661 5027 12673
rect 4975 12627 4983 12661
rect 5017 12627 5027 12661
rect 4975 12566 5027 12627
rect 4975 12532 4983 12566
rect 5017 12532 5027 12566
rect 4975 12499 5027 12532
rect 5145 12661 5197 12673
rect 5145 12627 5155 12661
rect 5189 12627 5197 12661
rect 5145 12566 5197 12627
rect 5145 12532 5155 12566
rect 5189 12532 5197 12566
rect 5145 12499 5197 12532
rect 5619 12661 5671 12673
rect 5619 12627 5627 12661
rect 5661 12627 5671 12661
rect 5619 12499 5671 12627
rect 6617 12661 6669 12673
rect 6617 12627 6627 12661
rect 6661 12627 6669 12661
rect 6617 12499 6669 12627
rect 6724 12647 6784 12673
rect 6724 12613 6739 12647
rect 6773 12613 6784 12647
rect 6724 12579 6784 12613
rect 6724 12545 6739 12579
rect 6773 12545 6784 12579
rect 6724 12473 6784 12545
rect 6814 12653 6870 12673
rect 6814 12619 6825 12653
rect 6859 12619 6870 12653
rect 6814 12585 6870 12619
rect 6814 12551 6825 12585
rect 6859 12551 6870 12585
rect 6814 12517 6870 12551
rect 6814 12483 6825 12517
rect 6859 12483 6870 12517
rect 6814 12473 6870 12483
rect 6900 12661 6956 12673
rect 6900 12627 6911 12661
rect 6945 12627 6956 12661
rect 6900 12473 6956 12627
rect 6986 12626 7042 12673
rect 6986 12592 6997 12626
rect 7031 12592 7042 12626
rect 6986 12473 7042 12592
rect 7072 12661 7138 12673
rect 7072 12627 7093 12661
rect 7127 12627 7138 12661
rect 7072 12593 7138 12627
rect 7072 12559 7093 12593
rect 7127 12559 7138 12593
rect 7072 12473 7138 12559
rect 7168 12653 7221 12673
rect 7367 12661 7419 12673
rect 7168 12619 7179 12653
rect 7213 12619 7221 12653
rect 7168 12531 7221 12619
rect 7168 12497 7179 12531
rect 7213 12497 7221 12531
rect 7168 12473 7221 12497
rect 7367 12627 7375 12661
rect 7409 12627 7419 12661
rect 7367 12559 7419 12627
rect 7367 12525 7375 12559
rect 7409 12525 7419 12559
rect 7367 12499 7419 12525
rect 7629 12661 7681 12673
rect 7629 12627 7639 12661
rect 7673 12627 7681 12661
rect 7629 12559 7681 12627
rect 7629 12525 7639 12559
rect 7673 12525 7681 12559
rect 7629 12499 7681 12525
rect 7735 12661 7787 12673
rect 7735 12627 7743 12661
rect 7777 12627 7787 12661
rect 7735 12499 7787 12627
rect 8733 12661 8785 12673
rect 8733 12627 8743 12661
rect 8777 12627 8785 12661
rect 8733 12499 8785 12627
rect 8840 12647 8900 12673
rect 8840 12613 8855 12647
rect 8889 12613 8900 12647
rect 8840 12579 8900 12613
rect 8840 12545 8855 12579
rect 8889 12545 8900 12579
rect 8840 12473 8900 12545
rect 8930 12653 8986 12673
rect 8930 12619 8941 12653
rect 8975 12619 8986 12653
rect 8930 12585 8986 12619
rect 8930 12551 8941 12585
rect 8975 12551 8986 12585
rect 8930 12517 8986 12551
rect 8930 12483 8941 12517
rect 8975 12483 8986 12517
rect 8930 12473 8986 12483
rect 9016 12661 9072 12673
rect 9016 12627 9027 12661
rect 9061 12627 9072 12661
rect 9016 12473 9072 12627
rect 9102 12626 9158 12673
rect 9102 12592 9113 12626
rect 9147 12592 9158 12626
rect 9102 12473 9158 12592
rect 9188 12661 9254 12673
rect 9188 12627 9209 12661
rect 9243 12627 9254 12661
rect 9188 12593 9254 12627
rect 9188 12559 9209 12593
rect 9243 12559 9254 12593
rect 9188 12473 9254 12559
rect 9284 12653 9337 12673
rect 9284 12619 9295 12653
rect 9329 12619 9337 12653
rect 9284 12531 9337 12619
rect 9284 12497 9295 12531
rect 9329 12497 9337 12531
rect 9483 12661 9535 12673
rect 9483 12627 9491 12661
rect 9525 12627 9535 12661
rect 9483 12559 9535 12627
rect 9483 12525 9491 12559
rect 9525 12525 9535 12559
rect 9483 12499 9535 12525
rect 9745 12661 9797 12673
rect 9745 12627 9755 12661
rect 9789 12627 9797 12661
rect 9745 12559 9797 12627
rect 9745 12525 9755 12559
rect 9789 12525 9797 12559
rect 9745 12499 9797 12525
rect 9284 12473 9337 12497
rect 9944 12647 10004 12673
rect 9944 12613 9959 12647
rect 9993 12613 10004 12647
rect 9944 12579 10004 12613
rect 9944 12545 9959 12579
rect 9993 12545 10004 12579
rect 9944 12473 10004 12545
rect 10034 12653 10090 12673
rect 10034 12619 10045 12653
rect 10079 12619 10090 12653
rect 10034 12585 10090 12619
rect 10034 12551 10045 12585
rect 10079 12551 10090 12585
rect 10034 12517 10090 12551
rect 10034 12483 10045 12517
rect 10079 12483 10090 12517
rect 10034 12473 10090 12483
rect 10120 12661 10176 12673
rect 10120 12627 10131 12661
rect 10165 12627 10176 12661
rect 10120 12473 10176 12627
rect 10206 12626 10262 12673
rect 10206 12592 10217 12626
rect 10251 12592 10262 12626
rect 10206 12473 10262 12592
rect 10292 12661 10358 12673
rect 10292 12627 10313 12661
rect 10347 12627 10358 12661
rect 10292 12593 10358 12627
rect 10292 12559 10313 12593
rect 10347 12559 10358 12593
rect 10292 12473 10358 12559
rect 10388 12653 10441 12673
rect 10388 12619 10399 12653
rect 10433 12619 10441 12653
rect 10388 12531 10441 12619
rect 10388 12497 10399 12531
rect 10433 12497 10441 12531
rect 10388 12473 10441 12497
rect 10495 12661 10547 12673
rect 10495 12627 10503 12661
rect 10537 12627 10547 12661
rect 10495 12593 10547 12627
rect 10495 12559 10503 12593
rect 10537 12559 10547 12593
rect 10495 12525 10547 12559
rect 10495 12491 10503 12525
rect 10537 12491 10547 12525
rect 10495 12473 10547 12491
rect 10577 12661 10629 12673
rect 10577 12627 10587 12661
rect 10621 12634 10629 12661
rect 12055 12661 12107 12673
rect 12055 12634 12063 12661
rect 10621 12627 10656 12634
rect 10577 12593 10656 12627
rect 10577 12559 10587 12593
rect 10621 12559 10656 12593
rect 10577 12550 10656 12559
rect 10686 12550 10759 12634
rect 10789 12601 10973 12634
rect 10789 12567 10823 12601
rect 10857 12567 10898 12601
rect 10932 12567 10973 12601
rect 10789 12550 10973 12567
rect 11003 12550 11045 12634
rect 11075 12601 11141 12634
rect 11075 12567 11095 12601
rect 11129 12567 11141 12601
rect 11075 12550 11141 12567
rect 11171 12601 11227 12634
rect 11171 12567 11181 12601
rect 11215 12567 11227 12601
rect 11171 12550 11227 12567
rect 11457 12601 11513 12634
rect 11457 12567 11469 12601
rect 11503 12567 11513 12601
rect 11457 12550 11513 12567
rect 11543 12601 11609 12634
rect 11543 12567 11555 12601
rect 11589 12567 11609 12601
rect 11543 12550 11609 12567
rect 11639 12550 11681 12634
rect 11711 12601 11895 12634
rect 11711 12567 11752 12601
rect 11786 12567 11827 12601
rect 11861 12567 11895 12601
rect 11711 12550 11895 12567
rect 11925 12550 11998 12634
rect 12028 12627 12063 12634
rect 12097 12627 12107 12661
rect 12028 12593 12107 12627
rect 12028 12559 12063 12593
rect 12097 12559 12107 12593
rect 12028 12550 12107 12559
rect 10577 12525 10629 12550
rect 10577 12491 10587 12525
rect 10621 12491 10629 12525
rect 10577 12473 10629 12491
rect 12055 12525 12107 12550
rect 12055 12491 12063 12525
rect 12097 12491 12107 12525
rect 12055 12473 12107 12491
rect 12137 12661 12189 12673
rect 12137 12627 12147 12661
rect 12181 12627 12189 12661
rect 12137 12593 12189 12627
rect 12137 12559 12147 12593
rect 12181 12559 12189 12593
rect 12137 12525 12189 12559
rect 12137 12491 12147 12525
rect 12181 12491 12189 12525
rect 12137 12473 12189 12491
rect 12704 12647 12764 12673
rect 12704 12613 12719 12647
rect 12753 12613 12764 12647
rect 12704 12579 12764 12613
rect 12704 12545 12719 12579
rect 12753 12545 12764 12579
rect 12704 12473 12764 12545
rect 12794 12653 12850 12673
rect 12794 12619 12805 12653
rect 12839 12619 12850 12653
rect 12794 12585 12850 12619
rect 12794 12551 12805 12585
rect 12839 12551 12850 12585
rect 12794 12517 12850 12551
rect 12794 12483 12805 12517
rect 12839 12483 12850 12517
rect 12794 12473 12850 12483
rect 12880 12661 12936 12673
rect 12880 12627 12891 12661
rect 12925 12627 12936 12661
rect 12880 12473 12936 12627
rect 12966 12626 13022 12673
rect 12966 12592 12977 12626
rect 13011 12592 13022 12626
rect 12966 12473 13022 12592
rect 13052 12661 13118 12673
rect 13052 12627 13073 12661
rect 13107 12627 13118 12661
rect 13052 12593 13118 12627
rect 13052 12559 13073 12593
rect 13107 12559 13118 12593
rect 13052 12473 13118 12559
rect 13148 12653 13201 12673
rect 13148 12619 13159 12653
rect 13193 12619 13201 12653
rect 13148 12531 13201 12619
rect 13148 12497 13159 12531
rect 13193 12497 13201 12531
rect 13148 12473 13201 12497
rect 13255 12653 13308 12673
rect 13255 12619 13263 12653
rect 13297 12619 13308 12653
rect 13255 12531 13308 12619
rect 13255 12497 13263 12531
rect 13297 12497 13308 12531
rect 13255 12473 13308 12497
rect 13338 12661 13404 12673
rect 13338 12627 13349 12661
rect 13383 12627 13404 12661
rect 13338 12593 13404 12627
rect 13338 12559 13349 12593
rect 13383 12559 13404 12593
rect 13338 12473 13404 12559
rect 13434 12626 13490 12673
rect 13434 12592 13445 12626
rect 13479 12592 13490 12626
rect 13434 12473 13490 12592
rect 13520 12661 13576 12673
rect 13520 12627 13531 12661
rect 13565 12627 13576 12661
rect 13520 12473 13576 12627
rect 13606 12653 13662 12673
rect 13606 12619 13617 12653
rect 13651 12619 13662 12653
rect 13606 12585 13662 12619
rect 13606 12551 13617 12585
rect 13651 12551 13662 12585
rect 13606 12517 13662 12551
rect 13606 12483 13617 12517
rect 13651 12483 13662 12517
rect 13606 12473 13662 12483
rect 13692 12647 13752 12673
rect 13692 12613 13703 12647
rect 13737 12613 13752 12647
rect 13692 12579 13752 12613
rect 13692 12545 13703 12579
rect 13737 12545 13752 12579
rect 13692 12473 13752 12545
rect 13807 12653 13859 12673
rect 13807 12619 13815 12653
rect 13849 12619 13859 12653
rect 13807 12585 13859 12619
rect 13807 12551 13815 12585
rect 13849 12551 13859 12585
rect 13807 12515 13859 12551
rect 13889 12653 13947 12673
rect 13889 12619 13901 12653
rect 13935 12619 13947 12653
rect 13889 12585 13947 12619
rect 13889 12551 13901 12585
rect 13935 12551 13947 12585
rect 13889 12515 13947 12551
rect 13977 12653 14029 12673
rect 13977 12619 13987 12653
rect 14021 12619 14029 12653
rect 13977 12572 14029 12619
rect 14105 12635 14157 12673
rect 14105 12601 14113 12635
rect 14147 12601 14157 12635
rect 14105 12589 14157 12601
rect 14187 12661 14241 12673
rect 14187 12627 14197 12661
rect 14231 12627 14241 12661
rect 14187 12589 14241 12627
rect 14341 12635 14393 12673
rect 14341 12601 14351 12635
rect 14385 12601 14393 12635
rect 14341 12589 14393 12601
rect 14447 12635 14499 12673
rect 14447 12601 14455 12635
rect 14489 12601 14499 12635
rect 14447 12589 14499 12601
rect 14599 12661 14664 12673
rect 14599 12627 14614 12661
rect 14648 12627 14664 12661
rect 14599 12589 14664 12627
rect 13977 12538 13987 12572
rect 14021 12538 14029 12572
rect 13977 12515 14029 12538
rect 14614 12473 14664 12589
rect 14694 12635 14746 12673
rect 14694 12601 14704 12635
rect 14738 12601 14746 12635
rect 14694 12473 14746 12601
rect 15095 12653 15147 12667
rect 15095 12619 15103 12653
rect 15137 12619 15147 12653
rect 15095 12585 15147 12619
rect 15095 12551 15103 12585
rect 15137 12551 15147 12585
rect 15095 12539 15147 12551
rect 15177 12637 15231 12667
rect 15177 12603 15187 12637
rect 15221 12603 15231 12637
rect 15177 12539 15231 12603
rect 15261 12653 15313 12667
rect 15261 12619 15271 12653
rect 15305 12619 15313 12653
rect 15261 12585 15313 12619
rect 15446 12661 15498 12673
rect 15446 12627 15454 12661
rect 15488 12627 15498 12661
rect 15446 12589 15498 12627
rect 15528 12653 15590 12673
rect 15528 12619 15538 12653
rect 15572 12619 15590 12653
rect 15528 12589 15590 12619
rect 15620 12659 15689 12673
rect 15620 12625 15631 12659
rect 15665 12625 15689 12659
rect 15620 12589 15689 12625
rect 15719 12635 15829 12673
rect 15719 12601 15785 12635
rect 15819 12601 15829 12635
rect 15719 12589 15829 12601
rect 15859 12651 15926 12673
rect 15859 12617 15882 12651
rect 15916 12617 15926 12651
rect 15859 12589 15926 12617
rect 15956 12635 16008 12673
rect 15956 12601 15966 12635
rect 16000 12601 16008 12635
rect 15956 12589 16008 12601
rect 16071 12661 16123 12673
rect 16071 12627 16079 12661
rect 16113 12627 16123 12661
rect 15261 12551 15271 12585
rect 15305 12551 15313 12585
rect 15261 12539 15313 12551
rect 16071 12505 16123 12627
rect 16153 12653 16222 12673
rect 16153 12619 16167 12653
rect 16201 12619 16222 12653
rect 16153 12589 16222 12619
rect 16252 12660 16308 12673
rect 16252 12626 16264 12660
rect 16298 12626 16308 12660
rect 16252 12589 16308 12626
rect 16338 12589 16392 12673
rect 16422 12661 16500 12673
rect 16422 12627 16456 12661
rect 16490 12627 16500 12661
rect 16422 12589 16500 12627
rect 16530 12635 16584 12673
rect 16530 12601 16540 12635
rect 16574 12601 16584 12635
rect 16530 12589 16584 12601
rect 16614 12661 16668 12673
rect 16614 12627 16626 12661
rect 16660 12627 16668 12661
rect 16614 12589 16668 12627
rect 16733 12661 16799 12673
rect 16733 12627 16755 12661
rect 16789 12627 16799 12661
rect 16733 12593 16799 12627
rect 16153 12505 16207 12589
rect 16733 12559 16755 12593
rect 16789 12559 16799 12593
rect 16733 12545 16799 12559
rect 16749 12473 16799 12545
rect 16829 12625 16881 12673
rect 16829 12591 16839 12625
rect 16873 12591 16881 12625
rect 16829 12557 16881 12591
rect 16829 12523 16839 12557
rect 16873 12523 16881 12557
rect 16829 12473 16881 12523
rect 17027 12653 17080 12673
rect 17027 12619 17035 12653
rect 17069 12619 17080 12653
rect 17027 12531 17080 12619
rect 17027 12497 17035 12531
rect 17069 12497 17080 12531
rect 17027 12473 17080 12497
rect 17110 12661 17176 12673
rect 17110 12627 17121 12661
rect 17155 12627 17176 12661
rect 17110 12593 17176 12627
rect 17110 12559 17121 12593
rect 17155 12559 17176 12593
rect 17110 12473 17176 12559
rect 17206 12626 17262 12673
rect 17206 12592 17217 12626
rect 17251 12592 17262 12626
rect 17206 12473 17262 12592
rect 17292 12661 17348 12673
rect 17292 12627 17303 12661
rect 17337 12627 17348 12661
rect 17292 12473 17348 12627
rect 17378 12653 17434 12673
rect 17378 12619 17389 12653
rect 17423 12619 17434 12653
rect 17378 12585 17434 12619
rect 17378 12551 17389 12585
rect 17423 12551 17434 12585
rect 17378 12517 17434 12551
rect 17378 12483 17389 12517
rect 17423 12483 17434 12517
rect 17378 12473 17434 12483
rect 17464 12647 17524 12673
rect 17763 12661 17815 12673
rect 17464 12613 17475 12647
rect 17509 12613 17524 12647
rect 17464 12579 17524 12613
rect 17464 12545 17475 12579
rect 17509 12545 17524 12579
rect 17464 12473 17524 12545
rect 17763 12627 17771 12661
rect 17805 12627 17815 12661
rect 17763 12559 17815 12627
rect 17763 12525 17771 12559
rect 17805 12525 17815 12559
rect 17763 12499 17815 12525
rect 18209 12661 18261 12673
rect 18209 12627 18219 12661
rect 18253 12627 18261 12661
rect 18209 12559 18261 12627
rect 18209 12525 18219 12559
rect 18253 12525 18261 12559
rect 18209 12499 18261 12525
rect 18315 12661 18367 12673
rect 18315 12627 18323 12661
rect 18357 12627 18367 12661
rect 18315 12499 18367 12627
rect 19313 12661 19365 12673
rect 19313 12627 19323 12661
rect 19357 12627 19365 12661
rect 19313 12499 19365 12627
rect 19419 12653 19472 12673
rect 19419 12619 19427 12653
rect 19461 12619 19472 12653
rect 19419 12531 19472 12619
rect 19419 12497 19427 12531
rect 19461 12497 19472 12531
rect 19419 12473 19472 12497
rect 19502 12661 19568 12673
rect 19502 12627 19513 12661
rect 19547 12627 19568 12661
rect 19502 12593 19568 12627
rect 19502 12559 19513 12593
rect 19547 12559 19568 12593
rect 19502 12473 19568 12559
rect 19598 12626 19654 12673
rect 19598 12592 19609 12626
rect 19643 12592 19654 12626
rect 19598 12473 19654 12592
rect 19684 12661 19740 12673
rect 19684 12627 19695 12661
rect 19729 12627 19740 12661
rect 19684 12473 19740 12627
rect 19770 12653 19826 12673
rect 19770 12619 19781 12653
rect 19815 12619 19826 12653
rect 19770 12585 19826 12619
rect 19770 12551 19781 12585
rect 19815 12551 19826 12585
rect 19770 12517 19826 12551
rect 19770 12483 19781 12517
rect 19815 12483 19826 12517
rect 19770 12473 19826 12483
rect 19856 12647 19916 12673
rect 19856 12613 19867 12647
rect 19901 12613 19916 12647
rect 19856 12579 19916 12613
rect 19856 12545 19867 12579
rect 19901 12545 19916 12579
rect 19856 12473 19916 12545
rect 19971 12661 20023 12673
rect 19971 12627 19979 12661
rect 20013 12627 20023 12661
rect 19971 12566 20023 12627
rect 19971 12532 19979 12566
rect 20013 12532 20023 12566
rect 19971 12499 20023 12532
rect 20141 12661 20193 12673
rect 20141 12627 20151 12661
rect 20185 12627 20193 12661
rect 20141 12566 20193 12627
rect 20141 12532 20151 12566
rect 20185 12532 20193 12566
rect 20141 12499 20193 12532
rect 29756 6738 29814 6750
rect 29756 6162 29768 6738
rect 29802 6162 29814 6738
rect 29756 6150 29814 6162
rect 30014 6738 30072 6750
rect 30014 6162 30026 6738
rect 30060 6162 30072 6738
rect 30014 6150 30072 6162
rect 30136 6738 30194 6750
rect 30136 6162 30148 6738
rect 30182 6162 30194 6738
rect 30136 6150 30194 6162
rect 30394 6738 30452 6750
rect 30394 6162 30406 6738
rect 30440 6162 30452 6738
rect 30394 6150 30452 6162
rect 30652 6738 30710 6750
rect 30652 6162 30664 6738
rect 30698 6162 30710 6738
rect 30652 6150 30710 6162
rect 30776 6738 30834 6750
rect 30776 6162 30788 6738
rect 30822 6162 30834 6738
rect 30776 6150 30834 6162
rect 31034 6738 31092 6750
rect 31034 6162 31046 6738
rect 31080 6162 31092 6738
rect 31034 6150 31092 6162
rect 31292 6738 31350 6750
rect 31292 6162 31304 6738
rect 31338 6162 31350 6738
rect 31292 6150 31350 6162
rect 31550 6738 31608 6750
rect 31550 6162 31562 6738
rect 31596 6162 31608 6738
rect 31550 6150 31608 6162
rect 31676 6738 31734 6750
rect 31676 6162 31688 6738
rect 31722 6162 31734 6738
rect 31676 6150 31734 6162
rect 31934 6738 31992 6750
rect 31934 6162 31946 6738
rect 31980 6162 31992 6738
rect 31934 6150 31992 6162
rect 32192 6738 32250 6750
rect 32192 6162 32204 6738
rect 32238 6162 32250 6738
rect 32192 6150 32250 6162
rect 32450 6738 32508 6750
rect 32450 6162 32462 6738
rect 32496 6162 32508 6738
rect 32450 6150 32508 6162
rect 32708 6738 32766 6750
rect 32708 6162 32720 6738
rect 32754 6162 32766 6738
rect 32708 6150 32766 6162
rect 32966 6738 33024 6750
rect 32966 6162 32978 6738
rect 33012 6162 33024 6738
rect 32966 6150 33024 6162
rect 33224 6738 33282 6750
rect 33224 6162 33236 6738
rect 33270 6162 33282 6738
rect 33224 6150 33282 6162
rect 33482 6738 33540 6750
rect 33482 6162 33494 6738
rect 33528 6162 33540 6738
rect 33482 6150 33540 6162
rect 33740 6738 33798 6750
rect 33740 6162 33752 6738
rect 33786 6162 33798 6738
rect 33740 6150 33798 6162
rect 33998 6738 34056 6750
rect 33998 6162 34010 6738
rect 34044 6162 34056 6738
rect 33998 6150 34056 6162
rect 34256 6738 34314 6750
rect 34256 6162 34268 6738
rect 34302 6162 34314 6738
rect 34256 6150 34314 6162
rect 34376 6738 34434 6750
rect 34376 6162 34388 6738
rect 34422 6162 34434 6738
rect 34376 6150 34434 6162
rect 34634 6738 34692 6750
rect 34634 6162 34646 6738
rect 34680 6162 34692 6738
rect 34634 6150 34692 6162
rect 30016 5718 30074 5730
rect 30016 5142 30028 5718
rect 30062 5142 30074 5718
rect 30016 5130 30074 5142
rect 30104 5718 30162 5730
rect 30104 5142 30116 5718
rect 30150 5142 30162 5718
rect 30104 5130 30162 5142
rect 30236 5718 30298 5730
rect 30236 5142 30248 5718
rect 30282 5142 30298 5718
rect 30236 5130 30298 5142
rect 30328 5718 30394 5730
rect 30328 5142 30344 5718
rect 30378 5142 30394 5718
rect 30328 5130 30394 5142
rect 30424 5718 30490 5730
rect 30424 5142 30440 5718
rect 30474 5142 30490 5718
rect 30424 5130 30490 5142
rect 30520 5718 30582 5730
rect 30520 5142 30536 5718
rect 30570 5142 30582 5718
rect 30520 5130 30582 5142
rect 30636 5718 30698 5730
rect 30636 5142 30648 5718
rect 30682 5142 30698 5718
rect 30636 5130 30698 5142
rect 30728 5718 30794 5730
rect 30728 5142 30744 5718
rect 30778 5142 30794 5718
rect 30728 5130 30794 5142
rect 30824 5718 30890 5730
rect 30824 5142 30840 5718
rect 30874 5142 30890 5718
rect 30824 5130 30890 5142
rect 30920 5718 30982 5730
rect 30920 5142 30936 5718
rect 30970 5142 30982 5718
rect 30920 5130 30982 5142
rect 31036 5718 31094 5730
rect 31036 5142 31048 5718
rect 31082 5142 31094 5718
rect 31036 5130 31094 5142
rect 31124 5718 31182 5730
rect 31124 5142 31136 5718
rect 31170 5142 31182 5718
rect 31124 5130 31182 5142
rect 1426 4218 1484 4230
rect 1426 3242 1438 4218
rect 1472 3242 1484 4218
rect 1426 3230 1484 3242
rect 1514 4218 1572 4230
rect 1514 3242 1526 4218
rect 1560 3242 1572 4218
rect 1839 4211 1901 4223
rect 1514 3230 1572 3242
rect 1626 3818 1684 3830
rect 1626 3242 1638 3818
rect 1672 3242 1684 3818
rect 1626 3230 1684 3242
rect 1714 3818 1772 3830
rect 1714 3242 1726 3818
rect 1760 3242 1772 3818
rect 1714 3230 1772 3242
rect 1839 3235 1851 4211
rect 1885 3235 1901 4211
rect 1839 3223 1901 3235
rect 1931 4211 1997 4223
rect 1931 3235 1947 4211
rect 1981 3235 1997 4211
rect 1931 3223 1997 3235
rect 2027 4211 2093 4223
rect 2027 3235 2043 4211
rect 2077 3235 2093 4211
rect 2027 3223 2093 3235
rect 2123 4211 2189 4223
rect 2123 3235 2139 4211
rect 2173 3235 2189 4211
rect 2123 3223 2189 3235
rect 2219 4211 2285 4223
rect 2219 3235 2235 4211
rect 2269 3235 2285 4211
rect 2219 3223 2285 3235
rect 2315 4211 2381 4223
rect 2315 3235 2331 4211
rect 2365 3235 2381 4211
rect 2315 3223 2381 3235
rect 2411 4211 2477 4223
rect 2411 3235 2427 4211
rect 2461 3235 2477 4211
rect 2411 3223 2477 3235
rect 2507 4211 2573 4223
rect 2507 3235 2523 4211
rect 2557 3235 2573 4211
rect 2507 3223 2573 3235
rect 2603 4211 2669 4223
rect 2603 3235 2619 4211
rect 2653 3235 2669 4211
rect 2603 3223 2669 3235
rect 2699 4211 2765 4223
rect 2699 3235 2715 4211
rect 2749 3235 2765 4211
rect 2699 3223 2765 3235
rect 2795 4211 2861 4223
rect 2795 3235 2811 4211
rect 2845 3235 2861 4211
rect 2795 3223 2861 3235
rect 2891 4211 2957 4223
rect 2891 3235 2907 4211
rect 2941 3235 2957 4211
rect 2891 3223 2957 3235
rect 2987 4211 3049 4223
rect 2987 3235 3003 4211
rect 3037 3235 3049 4211
rect 2987 3223 3049 3235
rect 3126 4218 3184 4230
rect 3126 3242 3138 4218
rect 3172 3242 3184 4218
rect 3126 3230 3184 3242
rect 3214 4218 3272 4230
rect 3214 3242 3226 4218
rect 3260 3242 3272 4218
rect 3214 3230 3272 3242
rect 4726 4218 4784 4230
rect 4726 3242 4738 4218
rect 4772 3242 4784 4218
rect 4726 3230 4784 3242
rect 4814 4218 4872 4230
rect 4814 3242 4826 4218
rect 4860 3242 4872 4218
rect 5139 4211 5201 4223
rect 4814 3230 4872 3242
rect 4926 3818 4984 3830
rect 4926 3242 4938 3818
rect 4972 3242 4984 3818
rect 4926 3230 4984 3242
rect 5014 3818 5072 3830
rect 5014 3242 5026 3818
rect 5060 3242 5072 3818
rect 5014 3230 5072 3242
rect 5139 3235 5151 4211
rect 5185 3235 5201 4211
rect 5139 3223 5201 3235
rect 5231 4211 5297 4223
rect 5231 3235 5247 4211
rect 5281 3235 5297 4211
rect 5231 3223 5297 3235
rect 5327 4211 5393 4223
rect 5327 3235 5343 4211
rect 5377 3235 5393 4211
rect 5327 3223 5393 3235
rect 5423 4211 5489 4223
rect 5423 3235 5439 4211
rect 5473 3235 5489 4211
rect 5423 3223 5489 3235
rect 5519 4211 5585 4223
rect 5519 3235 5535 4211
rect 5569 3235 5585 4211
rect 5519 3223 5585 3235
rect 5615 4211 5681 4223
rect 5615 3235 5631 4211
rect 5665 3235 5681 4211
rect 5615 3223 5681 3235
rect 5711 4211 5777 4223
rect 5711 3235 5727 4211
rect 5761 3235 5777 4211
rect 5711 3223 5777 3235
rect 5807 4211 5873 4223
rect 5807 3235 5823 4211
rect 5857 3235 5873 4211
rect 5807 3223 5873 3235
rect 5903 4211 5969 4223
rect 5903 3235 5919 4211
rect 5953 3235 5969 4211
rect 5903 3223 5969 3235
rect 5999 4211 6065 4223
rect 5999 3235 6015 4211
rect 6049 3235 6065 4211
rect 5999 3223 6065 3235
rect 6095 4211 6161 4223
rect 6095 3235 6111 4211
rect 6145 3235 6161 4211
rect 6095 3223 6161 3235
rect 6191 4211 6257 4223
rect 6191 3235 6207 4211
rect 6241 3235 6257 4211
rect 6191 3223 6257 3235
rect 6287 4211 6349 4223
rect 6287 3235 6303 4211
rect 6337 3235 6349 4211
rect 6287 3223 6349 3235
rect 6426 4218 6484 4230
rect 6426 3242 6438 4218
rect 6472 3242 6484 4218
rect 6426 3230 6484 3242
rect 6514 4218 6572 4230
rect 6514 3242 6526 4218
rect 6560 3242 6572 4218
rect 6514 3230 6572 3242
rect 8026 4218 8084 4230
rect 8026 3242 8038 4218
rect 8072 3242 8084 4218
rect 8026 3230 8084 3242
rect 8114 4218 8172 4230
rect 8114 3242 8126 4218
rect 8160 3242 8172 4218
rect 8439 4211 8501 4223
rect 8114 3230 8172 3242
rect 8226 3818 8284 3830
rect 8226 3242 8238 3818
rect 8272 3242 8284 3818
rect 8226 3230 8284 3242
rect 8314 3818 8372 3830
rect 8314 3242 8326 3818
rect 8360 3242 8372 3818
rect 8314 3230 8372 3242
rect 8439 3235 8451 4211
rect 8485 3235 8501 4211
rect 8439 3223 8501 3235
rect 8531 4211 8597 4223
rect 8531 3235 8547 4211
rect 8581 3235 8597 4211
rect 8531 3223 8597 3235
rect 8627 4211 8693 4223
rect 8627 3235 8643 4211
rect 8677 3235 8693 4211
rect 8627 3223 8693 3235
rect 8723 4211 8789 4223
rect 8723 3235 8739 4211
rect 8773 3235 8789 4211
rect 8723 3223 8789 3235
rect 8819 4211 8885 4223
rect 8819 3235 8835 4211
rect 8869 3235 8885 4211
rect 8819 3223 8885 3235
rect 8915 4211 8981 4223
rect 8915 3235 8931 4211
rect 8965 3235 8981 4211
rect 8915 3223 8981 3235
rect 9011 4211 9077 4223
rect 9011 3235 9027 4211
rect 9061 3235 9077 4211
rect 9011 3223 9077 3235
rect 9107 4211 9173 4223
rect 9107 3235 9123 4211
rect 9157 3235 9173 4211
rect 9107 3223 9173 3235
rect 9203 4211 9269 4223
rect 9203 3235 9219 4211
rect 9253 3235 9269 4211
rect 9203 3223 9269 3235
rect 9299 4211 9365 4223
rect 9299 3235 9315 4211
rect 9349 3235 9365 4211
rect 9299 3223 9365 3235
rect 9395 4211 9461 4223
rect 9395 3235 9411 4211
rect 9445 3235 9461 4211
rect 9395 3223 9461 3235
rect 9491 4211 9557 4223
rect 9491 3235 9507 4211
rect 9541 3235 9557 4211
rect 9491 3223 9557 3235
rect 9587 4211 9649 4223
rect 9587 3235 9603 4211
rect 9637 3235 9649 4211
rect 9587 3223 9649 3235
rect 9726 4218 9784 4230
rect 9726 3242 9738 4218
rect 9772 3242 9784 4218
rect 9726 3230 9784 3242
rect 9814 4218 9872 4230
rect 9814 3242 9826 4218
rect 9860 3242 9872 4218
rect 9814 3230 9872 3242
rect 11326 4218 11384 4230
rect 11326 3242 11338 4218
rect 11372 3242 11384 4218
rect 11326 3230 11384 3242
rect 11414 4218 11472 4230
rect 11414 3242 11426 4218
rect 11460 3242 11472 4218
rect 11739 4211 11801 4223
rect 11414 3230 11472 3242
rect 11526 3818 11584 3830
rect 11526 3242 11538 3818
rect 11572 3242 11584 3818
rect 11526 3230 11584 3242
rect 11614 3818 11672 3830
rect 11614 3242 11626 3818
rect 11660 3242 11672 3818
rect 11614 3230 11672 3242
rect 11739 3235 11751 4211
rect 11785 3235 11801 4211
rect 11739 3223 11801 3235
rect 11831 4211 11897 4223
rect 11831 3235 11847 4211
rect 11881 3235 11897 4211
rect 11831 3223 11897 3235
rect 11927 4211 11993 4223
rect 11927 3235 11943 4211
rect 11977 3235 11993 4211
rect 11927 3223 11993 3235
rect 12023 4211 12089 4223
rect 12023 3235 12039 4211
rect 12073 3235 12089 4211
rect 12023 3223 12089 3235
rect 12119 4211 12185 4223
rect 12119 3235 12135 4211
rect 12169 3235 12185 4211
rect 12119 3223 12185 3235
rect 12215 4211 12281 4223
rect 12215 3235 12231 4211
rect 12265 3235 12281 4211
rect 12215 3223 12281 3235
rect 12311 4211 12377 4223
rect 12311 3235 12327 4211
rect 12361 3235 12377 4211
rect 12311 3223 12377 3235
rect 12407 4211 12473 4223
rect 12407 3235 12423 4211
rect 12457 3235 12473 4211
rect 12407 3223 12473 3235
rect 12503 4211 12569 4223
rect 12503 3235 12519 4211
rect 12553 3235 12569 4211
rect 12503 3223 12569 3235
rect 12599 4211 12665 4223
rect 12599 3235 12615 4211
rect 12649 3235 12665 4211
rect 12599 3223 12665 3235
rect 12695 4211 12761 4223
rect 12695 3235 12711 4211
rect 12745 3235 12761 4211
rect 12695 3223 12761 3235
rect 12791 4211 12857 4223
rect 12791 3235 12807 4211
rect 12841 3235 12857 4211
rect 12791 3223 12857 3235
rect 12887 4211 12949 4223
rect 12887 3235 12903 4211
rect 12937 3235 12949 4211
rect 12887 3223 12949 3235
rect 13026 4218 13084 4230
rect 13026 3242 13038 4218
rect 13072 3242 13084 4218
rect 13026 3230 13084 3242
rect 13114 4218 13172 4230
rect 13114 3242 13126 4218
rect 13160 3242 13172 4218
rect 13114 3230 13172 3242
rect 14926 4218 14984 4230
rect 14926 3242 14938 4218
rect 14972 3242 14984 4218
rect 14926 3230 14984 3242
rect 15014 4218 15072 4230
rect 15014 3242 15026 4218
rect 15060 3242 15072 4218
rect 15339 4211 15401 4223
rect 15014 3230 15072 3242
rect 15126 3818 15184 3830
rect 15126 3242 15138 3818
rect 15172 3242 15184 3818
rect 15126 3230 15184 3242
rect 15214 3818 15272 3830
rect 15214 3242 15226 3818
rect 15260 3242 15272 3818
rect 15214 3230 15272 3242
rect 15339 3235 15351 4211
rect 15385 3235 15401 4211
rect 15339 3223 15401 3235
rect 15431 4211 15497 4223
rect 15431 3235 15447 4211
rect 15481 3235 15497 4211
rect 15431 3223 15497 3235
rect 15527 4211 15593 4223
rect 15527 3235 15543 4211
rect 15577 3235 15593 4211
rect 15527 3223 15593 3235
rect 15623 4211 15689 4223
rect 15623 3235 15639 4211
rect 15673 3235 15689 4211
rect 15623 3223 15689 3235
rect 15719 4211 15785 4223
rect 15719 3235 15735 4211
rect 15769 3235 15785 4211
rect 15719 3223 15785 3235
rect 15815 4211 15881 4223
rect 15815 3235 15831 4211
rect 15865 3235 15881 4211
rect 15815 3223 15881 3235
rect 15911 4211 15977 4223
rect 15911 3235 15927 4211
rect 15961 3235 15977 4211
rect 15911 3223 15977 3235
rect 16007 4211 16073 4223
rect 16007 3235 16023 4211
rect 16057 3235 16073 4211
rect 16007 3223 16073 3235
rect 16103 4211 16169 4223
rect 16103 3235 16119 4211
rect 16153 3235 16169 4211
rect 16103 3223 16169 3235
rect 16199 4211 16265 4223
rect 16199 3235 16215 4211
rect 16249 3235 16265 4211
rect 16199 3223 16265 3235
rect 16295 4211 16361 4223
rect 16295 3235 16311 4211
rect 16345 3235 16361 4211
rect 16295 3223 16361 3235
rect 16391 4211 16457 4223
rect 16391 3235 16407 4211
rect 16441 3235 16457 4211
rect 16391 3223 16457 3235
rect 16487 4211 16549 4223
rect 16487 3235 16503 4211
rect 16537 3235 16549 4211
rect 16487 3223 16549 3235
rect 16626 4218 16684 4230
rect 16626 3242 16638 4218
rect 16672 3242 16684 4218
rect 16626 3230 16684 3242
rect 16714 4218 16772 4230
rect 16714 3242 16726 4218
rect 16760 3242 16772 4218
rect 16714 3230 16772 3242
rect 18426 4218 18484 4230
rect 18426 3242 18438 4218
rect 18472 3242 18484 4218
rect 18426 3230 18484 3242
rect 18514 4218 18572 4230
rect 18514 3242 18526 4218
rect 18560 3242 18572 4218
rect 18839 4211 18901 4223
rect 18514 3230 18572 3242
rect 18626 3818 18684 3830
rect 18626 3242 18638 3818
rect 18672 3242 18684 3818
rect 18626 3230 18684 3242
rect 18714 3818 18772 3830
rect 18714 3242 18726 3818
rect 18760 3242 18772 3818
rect 18714 3230 18772 3242
rect 18839 3235 18851 4211
rect 18885 3235 18901 4211
rect 18839 3223 18901 3235
rect 18931 4211 18997 4223
rect 18931 3235 18947 4211
rect 18981 3235 18997 4211
rect 18931 3223 18997 3235
rect 19027 4211 19093 4223
rect 19027 3235 19043 4211
rect 19077 3235 19093 4211
rect 19027 3223 19093 3235
rect 19123 4211 19189 4223
rect 19123 3235 19139 4211
rect 19173 3235 19189 4211
rect 19123 3223 19189 3235
rect 19219 4211 19285 4223
rect 19219 3235 19235 4211
rect 19269 3235 19285 4211
rect 19219 3223 19285 3235
rect 19315 4211 19381 4223
rect 19315 3235 19331 4211
rect 19365 3235 19381 4211
rect 19315 3223 19381 3235
rect 19411 4211 19477 4223
rect 19411 3235 19427 4211
rect 19461 3235 19477 4211
rect 19411 3223 19477 3235
rect 19507 4211 19573 4223
rect 19507 3235 19523 4211
rect 19557 3235 19573 4211
rect 19507 3223 19573 3235
rect 19603 4211 19669 4223
rect 19603 3235 19619 4211
rect 19653 3235 19669 4211
rect 19603 3223 19669 3235
rect 19699 4211 19765 4223
rect 19699 3235 19715 4211
rect 19749 3235 19765 4211
rect 19699 3223 19765 3235
rect 19795 4211 19861 4223
rect 19795 3235 19811 4211
rect 19845 3235 19861 4211
rect 19795 3223 19861 3235
rect 19891 4211 19957 4223
rect 19891 3235 19907 4211
rect 19941 3235 19957 4211
rect 19891 3223 19957 3235
rect 19987 4211 20049 4223
rect 19987 3235 20003 4211
rect 20037 3235 20049 4211
rect 19987 3223 20049 3235
rect 20126 4218 20184 4230
rect 20126 3242 20138 4218
rect 20172 3242 20184 4218
rect 20126 3230 20184 3242
rect 20214 4218 20272 4230
rect 20214 3242 20226 4218
rect 20260 3242 20272 4218
rect 20214 3230 20272 3242
rect 22126 4218 22184 4230
rect 22126 3242 22138 4218
rect 22172 3242 22184 4218
rect 22126 3230 22184 3242
rect 22214 4218 22272 4230
rect 22214 3242 22226 4218
rect 22260 3242 22272 4218
rect 22539 4211 22601 4223
rect 22214 3230 22272 3242
rect 22326 3818 22384 3830
rect 22326 3242 22338 3818
rect 22372 3242 22384 3818
rect 22326 3230 22384 3242
rect 22414 3818 22472 3830
rect 22414 3242 22426 3818
rect 22460 3242 22472 3818
rect 22414 3230 22472 3242
rect 22539 3235 22551 4211
rect 22585 3235 22601 4211
rect 22539 3223 22601 3235
rect 22631 4211 22697 4223
rect 22631 3235 22647 4211
rect 22681 3235 22697 4211
rect 22631 3223 22697 3235
rect 22727 4211 22793 4223
rect 22727 3235 22743 4211
rect 22777 3235 22793 4211
rect 22727 3223 22793 3235
rect 22823 4211 22889 4223
rect 22823 3235 22839 4211
rect 22873 3235 22889 4211
rect 22823 3223 22889 3235
rect 22919 4211 22985 4223
rect 22919 3235 22935 4211
rect 22969 3235 22985 4211
rect 22919 3223 22985 3235
rect 23015 4211 23081 4223
rect 23015 3235 23031 4211
rect 23065 3235 23081 4211
rect 23015 3223 23081 3235
rect 23111 4211 23177 4223
rect 23111 3235 23127 4211
rect 23161 3235 23177 4211
rect 23111 3223 23177 3235
rect 23207 4211 23273 4223
rect 23207 3235 23223 4211
rect 23257 3235 23273 4211
rect 23207 3223 23273 3235
rect 23303 4211 23369 4223
rect 23303 3235 23319 4211
rect 23353 3235 23369 4211
rect 23303 3223 23369 3235
rect 23399 4211 23465 4223
rect 23399 3235 23415 4211
rect 23449 3235 23465 4211
rect 23399 3223 23465 3235
rect 23495 4211 23561 4223
rect 23495 3235 23511 4211
rect 23545 3235 23561 4211
rect 23495 3223 23561 3235
rect 23591 4211 23657 4223
rect 23591 3235 23607 4211
rect 23641 3235 23657 4211
rect 23591 3223 23657 3235
rect 23687 4211 23749 4223
rect 23687 3235 23703 4211
rect 23737 3235 23749 4211
rect 23687 3223 23749 3235
rect 23826 4218 23884 4230
rect 23826 3242 23838 4218
rect 23872 3242 23884 4218
rect 23826 3230 23884 3242
rect 23914 4218 23972 4230
rect 23914 3242 23926 4218
rect 23960 3242 23972 4218
rect 23914 3230 23972 3242
rect 25926 4218 25984 4230
rect 25926 3242 25938 4218
rect 25972 3242 25984 4218
rect 25926 3230 25984 3242
rect 26014 4218 26072 4230
rect 26014 3242 26026 4218
rect 26060 3242 26072 4218
rect 26339 4211 26401 4223
rect 26014 3230 26072 3242
rect 26126 3818 26184 3830
rect 26126 3242 26138 3818
rect 26172 3242 26184 3818
rect 26126 3230 26184 3242
rect 26214 3818 26272 3830
rect 26214 3242 26226 3818
rect 26260 3242 26272 3818
rect 26214 3230 26272 3242
rect 26339 3235 26351 4211
rect 26385 3235 26401 4211
rect 26339 3223 26401 3235
rect 26431 4211 26497 4223
rect 26431 3235 26447 4211
rect 26481 3235 26497 4211
rect 26431 3223 26497 3235
rect 26527 4211 26593 4223
rect 26527 3235 26543 4211
rect 26577 3235 26593 4211
rect 26527 3223 26593 3235
rect 26623 4211 26689 4223
rect 26623 3235 26639 4211
rect 26673 3235 26689 4211
rect 26623 3223 26689 3235
rect 26719 4211 26785 4223
rect 26719 3235 26735 4211
rect 26769 3235 26785 4211
rect 26719 3223 26785 3235
rect 26815 4211 26881 4223
rect 26815 3235 26831 4211
rect 26865 3235 26881 4211
rect 26815 3223 26881 3235
rect 26911 4211 26977 4223
rect 26911 3235 26927 4211
rect 26961 3235 26977 4211
rect 26911 3223 26977 3235
rect 27007 4211 27073 4223
rect 27007 3235 27023 4211
rect 27057 3235 27073 4211
rect 27007 3223 27073 3235
rect 27103 4211 27169 4223
rect 27103 3235 27119 4211
rect 27153 3235 27169 4211
rect 27103 3223 27169 3235
rect 27199 4211 27265 4223
rect 27199 3235 27215 4211
rect 27249 3235 27265 4211
rect 27199 3223 27265 3235
rect 27295 4211 27361 4223
rect 27295 3235 27311 4211
rect 27345 3235 27361 4211
rect 27295 3223 27361 3235
rect 27391 4211 27457 4223
rect 27391 3235 27407 4211
rect 27441 3235 27457 4211
rect 27391 3223 27457 3235
rect 27487 4211 27549 4223
rect 27487 3235 27503 4211
rect 27537 3235 27549 4211
rect 27487 3223 27549 3235
rect 27626 4218 27684 4230
rect 27626 3242 27638 4218
rect 27672 3242 27684 4218
rect 27626 3230 27684 3242
rect 27714 4218 27772 4230
rect 27714 3242 27726 4218
rect 27760 3242 27772 4218
rect 27714 3230 27772 3242
<< ndiffc >>
rect 4983 27294 5017 27328
rect 5155 27294 5189 27328
rect 5259 27294 5293 27328
rect 5431 27294 5465 27328
rect 5542 27311 5576 27345
rect 5628 27289 5662 27323
rect 5714 27311 5748 27345
rect 5800 27289 5834 27323
rect 5897 27311 5931 27345
rect 5983 27307 6017 27341
rect 6179 27296 6213 27330
rect 7179 27296 7213 27330
rect 7375 27294 7409 27328
rect 7547 27294 7581 27328
rect 7651 27296 7685 27330
rect 8651 27296 8685 27330
rect 8755 27296 8789 27330
rect 9755 27296 9789 27330
rect 10135 27302 10169 27336
rect 10221 27315 10255 27349
rect 10307 27285 10341 27319
rect 10595 27296 10629 27330
rect 11227 27296 11261 27330
rect 11331 27296 11365 27330
rect 12331 27296 12365 27330
rect 12527 27294 12561 27328
rect 12699 27294 12733 27328
rect 12803 27296 12837 27330
rect 13803 27296 13837 27330
rect 13907 27296 13941 27330
rect 14907 27296 14941 27330
rect 15103 27294 15137 27328
rect 15275 27294 15309 27328
rect 15379 27296 15413 27330
rect 16379 27296 16413 27330
rect 16483 27296 16517 27330
rect 17483 27296 17517 27330
rect 17771 27296 17805 27330
rect 18403 27296 18437 27330
rect 18514 27311 18548 27345
rect 18600 27289 18634 27323
rect 18686 27311 18720 27345
rect 18772 27289 18806 27323
rect 18869 27311 18903 27345
rect 18955 27307 18989 27341
rect 19243 27296 19277 27330
rect 19875 27296 19909 27330
rect 19979 27294 20013 27328
rect 20151 27294 20185 27328
rect 4983 26400 5017 26434
rect 5155 26400 5189 26434
rect 5443 26398 5477 26432
rect 6075 26398 6109 26432
rect 6179 26398 6213 26432
rect 7179 26398 7213 26432
rect 7467 26398 7501 26432
rect 7915 26398 7949 26432
rect 8019 26398 8053 26432
rect 9019 26398 9053 26432
rect 9123 26398 9157 26432
rect 10123 26398 10157 26432
rect 10227 26398 10261 26432
rect 11227 26398 11261 26432
rect 11331 26398 11365 26432
rect 12331 26398 12365 26432
rect 12619 26398 12653 26432
rect 13067 26398 13101 26432
rect 13171 26398 13205 26432
rect 14171 26398 14205 26432
rect 14275 26398 14309 26432
rect 15275 26398 15309 26432
rect 15379 26398 15413 26432
rect 16379 26398 16413 26432
rect 16483 26398 16517 26432
rect 17483 26398 17517 26432
rect 17771 26398 17805 26432
rect 18771 26398 18805 26432
rect 18875 26398 18909 26432
rect 19875 26398 19909 26432
rect 19979 26400 20013 26434
rect 20151 26400 20185 26434
rect 4983 26206 5017 26240
rect 5155 26206 5189 26240
rect 5443 26208 5477 26242
rect 6443 26208 6477 26242
rect 6547 26208 6581 26242
rect 7547 26208 7581 26242
rect 7651 26208 7685 26242
rect 8651 26208 8685 26242
rect 8755 26208 8789 26242
rect 9755 26208 9789 26242
rect 10043 26208 10077 26242
rect 10491 26208 10525 26242
rect 10595 26208 10629 26242
rect 11595 26208 11629 26242
rect 11699 26208 11733 26242
rect 12699 26208 12733 26242
rect 12803 26208 12837 26242
rect 13803 26208 13837 26242
rect 13907 26208 13941 26242
rect 14907 26208 14941 26242
rect 15195 26201 15229 26235
rect 15459 26201 15493 26235
rect 15563 26208 15597 26242
rect 16563 26208 16597 26242
rect 16667 26208 16701 26242
rect 17667 26208 17701 26242
rect 17771 26208 17805 26242
rect 18771 26208 18805 26242
rect 18875 26208 18909 26242
rect 19875 26208 19909 26242
rect 19979 26206 20013 26240
rect 20151 26206 20185 26240
rect 4983 25312 5017 25346
rect 5155 25312 5189 25346
rect 5443 25310 5477 25344
rect 6075 25310 6109 25344
rect 6179 25310 6213 25344
rect 7179 25310 7213 25344
rect 7467 25310 7501 25344
rect 7915 25310 7949 25344
rect 8019 25310 8053 25344
rect 9019 25310 9053 25344
rect 9123 25310 9157 25344
rect 10123 25310 10157 25344
rect 10227 25310 10261 25344
rect 11227 25310 11261 25344
rect 11331 25310 11365 25344
rect 12331 25310 12365 25344
rect 12619 25310 12653 25344
rect 13067 25310 13101 25344
rect 13171 25310 13205 25344
rect 14171 25310 14205 25344
rect 14275 25310 14309 25344
rect 15275 25310 15309 25344
rect 15379 25310 15413 25344
rect 16379 25310 16413 25344
rect 16483 25310 16517 25344
rect 17483 25310 17517 25344
rect 17771 25310 17805 25344
rect 18771 25310 18805 25344
rect 18875 25310 18909 25344
rect 19875 25310 19909 25344
rect 19979 25312 20013 25346
rect 20151 25312 20185 25346
rect 4983 25118 5017 25152
rect 5155 25118 5189 25152
rect 5443 25120 5477 25154
rect 6443 25120 6477 25154
rect 6547 25120 6581 25154
rect 7547 25120 7581 25154
rect 7651 25120 7685 25154
rect 8651 25120 8685 25154
rect 8755 25120 8789 25154
rect 9755 25120 9789 25154
rect 10043 25120 10077 25154
rect 10491 25120 10525 25154
rect 10595 25120 10629 25154
rect 11595 25120 11629 25154
rect 11699 25120 11733 25154
rect 12699 25120 12733 25154
rect 12803 25120 12837 25154
rect 13803 25120 13837 25154
rect 13907 25120 13941 25154
rect 14907 25120 14941 25154
rect 15195 25113 15229 25147
rect 15459 25113 15493 25147
rect 15563 25120 15597 25154
rect 16563 25120 16597 25154
rect 16667 25120 16701 25154
rect 17667 25120 17701 25154
rect 17771 25120 17805 25154
rect 18771 25120 18805 25154
rect 18875 25120 18909 25154
rect 19875 25120 19909 25154
rect 19979 25118 20013 25152
rect 20151 25118 20185 25152
rect 4983 24224 5017 24258
rect 5155 24224 5189 24258
rect 5443 24222 5477 24256
rect 6075 24222 6109 24256
rect 6179 24222 6213 24256
rect 7179 24222 7213 24256
rect 7467 24222 7501 24256
rect 7915 24222 7949 24256
rect 8019 24222 8053 24256
rect 9019 24222 9053 24256
rect 9123 24222 9157 24256
rect 10123 24222 10157 24256
rect 10227 24222 10261 24256
rect 11227 24222 11261 24256
rect 11331 24222 11365 24256
rect 12331 24222 12365 24256
rect 12619 24222 12653 24256
rect 13067 24222 13101 24256
rect 13171 24222 13205 24256
rect 14171 24222 14205 24256
rect 14275 24222 14309 24256
rect 15275 24222 15309 24256
rect 15379 24222 15413 24256
rect 16379 24222 16413 24256
rect 16483 24222 16517 24256
rect 17483 24222 17517 24256
rect 17771 24222 17805 24256
rect 18771 24222 18805 24256
rect 18875 24222 18909 24256
rect 19875 24222 19909 24256
rect 19979 24224 20013 24258
rect 20151 24224 20185 24258
rect 4983 24030 5017 24064
rect 5155 24030 5189 24064
rect 5443 24032 5477 24066
rect 6443 24032 6477 24066
rect 6547 24032 6581 24066
rect 7547 24032 7581 24066
rect 7651 24032 7685 24066
rect 8651 24032 8685 24066
rect 8755 24032 8789 24066
rect 9755 24032 9789 24066
rect 10043 24032 10077 24066
rect 10491 24032 10525 24066
rect 10595 24032 10629 24066
rect 11595 24032 11629 24066
rect 11699 24032 11733 24066
rect 12699 24032 12733 24066
rect 12803 24032 12837 24066
rect 13803 24032 13837 24066
rect 13907 24032 13941 24066
rect 14907 24032 14941 24066
rect 15195 24025 15229 24059
rect 15459 24025 15493 24059
rect 15563 24032 15597 24066
rect 16563 24032 16597 24066
rect 16667 24032 16701 24066
rect 17667 24032 17701 24066
rect 17771 24032 17805 24066
rect 18771 24032 18805 24066
rect 18875 24032 18909 24066
rect 19875 24032 19909 24066
rect 19979 24030 20013 24064
rect 20151 24030 20185 24064
rect 4983 23136 5017 23170
rect 5155 23136 5189 23170
rect 5443 23134 5477 23168
rect 6075 23134 6109 23168
rect 6179 23134 6213 23168
rect 7179 23134 7213 23168
rect 7467 23134 7501 23168
rect 7915 23134 7949 23168
rect 8019 23134 8053 23168
rect 9019 23134 9053 23168
rect 9123 23134 9157 23168
rect 10123 23134 10157 23168
rect 10227 23134 10261 23168
rect 11227 23134 11261 23168
rect 11331 23134 11365 23168
rect 12331 23134 12365 23168
rect 12619 23134 12653 23168
rect 13067 23134 13101 23168
rect 13171 23134 13205 23168
rect 14171 23134 14205 23168
rect 14275 23134 14309 23168
rect 15275 23134 15309 23168
rect 15379 23134 15413 23168
rect 16379 23134 16413 23168
rect 16483 23134 16517 23168
rect 17483 23134 17517 23168
rect 17771 23134 17805 23168
rect 18771 23134 18805 23168
rect 18875 23134 18909 23168
rect 19875 23134 19909 23168
rect 19979 23136 20013 23170
rect 20151 23136 20185 23170
rect 4983 22942 5017 22976
rect 5155 22942 5189 22976
rect 5443 22944 5477 22978
rect 6443 22944 6477 22978
rect 6547 22944 6581 22978
rect 7547 22944 7581 22978
rect 7651 22944 7685 22978
rect 8651 22944 8685 22978
rect 8755 22944 8789 22978
rect 9755 22944 9789 22978
rect 10043 22944 10077 22978
rect 10491 22944 10525 22978
rect 10595 22944 10629 22978
rect 11595 22944 11629 22978
rect 11699 22944 11733 22978
rect 12699 22944 12733 22978
rect 12803 22944 12837 22978
rect 13803 22944 13837 22978
rect 13907 22944 13941 22978
rect 14907 22944 14941 22978
rect 15195 22937 15229 22971
rect 15459 22937 15493 22971
rect 15563 22944 15597 22978
rect 16563 22944 16597 22978
rect 16667 22944 16701 22978
rect 17667 22944 17701 22978
rect 17771 22944 17805 22978
rect 18771 22944 18805 22978
rect 18875 22944 18909 22978
rect 19875 22944 19909 22978
rect 19979 22942 20013 22976
rect 20151 22942 20185 22976
rect 4983 22048 5017 22082
rect 5155 22048 5189 22082
rect 5443 22046 5477 22080
rect 6075 22046 6109 22080
rect 6179 22046 6213 22080
rect 7179 22046 7213 22080
rect 7467 22046 7501 22080
rect 7915 22046 7949 22080
rect 8019 22046 8053 22080
rect 9019 22046 9053 22080
rect 9123 22046 9157 22080
rect 10123 22046 10157 22080
rect 10227 22046 10261 22080
rect 11227 22046 11261 22080
rect 11331 22046 11365 22080
rect 12331 22046 12365 22080
rect 12619 22046 12653 22080
rect 13067 22046 13101 22080
rect 13171 22046 13205 22080
rect 14171 22046 14205 22080
rect 14275 22046 14309 22080
rect 15275 22046 15309 22080
rect 15379 22046 15413 22080
rect 16379 22046 16413 22080
rect 16483 22046 16517 22080
rect 17483 22046 17517 22080
rect 17771 22046 17805 22080
rect 18771 22046 18805 22080
rect 18875 22046 18909 22080
rect 19875 22046 19909 22080
rect 19979 22048 20013 22082
rect 20151 22048 20185 22082
rect 4983 21854 5017 21888
rect 5155 21854 5189 21888
rect 5443 21856 5477 21890
rect 6443 21856 6477 21890
rect 6547 21856 6581 21890
rect 7547 21856 7581 21890
rect 7651 21856 7685 21890
rect 8651 21856 8685 21890
rect 8755 21856 8789 21890
rect 9755 21856 9789 21890
rect 10043 21856 10077 21890
rect 10491 21856 10525 21890
rect 10595 21856 10629 21890
rect 11595 21856 11629 21890
rect 11699 21856 11733 21890
rect 12699 21856 12733 21890
rect 12803 21856 12837 21890
rect 13803 21856 13837 21890
rect 13907 21856 13941 21890
rect 14907 21856 14941 21890
rect 15195 21849 15229 21883
rect 15459 21849 15493 21883
rect 15563 21856 15597 21890
rect 16563 21856 16597 21890
rect 16667 21856 16701 21890
rect 17667 21856 17701 21890
rect 17771 21856 17805 21890
rect 18771 21856 18805 21890
rect 18875 21856 18909 21890
rect 19875 21856 19909 21890
rect 19979 21854 20013 21888
rect 20151 21854 20185 21888
rect 4983 20960 5017 20994
rect 5155 20960 5189 20994
rect 5443 20958 5477 20992
rect 6075 20958 6109 20992
rect 6179 20958 6213 20992
rect 7179 20958 7213 20992
rect 7467 20958 7501 20992
rect 7915 20958 7949 20992
rect 8019 20958 8053 20992
rect 9019 20958 9053 20992
rect 9123 20958 9157 20992
rect 10123 20958 10157 20992
rect 10227 20958 10261 20992
rect 11227 20958 11261 20992
rect 11331 20958 11365 20992
rect 12331 20958 12365 20992
rect 12619 20958 12653 20992
rect 13067 20958 13101 20992
rect 13171 20958 13205 20992
rect 14171 20958 14205 20992
rect 14275 20958 14309 20992
rect 15275 20958 15309 20992
rect 15379 20958 15413 20992
rect 16379 20958 16413 20992
rect 16483 20958 16517 20992
rect 17483 20958 17517 20992
rect 17771 20958 17805 20992
rect 18771 20958 18805 20992
rect 18875 20958 18909 20992
rect 19875 20958 19909 20992
rect 19979 20960 20013 20994
rect 20151 20960 20185 20994
rect 4983 20766 5017 20800
rect 5155 20766 5189 20800
rect 5443 20768 5477 20802
rect 6443 20768 6477 20802
rect 6547 20768 6581 20802
rect 7547 20768 7581 20802
rect 7651 20768 7685 20802
rect 8651 20768 8685 20802
rect 8755 20768 8789 20802
rect 9755 20768 9789 20802
rect 10043 20768 10077 20802
rect 10491 20768 10525 20802
rect 10595 20768 10629 20802
rect 11595 20768 11629 20802
rect 11699 20768 11733 20802
rect 12699 20768 12733 20802
rect 12803 20768 12837 20802
rect 13803 20768 13837 20802
rect 13907 20768 13941 20802
rect 14907 20768 14941 20802
rect 15195 20761 15229 20795
rect 15459 20761 15493 20795
rect 15563 20768 15597 20802
rect 16563 20768 16597 20802
rect 16667 20768 16701 20802
rect 17667 20768 17701 20802
rect 17771 20768 17805 20802
rect 18771 20768 18805 20802
rect 18875 20768 18909 20802
rect 19875 20768 19909 20802
rect 19979 20766 20013 20800
rect 20151 20766 20185 20800
rect 4983 19872 5017 19906
rect 5155 19872 5189 19906
rect 5443 19870 5477 19904
rect 6075 19870 6109 19904
rect 6179 19870 6213 19904
rect 7179 19870 7213 19904
rect 7467 19870 7501 19904
rect 7915 19870 7949 19904
rect 8019 19870 8053 19904
rect 9019 19870 9053 19904
rect 9123 19870 9157 19904
rect 10123 19870 10157 19904
rect 10227 19870 10261 19904
rect 11227 19870 11261 19904
rect 11331 19870 11365 19904
rect 12331 19870 12365 19904
rect 12619 19870 12653 19904
rect 13067 19870 13101 19904
rect 13171 19870 13205 19904
rect 14171 19870 14205 19904
rect 14275 19870 14309 19904
rect 15275 19870 15309 19904
rect 15379 19870 15413 19904
rect 16379 19870 16413 19904
rect 16483 19870 16517 19904
rect 17483 19870 17517 19904
rect 17771 19870 17805 19904
rect 18771 19870 18805 19904
rect 18875 19870 18909 19904
rect 19875 19870 19909 19904
rect 19979 19872 20013 19906
rect 20151 19872 20185 19906
rect 4983 19678 5017 19712
rect 5155 19678 5189 19712
rect 5443 19680 5477 19714
rect 6443 19680 6477 19714
rect 6547 19680 6581 19714
rect 7547 19680 7581 19714
rect 7651 19680 7685 19714
rect 8651 19680 8685 19714
rect 8755 19680 8789 19714
rect 9755 19680 9789 19714
rect 10043 19680 10077 19714
rect 10491 19680 10525 19714
rect 10595 19680 10629 19714
rect 11595 19680 11629 19714
rect 11699 19680 11733 19714
rect 12699 19680 12733 19714
rect 12803 19680 12837 19714
rect 13803 19680 13837 19714
rect 13907 19680 13941 19714
rect 14907 19680 14941 19714
rect 15195 19673 15229 19707
rect 15459 19673 15493 19707
rect 15563 19680 15597 19714
rect 16563 19680 16597 19714
rect 16667 19680 16701 19714
rect 17667 19680 17701 19714
rect 17771 19680 17805 19714
rect 18771 19680 18805 19714
rect 18875 19680 18909 19714
rect 19875 19680 19909 19714
rect 19979 19678 20013 19712
rect 20151 19678 20185 19712
rect 4983 18784 5017 18818
rect 5155 18784 5189 18818
rect 5443 18782 5477 18816
rect 6075 18782 6109 18816
rect 6179 18782 6213 18816
rect 7179 18782 7213 18816
rect 7467 18782 7501 18816
rect 7915 18782 7949 18816
rect 8019 18782 8053 18816
rect 9019 18782 9053 18816
rect 9123 18782 9157 18816
rect 10123 18782 10157 18816
rect 10227 18782 10261 18816
rect 11227 18782 11261 18816
rect 11331 18782 11365 18816
rect 12331 18782 12365 18816
rect 12619 18782 12653 18816
rect 13067 18782 13101 18816
rect 13171 18782 13205 18816
rect 14171 18782 14205 18816
rect 14275 18782 14309 18816
rect 15275 18782 15309 18816
rect 15379 18782 15413 18816
rect 16379 18782 16413 18816
rect 16483 18782 16517 18816
rect 17483 18782 17517 18816
rect 17771 18782 17805 18816
rect 18771 18782 18805 18816
rect 18875 18782 18909 18816
rect 19875 18782 19909 18816
rect 19979 18784 20013 18818
rect 20151 18784 20185 18818
rect 4983 18590 5017 18624
rect 5155 18590 5189 18624
rect 5443 18592 5477 18626
rect 6443 18592 6477 18626
rect 6547 18592 6581 18626
rect 7547 18592 7581 18626
rect 7651 18592 7685 18626
rect 8651 18592 8685 18626
rect 8755 18592 8789 18626
rect 9755 18592 9789 18626
rect 10043 18592 10077 18626
rect 10491 18592 10525 18626
rect 10595 18592 10629 18626
rect 11595 18592 11629 18626
rect 11699 18592 11733 18626
rect 12699 18592 12733 18626
rect 12803 18592 12837 18626
rect 13803 18592 13837 18626
rect 13907 18592 13941 18626
rect 14907 18592 14941 18626
rect 15195 18585 15229 18619
rect 15459 18585 15493 18619
rect 15563 18592 15597 18626
rect 16563 18592 16597 18626
rect 16667 18592 16701 18626
rect 17667 18592 17701 18626
rect 17771 18592 17805 18626
rect 18771 18592 18805 18626
rect 18875 18592 18909 18626
rect 19875 18592 19909 18626
rect 19979 18590 20013 18624
rect 20151 18590 20185 18624
rect 4983 17696 5017 17730
rect 5155 17696 5189 17730
rect 5443 17694 5477 17728
rect 6075 17694 6109 17728
rect 6179 17694 6213 17728
rect 7179 17694 7213 17728
rect 7467 17694 7501 17728
rect 7915 17694 7949 17728
rect 8019 17694 8053 17728
rect 9019 17694 9053 17728
rect 9123 17694 9157 17728
rect 10123 17694 10157 17728
rect 10227 17694 10261 17728
rect 11227 17694 11261 17728
rect 11331 17694 11365 17728
rect 12331 17694 12365 17728
rect 12619 17694 12653 17728
rect 13067 17694 13101 17728
rect 13171 17694 13205 17728
rect 14171 17694 14205 17728
rect 14275 17694 14309 17728
rect 15275 17694 15309 17728
rect 15379 17694 15413 17728
rect 16379 17694 16413 17728
rect 16483 17694 16517 17728
rect 17483 17694 17517 17728
rect 17771 17694 17805 17728
rect 18771 17694 18805 17728
rect 18875 17694 18909 17728
rect 19875 17694 19909 17728
rect 19979 17696 20013 17730
rect 20151 17696 20185 17730
rect 4983 17502 5017 17536
rect 5155 17502 5189 17536
rect 5443 17504 5477 17538
rect 6443 17504 6477 17538
rect 6547 17504 6581 17538
rect 7547 17504 7581 17538
rect 7651 17504 7685 17538
rect 8651 17504 8685 17538
rect 8755 17504 8789 17538
rect 9755 17504 9789 17538
rect 10043 17504 10077 17538
rect 10491 17504 10525 17538
rect 10595 17504 10629 17538
rect 11595 17504 11629 17538
rect 11699 17504 11733 17538
rect 12699 17504 12733 17538
rect 12803 17504 12837 17538
rect 13803 17504 13837 17538
rect 13907 17504 13941 17538
rect 14907 17504 14941 17538
rect 15195 17497 15229 17531
rect 15459 17497 15493 17531
rect 15563 17504 15597 17538
rect 16563 17504 16597 17538
rect 16667 17504 16701 17538
rect 17667 17504 17701 17538
rect 17771 17504 17805 17538
rect 18771 17504 18805 17538
rect 18875 17504 18909 17538
rect 19875 17504 19909 17538
rect 19979 17502 20013 17536
rect 20151 17502 20185 17536
rect 4983 16608 5017 16642
rect 5155 16608 5189 16642
rect 5443 16606 5477 16640
rect 6075 16606 6109 16640
rect 6179 16606 6213 16640
rect 7179 16606 7213 16640
rect 7467 16606 7501 16640
rect 7915 16606 7949 16640
rect 8019 16606 8053 16640
rect 9019 16606 9053 16640
rect 9123 16606 9157 16640
rect 10123 16606 10157 16640
rect 10227 16606 10261 16640
rect 11227 16606 11261 16640
rect 11331 16606 11365 16640
rect 12331 16606 12365 16640
rect 12619 16606 12653 16640
rect 13067 16606 13101 16640
rect 13171 16606 13205 16640
rect 14171 16606 14205 16640
rect 14275 16606 14309 16640
rect 15275 16606 15309 16640
rect 15379 16606 15413 16640
rect 16379 16606 16413 16640
rect 16483 16606 16517 16640
rect 17483 16606 17517 16640
rect 17771 16606 17805 16640
rect 18771 16606 18805 16640
rect 18875 16606 18909 16640
rect 19875 16606 19909 16640
rect 19979 16608 20013 16642
rect 20151 16608 20185 16642
rect 4983 16414 5017 16448
rect 5155 16414 5189 16448
rect 5443 16416 5477 16450
rect 6443 16416 6477 16450
rect 6547 16416 6581 16450
rect 7547 16416 7581 16450
rect 7651 16416 7685 16450
rect 8651 16416 8685 16450
rect 8755 16416 8789 16450
rect 9755 16416 9789 16450
rect 10043 16416 10077 16450
rect 10491 16416 10525 16450
rect 10595 16416 10629 16450
rect 11595 16416 11629 16450
rect 11699 16416 11733 16450
rect 12699 16416 12733 16450
rect 12803 16416 12837 16450
rect 13803 16416 13837 16450
rect 13907 16416 13941 16450
rect 14907 16416 14941 16450
rect 15195 16409 15229 16443
rect 15459 16409 15493 16443
rect 15563 16416 15597 16450
rect 16563 16416 16597 16450
rect 16667 16416 16701 16450
rect 17667 16416 17701 16450
rect 17771 16416 17805 16450
rect 18771 16416 18805 16450
rect 18875 16416 18909 16450
rect 19875 16416 19909 16450
rect 19979 16414 20013 16448
rect 20151 16414 20185 16448
rect 4983 15520 5017 15554
rect 5155 15520 5189 15554
rect 5443 15518 5477 15552
rect 6075 15518 6109 15552
rect 6179 15518 6213 15552
rect 7179 15518 7213 15552
rect 7467 15518 7501 15552
rect 7915 15518 7949 15552
rect 8019 15518 8053 15552
rect 9019 15518 9053 15552
rect 9123 15518 9157 15552
rect 10123 15518 10157 15552
rect 10227 15518 10261 15552
rect 11227 15518 11261 15552
rect 11331 15518 11365 15552
rect 12331 15518 12365 15552
rect 12619 15518 12653 15552
rect 13067 15518 13101 15552
rect 13171 15518 13205 15552
rect 14171 15518 14205 15552
rect 14275 15518 14309 15552
rect 15275 15518 15309 15552
rect 15379 15518 15413 15552
rect 16379 15518 16413 15552
rect 16483 15518 16517 15552
rect 17483 15518 17517 15552
rect 17771 15518 17805 15552
rect 18771 15518 18805 15552
rect 18875 15518 18909 15552
rect 19875 15518 19909 15552
rect 19979 15520 20013 15554
rect 20151 15520 20185 15554
rect 4983 15326 5017 15360
rect 5155 15326 5189 15360
rect 5443 15328 5477 15362
rect 6443 15328 6477 15362
rect 6547 15328 6581 15362
rect 7547 15328 7581 15362
rect 7651 15328 7685 15362
rect 8651 15328 8685 15362
rect 8755 15328 8789 15362
rect 9755 15328 9789 15362
rect 10043 15328 10077 15362
rect 10491 15328 10525 15362
rect 10595 15328 10629 15362
rect 11595 15328 11629 15362
rect 11699 15328 11733 15362
rect 12699 15328 12733 15362
rect 12825 15321 12859 15355
rect 12909 15347 12943 15381
rect 13063 15321 13097 15355
rect 13167 15321 13201 15355
rect 13326 15347 13360 15381
rect 13416 15321 13450 15355
rect 13539 15321 13573 15355
rect 13803 15321 13837 15355
rect 13907 15328 13941 15362
rect 14907 15328 14941 15362
rect 15103 15326 15137 15360
rect 15275 15326 15309 15360
rect 15401 15321 15435 15355
rect 15485 15347 15519 15381
rect 15639 15321 15673 15355
rect 15743 15321 15777 15355
rect 15902 15347 15936 15381
rect 15992 15321 16026 15355
rect 16115 15328 16149 15362
rect 16563 15328 16597 15362
rect 16667 15328 16701 15362
rect 17667 15328 17701 15362
rect 17771 15328 17805 15362
rect 18771 15328 18805 15362
rect 18875 15328 18909 15362
rect 19875 15328 19909 15362
rect 19979 15326 20013 15360
rect 20151 15326 20185 15360
rect 4983 14432 5017 14466
rect 5155 14432 5189 14466
rect 5443 14430 5477 14464
rect 6075 14430 6109 14464
rect 6179 14430 6213 14464
rect 7179 14430 7213 14464
rect 7375 14430 7409 14464
rect 8375 14430 8409 14464
rect 8479 14430 8513 14464
rect 9479 14430 9513 14464
rect 9583 14430 9617 14464
rect 10583 14430 10617 14464
rect 10733 14426 10767 14460
rect 10817 14426 10851 14460
rect 10885 14426 10919 14460
rect 11120 14426 11154 14460
rect 11327 14411 11361 14445
rect 11411 14430 11445 14464
rect 11699 14430 11733 14464
rect 12331 14430 12365 14464
rect 12757 14426 12791 14460
rect 12841 14426 12875 14460
rect 12909 14426 12943 14460
rect 13144 14426 13178 14460
rect 13351 14411 13385 14445
rect 13435 14430 13469 14464
rect 13539 14430 13573 14464
rect 14171 14430 14205 14464
rect 14275 14424 14309 14458
rect 14361 14411 14395 14445
rect 14447 14441 14481 14475
rect 14551 14461 14585 14495
rect 14635 14411 14669 14445
rect 14759 14427 14793 14461
rect 14977 14407 15011 14441
rect 15189 14411 15223 14445
rect 15299 14407 15333 14441
rect 15411 14411 15445 14445
rect 15757 14413 15791 14447
rect 15864 14413 15898 14447
rect 15997 14407 16031 14441
rect 16119 14437 16153 14471
rect 16203 14411 16237 14445
rect 16287 14437 16321 14471
rect 16483 14430 16517 14464
rect 17483 14430 17517 14464
rect 17771 14430 17805 14464
rect 18771 14430 18805 14464
rect 18875 14430 18909 14464
rect 19875 14430 19909 14464
rect 19979 14432 20013 14466
rect 20151 14432 20185 14466
rect 4983 14238 5017 14272
rect 5155 14238 5189 14272
rect 5443 14240 5477 14274
rect 6443 14240 6477 14274
rect 6547 14240 6581 14274
rect 7547 14240 7581 14274
rect 7651 14240 7685 14274
rect 8651 14240 8685 14274
rect 8755 14240 8789 14274
rect 9755 14240 9789 14274
rect 10135 14209 10169 14243
rect 10219 14259 10253 14293
rect 10343 14243 10377 14277
rect 10561 14263 10595 14297
rect 10773 14259 10807 14293
rect 10883 14263 10917 14297
rect 10995 14259 11029 14293
rect 11341 14257 11375 14291
rect 11448 14257 11482 14291
rect 11581 14263 11615 14297
rect 11703 14233 11737 14267
rect 11787 14259 11821 14293
rect 11871 14233 11905 14267
rect 11975 14229 12009 14263
rect 12061 14259 12095 14293
rect 12147 14246 12181 14280
rect 12268 14255 12302 14289
rect 12354 14246 12388 14280
rect 12440 14255 12474 14289
rect 12526 14246 12560 14280
rect 12612 14255 12646 14289
rect 12698 14246 12732 14280
rect 12784 14255 12818 14289
rect 12870 14246 12904 14280
rect 12955 14255 12989 14289
rect 13041 14246 13075 14280
rect 13127 14255 13161 14289
rect 13213 14246 13247 14280
rect 13299 14255 13333 14289
rect 13385 14246 13419 14280
rect 13471 14255 13505 14289
rect 13557 14246 13591 14280
rect 13643 14246 13677 14280
rect 13729 14246 13763 14280
rect 13815 14246 13849 14280
rect 13901 14246 13935 14280
rect 13987 14259 14021 14293
rect 14297 14233 14331 14267
rect 14381 14259 14415 14293
rect 14535 14233 14569 14267
rect 14639 14233 14673 14267
rect 14798 14259 14832 14293
rect 14888 14233 14922 14267
rect 15195 14240 15229 14274
rect 15279 14259 15313 14293
rect 15486 14244 15520 14278
rect 15721 14244 15755 14278
rect 15789 14244 15823 14278
rect 15873 14244 15907 14278
rect 16023 14229 16057 14263
rect 16109 14259 16143 14293
rect 16195 14246 16229 14280
rect 16299 14229 16333 14263
rect 16385 14259 16419 14293
rect 16471 14246 16505 14280
rect 16667 14240 16701 14274
rect 17667 14240 17701 14274
rect 17771 14240 17805 14274
rect 18771 14240 18805 14274
rect 18875 14240 18909 14274
rect 19875 14240 19909 14274
rect 19979 14238 20013 14272
rect 20151 14238 20185 14272
rect 4983 13344 5017 13378
rect 5155 13344 5189 13378
rect 5443 13342 5477 13376
rect 6075 13342 6109 13376
rect 6179 13342 6213 13376
rect 7179 13342 7213 13376
rect 7467 13342 7501 13376
rect 8467 13342 8501 13376
rect 8571 13342 8605 13376
rect 9571 13342 9605 13376
rect 9675 13336 9709 13370
rect 9761 13323 9795 13357
rect 9847 13353 9881 13387
rect 9968 13327 10002 13361
rect 10054 13336 10088 13370
rect 10140 13327 10174 13361
rect 10226 13336 10260 13370
rect 10312 13327 10346 13361
rect 10398 13336 10432 13370
rect 10484 13327 10518 13361
rect 10570 13336 10604 13370
rect 10655 13327 10689 13361
rect 10741 13336 10775 13370
rect 10827 13327 10861 13361
rect 10913 13336 10947 13370
rect 10999 13327 11033 13361
rect 11085 13336 11119 13370
rect 11171 13327 11205 13361
rect 11257 13336 11291 13370
rect 11343 13336 11377 13370
rect 11429 13336 11463 13370
rect 11515 13336 11549 13370
rect 11601 13336 11635 13370
rect 11687 13323 11721 13357
rect 11883 13342 11917 13376
rect 12331 13342 12365 13376
rect 12527 13353 12561 13387
rect 12613 13323 12647 13357
rect 12699 13336 12733 13370
rect 12895 13373 12929 13407
rect 12979 13323 13013 13357
rect 13103 13339 13137 13373
rect 13321 13319 13355 13353
rect 13533 13323 13567 13357
rect 13643 13319 13677 13353
rect 13755 13323 13789 13357
rect 14101 13325 14135 13359
rect 14208 13325 14242 13359
rect 14341 13319 14375 13353
rect 14463 13349 14497 13383
rect 14547 13323 14581 13357
rect 14631 13349 14665 13383
rect 14735 13323 14769 13357
rect 14821 13336 14855 13370
rect 14907 13336 14941 13370
rect 14993 13336 15027 13370
rect 15079 13336 15113 13370
rect 15165 13336 15199 13370
rect 15251 13327 15285 13361
rect 15337 13336 15371 13370
rect 15423 13327 15457 13361
rect 15509 13336 15543 13370
rect 15595 13327 15629 13361
rect 15681 13336 15715 13370
rect 15767 13327 15801 13361
rect 15852 13336 15886 13370
rect 15938 13327 15972 13361
rect 16024 13336 16058 13370
rect 16110 13327 16144 13361
rect 16196 13336 16230 13370
rect 16282 13327 16316 13361
rect 16368 13336 16402 13370
rect 16454 13327 16488 13361
rect 16575 13342 16609 13376
rect 16659 13323 16693 13357
rect 16866 13338 16900 13372
rect 17101 13338 17135 13372
rect 17169 13338 17203 13372
rect 17253 13338 17287 13372
rect 17771 13342 17805 13376
rect 18771 13342 18805 13376
rect 18875 13342 18909 13376
rect 19875 13342 19909 13376
rect 19979 13344 20013 13378
rect 20151 13344 20185 13378
rect 4983 13150 5017 13184
rect 5155 13150 5189 13184
rect 5259 13152 5293 13186
rect 5707 13152 5741 13186
rect 5811 13152 5845 13186
rect 6811 13152 6845 13186
rect 6915 13152 6949 13186
rect 7915 13152 7949 13186
rect 8019 13152 8053 13186
rect 9019 13152 9053 13186
rect 9145 13145 9179 13179
rect 9229 13171 9263 13205
rect 9383 13145 9417 13179
rect 9487 13145 9521 13179
rect 9646 13171 9680 13205
rect 9736 13145 9770 13179
rect 10043 13145 10077 13179
rect 10307 13145 10341 13179
rect 10411 13121 10445 13155
rect 10495 13171 10529 13205
rect 10619 13155 10653 13189
rect 10837 13175 10871 13209
rect 11049 13171 11083 13205
rect 11159 13175 11193 13209
rect 11271 13171 11305 13205
rect 11617 13169 11651 13203
rect 11724 13169 11758 13203
rect 11857 13175 11891 13209
rect 11979 13145 12013 13179
rect 12063 13171 12097 13205
rect 12147 13145 12181 13179
rect 12251 13145 12285 13179
rect 12335 13171 12369 13205
rect 12419 13145 12453 13179
rect 12541 13175 12575 13209
rect 12674 13169 12708 13203
rect 12781 13169 12815 13203
rect 13127 13171 13161 13205
rect 13239 13175 13273 13209
rect 13349 13171 13383 13205
rect 13561 13175 13595 13209
rect 13779 13155 13813 13189
rect 13903 13171 13937 13205
rect 13987 13121 14021 13155
rect 14091 13152 14125 13186
rect 14175 13171 14209 13205
rect 14382 13156 14416 13190
rect 14617 13156 14651 13190
rect 14685 13156 14719 13190
rect 14769 13156 14803 13190
rect 15103 13121 15137 13155
rect 15187 13171 15221 13205
rect 15311 13155 15345 13189
rect 15529 13175 15563 13209
rect 15741 13171 15775 13205
rect 15851 13175 15885 13209
rect 15963 13171 15997 13205
rect 16309 13169 16343 13203
rect 16416 13169 16450 13203
rect 16549 13175 16583 13209
rect 16671 13145 16705 13179
rect 16755 13171 16789 13205
rect 16839 13145 16873 13179
rect 16962 13145 16996 13179
rect 17052 13171 17086 13205
rect 17211 13145 17245 13179
rect 17315 13145 17349 13179
rect 17469 13171 17503 13205
rect 17553 13145 17587 13179
rect 17771 13152 17805 13186
rect 18771 13152 18805 13186
rect 18875 13152 18909 13186
rect 19875 13152 19909 13186
rect 19979 13150 20013 13184
rect 20151 13150 20185 13184
rect 4983 12256 5017 12290
rect 5155 12256 5189 12290
rect 5627 12254 5661 12288
rect 6627 12254 6661 12288
rect 6738 12239 6772 12273
rect 6824 12261 6858 12295
rect 6910 12239 6944 12273
rect 6996 12261 7030 12295
rect 7093 12239 7127 12273
rect 7179 12243 7213 12277
rect 7375 12261 7409 12295
rect 7639 12261 7673 12295
rect 7743 12254 7777 12288
rect 8743 12254 8777 12288
rect 8854 12239 8888 12273
rect 8940 12261 8974 12295
rect 9026 12239 9060 12273
rect 9112 12261 9146 12295
rect 9209 12239 9243 12273
rect 9295 12243 9329 12277
rect 9491 12261 9525 12295
rect 9755 12261 9789 12295
rect 9958 12239 9992 12273
rect 10044 12261 10078 12295
rect 10130 12239 10164 12273
rect 10216 12261 10250 12295
rect 10313 12239 10347 12273
rect 10399 12243 10433 12277
rect 10503 12254 10537 12288
rect 10587 12235 10621 12269
rect 10794 12250 10828 12284
rect 11029 12250 11063 12284
rect 11097 12250 11131 12284
rect 11181 12250 11215 12284
rect 11469 12250 11503 12284
rect 11553 12250 11587 12284
rect 11621 12250 11655 12284
rect 11856 12250 11890 12284
rect 12063 12235 12097 12269
rect 12147 12254 12181 12288
rect 12718 12239 12752 12273
rect 12804 12261 12838 12295
rect 12890 12239 12924 12273
rect 12976 12261 13010 12295
rect 13073 12239 13107 12273
rect 13159 12243 13193 12277
rect 13263 12243 13297 12277
rect 13349 12239 13383 12273
rect 13446 12261 13480 12295
rect 13532 12239 13566 12273
rect 13618 12261 13652 12295
rect 13704 12239 13738 12273
rect 13815 12248 13849 12282
rect 13901 12235 13935 12269
rect 13987 12265 14021 12299
rect 14113 12261 14147 12295
rect 14197 12235 14231 12269
rect 14351 12261 14385 12295
rect 14455 12261 14489 12295
rect 14614 12235 14648 12269
rect 14704 12261 14738 12295
rect 15103 12261 15137 12295
rect 15187 12235 15221 12269
rect 15271 12261 15305 12295
rect 15393 12231 15427 12265
rect 15526 12237 15560 12271
rect 15633 12237 15667 12271
rect 15979 12235 16013 12269
rect 16091 12231 16125 12265
rect 16201 12235 16235 12269
rect 16413 12231 16447 12265
rect 16631 12251 16665 12285
rect 16755 12235 16789 12269
rect 16839 12285 16873 12319
rect 17035 12243 17069 12277
rect 17121 12239 17155 12273
rect 17218 12261 17252 12295
rect 17304 12239 17338 12273
rect 17390 12261 17424 12295
rect 17476 12239 17510 12273
rect 17771 12254 17805 12288
rect 18219 12254 18253 12288
rect 18323 12254 18357 12288
rect 19323 12254 19357 12288
rect 19427 12243 19461 12277
rect 19513 12239 19547 12273
rect 19610 12261 19644 12295
rect 19696 12239 19730 12273
rect 19782 12261 19816 12295
rect 19868 12239 19902 12273
rect 19979 12256 20013 12290
rect 20151 12256 20185 12290
rect 29872 4370 29906 4546
rect 30130 4370 30164 4546
rect 30252 4370 30286 4546
rect 30510 4370 30544 4546
rect 30652 4370 30686 4546
rect 30910 4370 30944 4546
rect 31032 4370 31066 4546
rect 31290 4370 31324 4546
rect 31548 4370 31582 4546
rect 31806 4370 31840 4546
rect 32064 4370 32098 4546
rect 32322 4370 32356 4546
rect 32580 4370 32614 4546
rect 32838 4370 32872 4546
rect 33096 4370 33130 4546
rect 33354 4370 33388 4546
rect 33472 4370 33506 4546
rect 33730 4370 33764 4546
rect 1442 1720 1476 2696
rect 1530 1720 1564 2696
rect 1642 2520 1676 2696
rect 1730 2520 1764 2696
rect 1855 1713 1889 2689
rect 1951 1713 1985 2689
rect 2047 1713 2081 2689
rect 2143 1713 2177 2689
rect 2239 1713 2273 2689
rect 2335 1713 2369 2689
rect 2431 1713 2465 2689
rect 2527 1713 2561 2689
rect 2623 1713 2657 2689
rect 2719 1713 2753 2689
rect 2815 1713 2849 2689
rect 2911 1713 2945 2689
rect 3007 1713 3041 2689
rect 3122 1720 3156 2696
rect 3210 1720 3244 2696
rect 4742 1720 4776 2696
rect 4830 1720 4864 2696
rect 4942 2520 4976 2696
rect 5030 2520 5064 2696
rect 5155 1713 5189 2689
rect 5251 1713 5285 2689
rect 5347 1713 5381 2689
rect 5443 1713 5477 2689
rect 5539 1713 5573 2689
rect 5635 1713 5669 2689
rect 5731 1713 5765 2689
rect 5827 1713 5861 2689
rect 5923 1713 5957 2689
rect 6019 1713 6053 2689
rect 6115 1713 6149 2689
rect 6211 1713 6245 2689
rect 6307 1713 6341 2689
rect 6422 1720 6456 2696
rect 6510 1720 6544 2696
rect 8042 1720 8076 2696
rect 8130 1720 8164 2696
rect 8242 2520 8276 2696
rect 8330 2520 8364 2696
rect 8455 1713 8489 2689
rect 8551 1713 8585 2689
rect 8647 1713 8681 2689
rect 8743 1713 8777 2689
rect 8839 1713 8873 2689
rect 8935 1713 8969 2689
rect 9031 1713 9065 2689
rect 9127 1713 9161 2689
rect 9223 1713 9257 2689
rect 9319 1713 9353 2689
rect 9415 1713 9449 2689
rect 9511 1713 9545 2689
rect 9607 1713 9641 2689
rect 9722 1720 9756 2696
rect 9810 1720 9844 2696
rect 11342 1720 11376 2696
rect 11430 1720 11464 2696
rect 11542 2520 11576 2696
rect 11630 2520 11664 2696
rect 11755 1713 11789 2689
rect 11851 1713 11885 2689
rect 11947 1713 11981 2689
rect 12043 1713 12077 2689
rect 12139 1713 12173 2689
rect 12235 1713 12269 2689
rect 12331 1713 12365 2689
rect 12427 1713 12461 2689
rect 12523 1713 12557 2689
rect 12619 1713 12653 2689
rect 12715 1713 12749 2689
rect 12811 1713 12845 2689
rect 12907 1713 12941 2689
rect 13022 1720 13056 2696
rect 13110 1720 13144 2696
rect 14942 1720 14976 2696
rect 15030 1720 15064 2696
rect 15142 2520 15176 2696
rect 15230 2520 15264 2696
rect 15355 1713 15389 2689
rect 15451 1713 15485 2689
rect 15547 1713 15581 2689
rect 15643 1713 15677 2689
rect 15739 1713 15773 2689
rect 15835 1713 15869 2689
rect 15931 1713 15965 2689
rect 16027 1713 16061 2689
rect 16123 1713 16157 2689
rect 16219 1713 16253 2689
rect 16315 1713 16349 2689
rect 16411 1713 16445 2689
rect 16507 1713 16541 2689
rect 16622 1720 16656 2696
rect 16710 1720 16744 2696
rect 18442 1720 18476 2696
rect 18530 1720 18564 2696
rect 18642 2520 18676 2696
rect 18730 2520 18764 2696
rect 18855 1713 18889 2689
rect 18951 1713 18985 2689
rect 19047 1713 19081 2689
rect 19143 1713 19177 2689
rect 19239 1713 19273 2689
rect 19335 1713 19369 2689
rect 19431 1713 19465 2689
rect 19527 1713 19561 2689
rect 19623 1713 19657 2689
rect 19719 1713 19753 2689
rect 19815 1713 19849 2689
rect 19911 1713 19945 2689
rect 20007 1713 20041 2689
rect 20122 1720 20156 2696
rect 20210 1720 20244 2696
rect 22142 1720 22176 2696
rect 22230 1720 22264 2696
rect 22342 2520 22376 2696
rect 22430 2520 22464 2696
rect 22555 1713 22589 2689
rect 22651 1713 22685 2689
rect 22747 1713 22781 2689
rect 22843 1713 22877 2689
rect 22939 1713 22973 2689
rect 23035 1713 23069 2689
rect 23131 1713 23165 2689
rect 23227 1713 23261 2689
rect 23323 1713 23357 2689
rect 23419 1713 23453 2689
rect 23515 1713 23549 2689
rect 23611 1713 23645 2689
rect 23707 1713 23741 2689
rect 23822 1720 23856 2696
rect 23910 1720 23944 2696
rect 25942 1720 25976 2696
rect 26030 1720 26064 2696
rect 26142 2520 26176 2696
rect 26230 2520 26264 2696
rect 26355 1713 26389 2689
rect 26451 1713 26485 2689
rect 26547 1713 26581 2689
rect 26643 1713 26677 2689
rect 26739 1713 26773 2689
rect 26835 1713 26869 2689
rect 26931 1713 26965 2689
rect 27027 1713 27061 2689
rect 27123 1713 27157 2689
rect 27219 1713 27253 2689
rect 27315 1713 27349 2689
rect 27411 1713 27445 2689
rect 27507 1713 27541 2689
rect 27622 1720 27656 2696
rect 27710 1720 27744 2696
<< pdiffc >>
rect 4983 27018 5017 27052
rect 4983 26923 5017 26957
rect 5155 27018 5189 27052
rect 5155 26923 5189 26957
rect 5259 27018 5293 27052
rect 5259 26923 5293 26957
rect 5431 27018 5465 27052
rect 5431 26923 5465 26957
rect 5543 27005 5577 27039
rect 5543 26937 5577 26971
rect 5629 27067 5663 27101
rect 5629 26999 5663 27033
rect 5629 26931 5663 26965
rect 5715 26923 5749 26957
rect 5801 26958 5835 26992
rect 5897 26991 5931 27025
rect 5897 26923 5931 26957
rect 5983 27053 6017 27087
rect 5983 26931 6017 26965
rect 6179 26923 6213 26957
rect 7179 26923 7213 26957
rect 7375 27018 7409 27052
rect 7375 26923 7409 26957
rect 7547 27018 7581 27052
rect 7547 26923 7581 26957
rect 7651 26923 7685 26957
rect 8651 26923 8685 26957
rect 8755 26923 8789 26957
rect 9755 26923 9789 26957
rect 10135 26999 10169 27033
rect 10135 26931 10169 26965
rect 10221 26999 10255 27033
rect 10221 26931 10255 26965
rect 10307 27012 10341 27046
rect 10307 26931 10341 26965
rect 10595 27025 10629 27059
rect 10595 26923 10629 26957
rect 11227 27025 11261 27059
rect 11227 26923 11261 26957
rect 11331 26923 11365 26957
rect 12331 26923 12365 26957
rect 12527 27018 12561 27052
rect 12527 26923 12561 26957
rect 12699 27018 12733 27052
rect 12699 26923 12733 26957
rect 12803 26923 12837 26957
rect 13803 26923 13837 26957
rect 13907 26923 13941 26957
rect 14907 26923 14941 26957
rect 15103 27018 15137 27052
rect 15103 26923 15137 26957
rect 15275 27018 15309 27052
rect 15275 26923 15309 26957
rect 15379 26923 15413 26957
rect 16379 26923 16413 26957
rect 16483 26923 16517 26957
rect 17483 26923 17517 26957
rect 17771 27025 17805 27059
rect 17771 26923 17805 26957
rect 18403 27025 18437 27059
rect 18403 26923 18437 26957
rect 18515 27005 18549 27039
rect 18515 26937 18549 26971
rect 18601 27067 18635 27101
rect 18601 26999 18635 27033
rect 18601 26931 18635 26965
rect 18687 26923 18721 26957
rect 18773 26958 18807 26992
rect 18869 26991 18903 27025
rect 18869 26923 18903 26957
rect 18955 27053 18989 27087
rect 18955 26931 18989 26965
rect 19243 27025 19277 27059
rect 19243 26923 19277 26957
rect 19875 27025 19909 27059
rect 19875 26923 19909 26957
rect 19979 27018 20013 27052
rect 19979 26923 20013 26957
rect 20151 27018 20185 27052
rect 20151 26923 20185 26957
rect 4983 26771 5017 26805
rect 4983 26676 5017 26710
rect 5155 26771 5189 26805
rect 5155 26676 5189 26710
rect 5443 26771 5477 26805
rect 5443 26669 5477 26703
rect 6075 26771 6109 26805
rect 6075 26669 6109 26703
rect 6179 26771 6213 26805
rect 7179 26771 7213 26805
rect 7467 26771 7501 26805
rect 7467 26669 7501 26703
rect 7915 26771 7949 26805
rect 7915 26669 7949 26703
rect 8019 26771 8053 26805
rect 9019 26771 9053 26805
rect 9123 26771 9157 26805
rect 10123 26771 10157 26805
rect 10227 26771 10261 26805
rect 11227 26771 11261 26805
rect 11331 26771 11365 26805
rect 12331 26771 12365 26805
rect 12619 26771 12653 26805
rect 12619 26669 12653 26703
rect 13067 26771 13101 26805
rect 13067 26669 13101 26703
rect 13171 26771 13205 26805
rect 14171 26771 14205 26805
rect 14275 26771 14309 26805
rect 15275 26771 15309 26805
rect 15379 26771 15413 26805
rect 16379 26771 16413 26805
rect 16483 26771 16517 26805
rect 17483 26771 17517 26805
rect 17771 26771 17805 26805
rect 18771 26771 18805 26805
rect 18875 26771 18909 26805
rect 19875 26771 19909 26805
rect 19979 26771 20013 26805
rect 19979 26676 20013 26710
rect 20151 26771 20185 26805
rect 20151 26676 20185 26710
rect 4983 25930 5017 25964
rect 4983 25835 5017 25869
rect 5155 25930 5189 25964
rect 5155 25835 5189 25869
rect 5443 25835 5477 25869
rect 6443 25835 6477 25869
rect 6547 25835 6581 25869
rect 7547 25835 7581 25869
rect 7651 25835 7685 25869
rect 8651 25835 8685 25869
rect 8755 25835 8789 25869
rect 9755 25835 9789 25869
rect 10043 25937 10077 25971
rect 10043 25835 10077 25869
rect 10491 25937 10525 25971
rect 10491 25835 10525 25869
rect 10595 25835 10629 25869
rect 11595 25835 11629 25869
rect 11699 25835 11733 25869
rect 12699 25835 12733 25869
rect 12803 25835 12837 25869
rect 13803 25835 13837 25869
rect 13907 25835 13941 25869
rect 14907 25835 14941 25869
rect 15195 25937 15229 25971
rect 15195 25835 15229 25869
rect 15459 25937 15493 25971
rect 15459 25835 15493 25869
rect 15563 25835 15597 25869
rect 16563 25835 16597 25869
rect 16667 25835 16701 25869
rect 17667 25835 17701 25869
rect 17771 25835 17805 25869
rect 18771 25835 18805 25869
rect 18875 25835 18909 25869
rect 19875 25835 19909 25869
rect 19979 25930 20013 25964
rect 19979 25835 20013 25869
rect 20151 25930 20185 25964
rect 20151 25835 20185 25869
rect 4983 25683 5017 25717
rect 4983 25588 5017 25622
rect 5155 25683 5189 25717
rect 5155 25588 5189 25622
rect 5443 25683 5477 25717
rect 5443 25581 5477 25615
rect 6075 25683 6109 25717
rect 6075 25581 6109 25615
rect 6179 25683 6213 25717
rect 7179 25683 7213 25717
rect 7467 25683 7501 25717
rect 7467 25581 7501 25615
rect 7915 25683 7949 25717
rect 7915 25581 7949 25615
rect 8019 25683 8053 25717
rect 9019 25683 9053 25717
rect 9123 25683 9157 25717
rect 10123 25683 10157 25717
rect 10227 25683 10261 25717
rect 11227 25683 11261 25717
rect 11331 25683 11365 25717
rect 12331 25683 12365 25717
rect 12619 25683 12653 25717
rect 12619 25581 12653 25615
rect 13067 25683 13101 25717
rect 13067 25581 13101 25615
rect 13171 25683 13205 25717
rect 14171 25683 14205 25717
rect 14275 25683 14309 25717
rect 15275 25683 15309 25717
rect 15379 25683 15413 25717
rect 16379 25683 16413 25717
rect 16483 25683 16517 25717
rect 17483 25683 17517 25717
rect 17771 25683 17805 25717
rect 18771 25683 18805 25717
rect 18875 25683 18909 25717
rect 19875 25683 19909 25717
rect 19979 25683 20013 25717
rect 19979 25588 20013 25622
rect 20151 25683 20185 25717
rect 20151 25588 20185 25622
rect 4983 24842 5017 24876
rect 4983 24747 5017 24781
rect 5155 24842 5189 24876
rect 5155 24747 5189 24781
rect 5443 24747 5477 24781
rect 6443 24747 6477 24781
rect 6547 24747 6581 24781
rect 7547 24747 7581 24781
rect 7651 24747 7685 24781
rect 8651 24747 8685 24781
rect 8755 24747 8789 24781
rect 9755 24747 9789 24781
rect 10043 24849 10077 24883
rect 10043 24747 10077 24781
rect 10491 24849 10525 24883
rect 10491 24747 10525 24781
rect 10595 24747 10629 24781
rect 11595 24747 11629 24781
rect 11699 24747 11733 24781
rect 12699 24747 12733 24781
rect 12803 24747 12837 24781
rect 13803 24747 13837 24781
rect 13907 24747 13941 24781
rect 14907 24747 14941 24781
rect 15195 24849 15229 24883
rect 15195 24747 15229 24781
rect 15459 24849 15493 24883
rect 15459 24747 15493 24781
rect 15563 24747 15597 24781
rect 16563 24747 16597 24781
rect 16667 24747 16701 24781
rect 17667 24747 17701 24781
rect 17771 24747 17805 24781
rect 18771 24747 18805 24781
rect 18875 24747 18909 24781
rect 19875 24747 19909 24781
rect 19979 24842 20013 24876
rect 19979 24747 20013 24781
rect 20151 24842 20185 24876
rect 20151 24747 20185 24781
rect 4983 24595 5017 24629
rect 4983 24500 5017 24534
rect 5155 24595 5189 24629
rect 5155 24500 5189 24534
rect 5443 24595 5477 24629
rect 5443 24493 5477 24527
rect 6075 24595 6109 24629
rect 6075 24493 6109 24527
rect 6179 24595 6213 24629
rect 7179 24595 7213 24629
rect 7467 24595 7501 24629
rect 7467 24493 7501 24527
rect 7915 24595 7949 24629
rect 7915 24493 7949 24527
rect 8019 24595 8053 24629
rect 9019 24595 9053 24629
rect 9123 24595 9157 24629
rect 10123 24595 10157 24629
rect 10227 24595 10261 24629
rect 11227 24595 11261 24629
rect 11331 24595 11365 24629
rect 12331 24595 12365 24629
rect 12619 24595 12653 24629
rect 12619 24493 12653 24527
rect 13067 24595 13101 24629
rect 13067 24493 13101 24527
rect 13171 24595 13205 24629
rect 14171 24595 14205 24629
rect 14275 24595 14309 24629
rect 15275 24595 15309 24629
rect 15379 24595 15413 24629
rect 16379 24595 16413 24629
rect 16483 24595 16517 24629
rect 17483 24595 17517 24629
rect 17771 24595 17805 24629
rect 18771 24595 18805 24629
rect 18875 24595 18909 24629
rect 19875 24595 19909 24629
rect 19979 24595 20013 24629
rect 19979 24500 20013 24534
rect 20151 24595 20185 24629
rect 20151 24500 20185 24534
rect 4983 23754 5017 23788
rect 4983 23659 5017 23693
rect 5155 23754 5189 23788
rect 5155 23659 5189 23693
rect 5443 23659 5477 23693
rect 6443 23659 6477 23693
rect 6547 23659 6581 23693
rect 7547 23659 7581 23693
rect 7651 23659 7685 23693
rect 8651 23659 8685 23693
rect 8755 23659 8789 23693
rect 9755 23659 9789 23693
rect 10043 23761 10077 23795
rect 10043 23659 10077 23693
rect 10491 23761 10525 23795
rect 10491 23659 10525 23693
rect 10595 23659 10629 23693
rect 11595 23659 11629 23693
rect 11699 23659 11733 23693
rect 12699 23659 12733 23693
rect 12803 23659 12837 23693
rect 13803 23659 13837 23693
rect 13907 23659 13941 23693
rect 14907 23659 14941 23693
rect 15195 23761 15229 23795
rect 15195 23659 15229 23693
rect 15459 23761 15493 23795
rect 15459 23659 15493 23693
rect 15563 23659 15597 23693
rect 16563 23659 16597 23693
rect 16667 23659 16701 23693
rect 17667 23659 17701 23693
rect 17771 23659 17805 23693
rect 18771 23659 18805 23693
rect 18875 23659 18909 23693
rect 19875 23659 19909 23693
rect 19979 23754 20013 23788
rect 19979 23659 20013 23693
rect 20151 23754 20185 23788
rect 20151 23659 20185 23693
rect 4983 23507 5017 23541
rect 4983 23412 5017 23446
rect 5155 23507 5189 23541
rect 5155 23412 5189 23446
rect 5443 23507 5477 23541
rect 5443 23405 5477 23439
rect 6075 23507 6109 23541
rect 6075 23405 6109 23439
rect 6179 23507 6213 23541
rect 7179 23507 7213 23541
rect 7467 23507 7501 23541
rect 7467 23405 7501 23439
rect 7915 23507 7949 23541
rect 7915 23405 7949 23439
rect 8019 23507 8053 23541
rect 9019 23507 9053 23541
rect 9123 23507 9157 23541
rect 10123 23507 10157 23541
rect 10227 23507 10261 23541
rect 11227 23507 11261 23541
rect 11331 23507 11365 23541
rect 12331 23507 12365 23541
rect 12619 23507 12653 23541
rect 12619 23405 12653 23439
rect 13067 23507 13101 23541
rect 13067 23405 13101 23439
rect 13171 23507 13205 23541
rect 14171 23507 14205 23541
rect 14275 23507 14309 23541
rect 15275 23507 15309 23541
rect 15379 23507 15413 23541
rect 16379 23507 16413 23541
rect 16483 23507 16517 23541
rect 17483 23507 17517 23541
rect 17771 23507 17805 23541
rect 18771 23507 18805 23541
rect 18875 23507 18909 23541
rect 19875 23507 19909 23541
rect 19979 23507 20013 23541
rect 19979 23412 20013 23446
rect 20151 23507 20185 23541
rect 20151 23412 20185 23446
rect 4983 22666 5017 22700
rect 4983 22571 5017 22605
rect 5155 22666 5189 22700
rect 5155 22571 5189 22605
rect 5443 22571 5477 22605
rect 6443 22571 6477 22605
rect 6547 22571 6581 22605
rect 7547 22571 7581 22605
rect 7651 22571 7685 22605
rect 8651 22571 8685 22605
rect 8755 22571 8789 22605
rect 9755 22571 9789 22605
rect 10043 22673 10077 22707
rect 10043 22571 10077 22605
rect 10491 22673 10525 22707
rect 10491 22571 10525 22605
rect 10595 22571 10629 22605
rect 11595 22571 11629 22605
rect 11699 22571 11733 22605
rect 12699 22571 12733 22605
rect 12803 22571 12837 22605
rect 13803 22571 13837 22605
rect 13907 22571 13941 22605
rect 14907 22571 14941 22605
rect 15195 22673 15229 22707
rect 15195 22571 15229 22605
rect 15459 22673 15493 22707
rect 15459 22571 15493 22605
rect 15563 22571 15597 22605
rect 16563 22571 16597 22605
rect 16667 22571 16701 22605
rect 17667 22571 17701 22605
rect 17771 22571 17805 22605
rect 18771 22571 18805 22605
rect 18875 22571 18909 22605
rect 19875 22571 19909 22605
rect 19979 22666 20013 22700
rect 19979 22571 20013 22605
rect 20151 22666 20185 22700
rect 20151 22571 20185 22605
rect 4983 22419 5017 22453
rect 4983 22324 5017 22358
rect 5155 22419 5189 22453
rect 5155 22324 5189 22358
rect 5443 22419 5477 22453
rect 5443 22317 5477 22351
rect 6075 22419 6109 22453
rect 6075 22317 6109 22351
rect 6179 22419 6213 22453
rect 7179 22419 7213 22453
rect 7467 22419 7501 22453
rect 7467 22317 7501 22351
rect 7915 22419 7949 22453
rect 7915 22317 7949 22351
rect 8019 22419 8053 22453
rect 9019 22419 9053 22453
rect 9123 22419 9157 22453
rect 10123 22419 10157 22453
rect 10227 22419 10261 22453
rect 11227 22419 11261 22453
rect 11331 22419 11365 22453
rect 12331 22419 12365 22453
rect 12619 22419 12653 22453
rect 12619 22317 12653 22351
rect 13067 22419 13101 22453
rect 13067 22317 13101 22351
rect 13171 22419 13205 22453
rect 14171 22419 14205 22453
rect 14275 22419 14309 22453
rect 15275 22419 15309 22453
rect 15379 22419 15413 22453
rect 16379 22419 16413 22453
rect 16483 22419 16517 22453
rect 17483 22419 17517 22453
rect 17771 22419 17805 22453
rect 18771 22419 18805 22453
rect 18875 22419 18909 22453
rect 19875 22419 19909 22453
rect 19979 22419 20013 22453
rect 19979 22324 20013 22358
rect 20151 22419 20185 22453
rect 20151 22324 20185 22358
rect 4983 21578 5017 21612
rect 4983 21483 5017 21517
rect 5155 21578 5189 21612
rect 5155 21483 5189 21517
rect 5443 21483 5477 21517
rect 6443 21483 6477 21517
rect 6547 21483 6581 21517
rect 7547 21483 7581 21517
rect 7651 21483 7685 21517
rect 8651 21483 8685 21517
rect 8755 21483 8789 21517
rect 9755 21483 9789 21517
rect 10043 21585 10077 21619
rect 10043 21483 10077 21517
rect 10491 21585 10525 21619
rect 10491 21483 10525 21517
rect 10595 21483 10629 21517
rect 11595 21483 11629 21517
rect 11699 21483 11733 21517
rect 12699 21483 12733 21517
rect 12803 21483 12837 21517
rect 13803 21483 13837 21517
rect 13907 21483 13941 21517
rect 14907 21483 14941 21517
rect 15195 21585 15229 21619
rect 15195 21483 15229 21517
rect 15459 21585 15493 21619
rect 15459 21483 15493 21517
rect 15563 21483 15597 21517
rect 16563 21483 16597 21517
rect 16667 21483 16701 21517
rect 17667 21483 17701 21517
rect 17771 21483 17805 21517
rect 18771 21483 18805 21517
rect 18875 21483 18909 21517
rect 19875 21483 19909 21517
rect 19979 21578 20013 21612
rect 19979 21483 20013 21517
rect 20151 21578 20185 21612
rect 20151 21483 20185 21517
rect 4983 21331 5017 21365
rect 4983 21236 5017 21270
rect 5155 21331 5189 21365
rect 5155 21236 5189 21270
rect 5443 21331 5477 21365
rect 5443 21229 5477 21263
rect 6075 21331 6109 21365
rect 6075 21229 6109 21263
rect 6179 21331 6213 21365
rect 7179 21331 7213 21365
rect 7467 21331 7501 21365
rect 7467 21229 7501 21263
rect 7915 21331 7949 21365
rect 7915 21229 7949 21263
rect 8019 21331 8053 21365
rect 9019 21331 9053 21365
rect 9123 21331 9157 21365
rect 10123 21331 10157 21365
rect 10227 21331 10261 21365
rect 11227 21331 11261 21365
rect 11331 21331 11365 21365
rect 12331 21331 12365 21365
rect 12619 21331 12653 21365
rect 12619 21229 12653 21263
rect 13067 21331 13101 21365
rect 13067 21229 13101 21263
rect 13171 21331 13205 21365
rect 14171 21331 14205 21365
rect 14275 21331 14309 21365
rect 15275 21331 15309 21365
rect 15379 21331 15413 21365
rect 16379 21331 16413 21365
rect 16483 21331 16517 21365
rect 17483 21331 17517 21365
rect 17771 21331 17805 21365
rect 18771 21331 18805 21365
rect 18875 21331 18909 21365
rect 19875 21331 19909 21365
rect 19979 21331 20013 21365
rect 19979 21236 20013 21270
rect 20151 21331 20185 21365
rect 20151 21236 20185 21270
rect 4983 20490 5017 20524
rect 4983 20395 5017 20429
rect 5155 20490 5189 20524
rect 5155 20395 5189 20429
rect 5443 20395 5477 20429
rect 6443 20395 6477 20429
rect 6547 20395 6581 20429
rect 7547 20395 7581 20429
rect 7651 20395 7685 20429
rect 8651 20395 8685 20429
rect 8755 20395 8789 20429
rect 9755 20395 9789 20429
rect 10043 20497 10077 20531
rect 10043 20395 10077 20429
rect 10491 20497 10525 20531
rect 10491 20395 10525 20429
rect 10595 20395 10629 20429
rect 11595 20395 11629 20429
rect 11699 20395 11733 20429
rect 12699 20395 12733 20429
rect 12803 20395 12837 20429
rect 13803 20395 13837 20429
rect 13907 20395 13941 20429
rect 14907 20395 14941 20429
rect 15195 20497 15229 20531
rect 15195 20395 15229 20429
rect 15459 20497 15493 20531
rect 15459 20395 15493 20429
rect 15563 20395 15597 20429
rect 16563 20395 16597 20429
rect 16667 20395 16701 20429
rect 17667 20395 17701 20429
rect 17771 20395 17805 20429
rect 18771 20395 18805 20429
rect 18875 20395 18909 20429
rect 19875 20395 19909 20429
rect 19979 20490 20013 20524
rect 19979 20395 20013 20429
rect 20151 20490 20185 20524
rect 20151 20395 20185 20429
rect 4983 20243 5017 20277
rect 4983 20148 5017 20182
rect 5155 20243 5189 20277
rect 5155 20148 5189 20182
rect 5443 20243 5477 20277
rect 5443 20141 5477 20175
rect 6075 20243 6109 20277
rect 6075 20141 6109 20175
rect 6179 20243 6213 20277
rect 7179 20243 7213 20277
rect 7467 20243 7501 20277
rect 7467 20141 7501 20175
rect 7915 20243 7949 20277
rect 7915 20141 7949 20175
rect 8019 20243 8053 20277
rect 9019 20243 9053 20277
rect 9123 20243 9157 20277
rect 10123 20243 10157 20277
rect 10227 20243 10261 20277
rect 11227 20243 11261 20277
rect 11331 20243 11365 20277
rect 12331 20243 12365 20277
rect 12619 20243 12653 20277
rect 12619 20141 12653 20175
rect 13067 20243 13101 20277
rect 13067 20141 13101 20175
rect 13171 20243 13205 20277
rect 14171 20243 14205 20277
rect 14275 20243 14309 20277
rect 15275 20243 15309 20277
rect 15379 20243 15413 20277
rect 16379 20243 16413 20277
rect 16483 20243 16517 20277
rect 17483 20243 17517 20277
rect 17771 20243 17805 20277
rect 18771 20243 18805 20277
rect 18875 20243 18909 20277
rect 19875 20243 19909 20277
rect 19979 20243 20013 20277
rect 19979 20148 20013 20182
rect 20151 20243 20185 20277
rect 20151 20148 20185 20182
rect 4983 19402 5017 19436
rect 4983 19307 5017 19341
rect 5155 19402 5189 19436
rect 5155 19307 5189 19341
rect 5443 19307 5477 19341
rect 6443 19307 6477 19341
rect 6547 19307 6581 19341
rect 7547 19307 7581 19341
rect 7651 19307 7685 19341
rect 8651 19307 8685 19341
rect 8755 19307 8789 19341
rect 9755 19307 9789 19341
rect 10043 19409 10077 19443
rect 10043 19307 10077 19341
rect 10491 19409 10525 19443
rect 10491 19307 10525 19341
rect 10595 19307 10629 19341
rect 11595 19307 11629 19341
rect 11699 19307 11733 19341
rect 12699 19307 12733 19341
rect 12803 19307 12837 19341
rect 13803 19307 13837 19341
rect 13907 19307 13941 19341
rect 14907 19307 14941 19341
rect 15195 19409 15229 19443
rect 15195 19307 15229 19341
rect 15459 19409 15493 19443
rect 15459 19307 15493 19341
rect 15563 19307 15597 19341
rect 16563 19307 16597 19341
rect 16667 19307 16701 19341
rect 17667 19307 17701 19341
rect 17771 19307 17805 19341
rect 18771 19307 18805 19341
rect 18875 19307 18909 19341
rect 19875 19307 19909 19341
rect 19979 19402 20013 19436
rect 19979 19307 20013 19341
rect 20151 19402 20185 19436
rect 20151 19307 20185 19341
rect 4983 19155 5017 19189
rect 4983 19060 5017 19094
rect 5155 19155 5189 19189
rect 5155 19060 5189 19094
rect 5443 19155 5477 19189
rect 5443 19053 5477 19087
rect 6075 19155 6109 19189
rect 6075 19053 6109 19087
rect 6179 19155 6213 19189
rect 7179 19155 7213 19189
rect 7467 19155 7501 19189
rect 7467 19053 7501 19087
rect 7915 19155 7949 19189
rect 7915 19053 7949 19087
rect 8019 19155 8053 19189
rect 9019 19155 9053 19189
rect 9123 19155 9157 19189
rect 10123 19155 10157 19189
rect 10227 19155 10261 19189
rect 11227 19155 11261 19189
rect 11331 19155 11365 19189
rect 12331 19155 12365 19189
rect 12619 19155 12653 19189
rect 12619 19053 12653 19087
rect 13067 19155 13101 19189
rect 13067 19053 13101 19087
rect 13171 19155 13205 19189
rect 14171 19155 14205 19189
rect 14275 19155 14309 19189
rect 15275 19155 15309 19189
rect 15379 19155 15413 19189
rect 16379 19155 16413 19189
rect 16483 19155 16517 19189
rect 17483 19155 17517 19189
rect 17771 19155 17805 19189
rect 18771 19155 18805 19189
rect 18875 19155 18909 19189
rect 19875 19155 19909 19189
rect 19979 19155 20013 19189
rect 19979 19060 20013 19094
rect 20151 19155 20185 19189
rect 20151 19060 20185 19094
rect 4983 18314 5017 18348
rect 4983 18219 5017 18253
rect 5155 18314 5189 18348
rect 5155 18219 5189 18253
rect 5443 18219 5477 18253
rect 6443 18219 6477 18253
rect 6547 18219 6581 18253
rect 7547 18219 7581 18253
rect 7651 18219 7685 18253
rect 8651 18219 8685 18253
rect 8755 18219 8789 18253
rect 9755 18219 9789 18253
rect 10043 18321 10077 18355
rect 10043 18219 10077 18253
rect 10491 18321 10525 18355
rect 10491 18219 10525 18253
rect 10595 18219 10629 18253
rect 11595 18219 11629 18253
rect 11699 18219 11733 18253
rect 12699 18219 12733 18253
rect 12803 18219 12837 18253
rect 13803 18219 13837 18253
rect 13907 18219 13941 18253
rect 14907 18219 14941 18253
rect 15195 18321 15229 18355
rect 15195 18219 15229 18253
rect 15459 18321 15493 18355
rect 15459 18219 15493 18253
rect 15563 18219 15597 18253
rect 16563 18219 16597 18253
rect 16667 18219 16701 18253
rect 17667 18219 17701 18253
rect 17771 18219 17805 18253
rect 18771 18219 18805 18253
rect 18875 18219 18909 18253
rect 19875 18219 19909 18253
rect 19979 18314 20013 18348
rect 19979 18219 20013 18253
rect 20151 18314 20185 18348
rect 20151 18219 20185 18253
rect 4983 18067 5017 18101
rect 4983 17972 5017 18006
rect 5155 18067 5189 18101
rect 5155 17972 5189 18006
rect 5443 18067 5477 18101
rect 5443 17965 5477 17999
rect 6075 18067 6109 18101
rect 6075 17965 6109 17999
rect 6179 18067 6213 18101
rect 7179 18067 7213 18101
rect 7467 18067 7501 18101
rect 7467 17965 7501 17999
rect 7915 18067 7949 18101
rect 7915 17965 7949 17999
rect 8019 18067 8053 18101
rect 9019 18067 9053 18101
rect 9123 18067 9157 18101
rect 10123 18067 10157 18101
rect 10227 18067 10261 18101
rect 11227 18067 11261 18101
rect 11331 18067 11365 18101
rect 12331 18067 12365 18101
rect 12619 18067 12653 18101
rect 12619 17965 12653 17999
rect 13067 18067 13101 18101
rect 13067 17965 13101 17999
rect 13171 18067 13205 18101
rect 14171 18067 14205 18101
rect 14275 18067 14309 18101
rect 15275 18067 15309 18101
rect 15379 18067 15413 18101
rect 16379 18067 16413 18101
rect 16483 18067 16517 18101
rect 17483 18067 17517 18101
rect 17771 18067 17805 18101
rect 18771 18067 18805 18101
rect 18875 18067 18909 18101
rect 19875 18067 19909 18101
rect 19979 18067 20013 18101
rect 19979 17972 20013 18006
rect 20151 18067 20185 18101
rect 20151 17972 20185 18006
rect 4983 17226 5017 17260
rect 4983 17131 5017 17165
rect 5155 17226 5189 17260
rect 5155 17131 5189 17165
rect 5443 17131 5477 17165
rect 6443 17131 6477 17165
rect 6547 17131 6581 17165
rect 7547 17131 7581 17165
rect 7651 17131 7685 17165
rect 8651 17131 8685 17165
rect 8755 17131 8789 17165
rect 9755 17131 9789 17165
rect 10043 17233 10077 17267
rect 10043 17131 10077 17165
rect 10491 17233 10525 17267
rect 10491 17131 10525 17165
rect 10595 17131 10629 17165
rect 11595 17131 11629 17165
rect 11699 17131 11733 17165
rect 12699 17131 12733 17165
rect 12803 17131 12837 17165
rect 13803 17131 13837 17165
rect 13907 17131 13941 17165
rect 14907 17131 14941 17165
rect 15195 17233 15229 17267
rect 15195 17131 15229 17165
rect 15459 17233 15493 17267
rect 15459 17131 15493 17165
rect 15563 17131 15597 17165
rect 16563 17131 16597 17165
rect 16667 17131 16701 17165
rect 17667 17131 17701 17165
rect 17771 17131 17805 17165
rect 18771 17131 18805 17165
rect 18875 17131 18909 17165
rect 19875 17131 19909 17165
rect 19979 17226 20013 17260
rect 19979 17131 20013 17165
rect 20151 17226 20185 17260
rect 20151 17131 20185 17165
rect 4983 16979 5017 17013
rect 4983 16884 5017 16918
rect 5155 16979 5189 17013
rect 5155 16884 5189 16918
rect 5443 16979 5477 17013
rect 5443 16877 5477 16911
rect 6075 16979 6109 17013
rect 6075 16877 6109 16911
rect 6179 16979 6213 17013
rect 7179 16979 7213 17013
rect 7467 16979 7501 17013
rect 7467 16877 7501 16911
rect 7915 16979 7949 17013
rect 7915 16877 7949 16911
rect 8019 16979 8053 17013
rect 9019 16979 9053 17013
rect 9123 16979 9157 17013
rect 10123 16979 10157 17013
rect 10227 16979 10261 17013
rect 11227 16979 11261 17013
rect 11331 16979 11365 17013
rect 12331 16979 12365 17013
rect 12619 16979 12653 17013
rect 12619 16877 12653 16911
rect 13067 16979 13101 17013
rect 13067 16877 13101 16911
rect 13171 16979 13205 17013
rect 14171 16979 14205 17013
rect 14275 16979 14309 17013
rect 15275 16979 15309 17013
rect 15379 16979 15413 17013
rect 16379 16979 16413 17013
rect 16483 16979 16517 17013
rect 17483 16979 17517 17013
rect 17771 16979 17805 17013
rect 18771 16979 18805 17013
rect 18875 16979 18909 17013
rect 19875 16979 19909 17013
rect 19979 16979 20013 17013
rect 19979 16884 20013 16918
rect 20151 16979 20185 17013
rect 20151 16884 20185 16918
rect 4983 16138 5017 16172
rect 4983 16043 5017 16077
rect 5155 16138 5189 16172
rect 5155 16043 5189 16077
rect 5443 16043 5477 16077
rect 6443 16043 6477 16077
rect 6547 16043 6581 16077
rect 7547 16043 7581 16077
rect 7651 16043 7685 16077
rect 8651 16043 8685 16077
rect 8755 16043 8789 16077
rect 9755 16043 9789 16077
rect 10043 16145 10077 16179
rect 10043 16043 10077 16077
rect 10491 16145 10525 16179
rect 10491 16043 10525 16077
rect 10595 16043 10629 16077
rect 11595 16043 11629 16077
rect 11699 16043 11733 16077
rect 12699 16043 12733 16077
rect 12803 16043 12837 16077
rect 13803 16043 13837 16077
rect 13907 16043 13941 16077
rect 14907 16043 14941 16077
rect 15195 16145 15229 16179
rect 15195 16043 15229 16077
rect 15459 16145 15493 16179
rect 15459 16043 15493 16077
rect 15563 16043 15597 16077
rect 16563 16043 16597 16077
rect 16667 16043 16701 16077
rect 17667 16043 17701 16077
rect 17771 16043 17805 16077
rect 18771 16043 18805 16077
rect 18875 16043 18909 16077
rect 19875 16043 19909 16077
rect 19979 16138 20013 16172
rect 19979 16043 20013 16077
rect 20151 16138 20185 16172
rect 20151 16043 20185 16077
rect 4983 15891 5017 15925
rect 4983 15796 5017 15830
rect 5155 15891 5189 15925
rect 5155 15796 5189 15830
rect 5443 15891 5477 15925
rect 5443 15789 5477 15823
rect 6075 15891 6109 15925
rect 6075 15789 6109 15823
rect 6179 15891 6213 15925
rect 7179 15891 7213 15925
rect 7467 15891 7501 15925
rect 7467 15789 7501 15823
rect 7915 15891 7949 15925
rect 7915 15789 7949 15823
rect 8019 15891 8053 15925
rect 9019 15891 9053 15925
rect 9123 15891 9157 15925
rect 10123 15891 10157 15925
rect 10227 15891 10261 15925
rect 11227 15891 11261 15925
rect 11331 15891 11365 15925
rect 12331 15891 12365 15925
rect 12619 15891 12653 15925
rect 12619 15789 12653 15823
rect 13067 15891 13101 15925
rect 13067 15789 13101 15823
rect 13171 15891 13205 15925
rect 14171 15891 14205 15925
rect 14275 15891 14309 15925
rect 15275 15891 15309 15925
rect 15379 15891 15413 15925
rect 16379 15891 16413 15925
rect 16483 15891 16517 15925
rect 17483 15891 17517 15925
rect 17771 15891 17805 15925
rect 18771 15891 18805 15925
rect 18875 15891 18909 15925
rect 19875 15891 19909 15925
rect 19979 15891 20013 15925
rect 19979 15796 20013 15830
rect 20151 15891 20185 15925
rect 20151 15796 20185 15830
rect 4983 15050 5017 15084
rect 4983 14955 5017 14989
rect 5155 15050 5189 15084
rect 5155 14955 5189 14989
rect 5443 14955 5477 14989
rect 6443 14955 6477 14989
rect 6547 14955 6581 14989
rect 7547 14955 7581 14989
rect 7651 14955 7685 14989
rect 8651 14955 8685 14989
rect 8755 14955 8789 14989
rect 9755 14955 9789 14989
rect 10043 15057 10077 15091
rect 10043 14955 10077 14989
rect 10491 15057 10525 15091
rect 10491 14955 10525 14989
rect 10595 14955 10629 14989
rect 11595 14955 11629 14989
rect 11699 14955 11733 14989
rect 12699 14955 12733 14989
rect 12825 14981 12859 15015
rect 12909 14955 12943 14989
rect 13063 14981 13097 15015
rect 13167 14981 13201 15015
rect 13326 14955 13360 14989
rect 13416 14981 13450 15015
rect 13539 15057 13573 15091
rect 13539 14955 13573 14989
rect 13803 15057 13837 15091
rect 13803 14955 13837 14989
rect 13907 14955 13941 14989
rect 14907 14955 14941 14989
rect 15103 15050 15137 15084
rect 15103 14955 15137 14989
rect 15275 15050 15309 15084
rect 15275 14955 15309 14989
rect 15401 14981 15435 15015
rect 15485 14955 15519 14989
rect 15639 14981 15673 15015
rect 15743 14981 15777 15015
rect 15902 14955 15936 14989
rect 15992 14981 16026 15015
rect 16115 15057 16149 15091
rect 16115 14955 16149 14989
rect 16563 15057 16597 15091
rect 16563 14955 16597 14989
rect 16667 14955 16701 14989
rect 17667 14955 17701 14989
rect 17771 14955 17805 14989
rect 18771 14955 18805 14989
rect 18875 14955 18909 14989
rect 19875 14955 19909 14989
rect 19979 15050 20013 15084
rect 19979 14955 20013 14989
rect 20151 15050 20185 15084
rect 20151 14955 20185 14989
rect 4983 14803 5017 14837
rect 4983 14708 5017 14742
rect 5155 14803 5189 14837
rect 5155 14708 5189 14742
rect 5443 14803 5477 14837
rect 5443 14701 5477 14735
rect 6075 14803 6109 14837
rect 6075 14701 6109 14735
rect 6179 14803 6213 14837
rect 7179 14803 7213 14837
rect 7375 14803 7409 14837
rect 8375 14803 8409 14837
rect 8479 14803 8513 14837
rect 9479 14803 9513 14837
rect 9583 14803 9617 14837
rect 10583 14803 10617 14837
rect 10733 14743 10767 14777
rect 10819 14743 10853 14777
rect 11016 14743 11050 14777
rect 11091 14743 11125 14777
rect 11327 14803 11361 14837
rect 11327 14735 11361 14769
rect 11327 14667 11361 14701
rect 11411 14803 11445 14837
rect 11411 14735 11445 14769
rect 11411 14667 11445 14701
rect 11699 14803 11733 14837
rect 11699 14701 11733 14735
rect 12331 14803 12365 14837
rect 12331 14701 12365 14735
rect 12757 14743 12791 14777
rect 12843 14743 12877 14777
rect 13040 14743 13074 14777
rect 13115 14743 13149 14777
rect 13351 14803 13385 14837
rect 13351 14735 13385 14769
rect 13351 14667 13385 14701
rect 13435 14803 13469 14837
rect 13435 14735 13469 14769
rect 13435 14667 13469 14701
rect 13539 14803 13573 14837
rect 13539 14701 13573 14735
rect 14171 14803 14205 14837
rect 14171 14701 14205 14735
rect 14275 14795 14309 14829
rect 14275 14727 14309 14761
rect 14361 14795 14395 14829
rect 14361 14727 14395 14761
rect 14447 14795 14481 14829
rect 14447 14714 14481 14748
rect 14551 14767 14585 14801
rect 14551 14699 14585 14733
rect 14635 14803 14669 14837
rect 14635 14735 14669 14769
rect 14764 14803 14798 14837
rect 14850 14777 14884 14811
rect 14934 14803 14968 14837
rect 15126 14802 15160 14836
rect 15223 14795 15257 14829
rect 15311 14803 15345 14837
rect 15424 14777 15458 14811
rect 15508 14793 15542 14827
rect 15605 14777 15639 14811
rect 15759 14801 15793 14835
rect 15852 14795 15886 14829
rect 15936 14803 15970 14837
rect 16119 14795 16153 14829
rect 16119 14727 16153 14761
rect 16203 14779 16237 14813
rect 16287 14795 16321 14829
rect 16287 14727 16321 14761
rect 16483 14803 16517 14837
rect 17483 14803 17517 14837
rect 17771 14803 17805 14837
rect 18771 14803 18805 14837
rect 18875 14803 18909 14837
rect 19875 14803 19909 14837
rect 19979 14803 20013 14837
rect 19979 14708 20013 14742
rect 20151 14803 20185 14837
rect 20151 14708 20185 14742
rect 4983 13962 5017 13996
rect 4983 13867 5017 13901
rect 5155 13962 5189 13996
rect 5155 13867 5189 13901
rect 5443 13867 5477 13901
rect 6443 13867 6477 13901
rect 6547 13867 6581 13901
rect 7547 13867 7581 13901
rect 7651 13867 7685 13901
rect 8651 13867 8685 13901
rect 8755 13867 8789 13901
rect 9755 13867 9789 13901
rect 10135 13971 10169 14005
rect 10135 13903 10169 13937
rect 10219 13935 10253 13969
rect 10219 13867 10253 13901
rect 10348 13867 10382 13901
rect 10434 13893 10468 13927
rect 10518 13867 10552 13901
rect 10710 13868 10744 13902
rect 10807 13875 10841 13909
rect 11703 13943 11737 13977
rect 10895 13867 10929 13901
rect 11008 13893 11042 13927
rect 11092 13877 11126 13911
rect 11189 13893 11223 13927
rect 11343 13869 11377 13903
rect 11436 13875 11470 13909
rect 11520 13867 11554 13901
rect 11703 13875 11737 13909
rect 11787 13891 11821 13925
rect 11871 13943 11905 13977
rect 11871 13875 11905 13909
rect 11975 13956 12009 13990
rect 11975 13875 12009 13909
rect 12061 13943 12095 13977
rect 12061 13875 12095 13909
rect 12147 13943 12181 13977
rect 12147 13875 12181 13909
rect 12268 13891 12302 13925
rect 12354 13997 12388 14031
rect 12354 13911 12388 13945
rect 12440 13891 12474 13925
rect 12526 13997 12560 14031
rect 12526 13911 12560 13945
rect 12612 13891 12646 13925
rect 12698 13997 12732 14031
rect 12698 13911 12732 13945
rect 12784 13891 12818 13925
rect 12870 13997 12904 14031
rect 12870 13911 12904 13945
rect 12955 13891 12989 13925
rect 13041 13997 13075 14031
rect 13041 13911 13075 13945
rect 13127 13891 13161 13925
rect 13213 13997 13247 14031
rect 13213 13911 13247 13945
rect 13299 13891 13333 13925
rect 13385 13997 13419 14031
rect 13385 13911 13419 13945
rect 13471 13891 13505 13925
rect 13557 13997 13591 14031
rect 13557 13911 13591 13945
rect 13643 13935 13677 13969
rect 13643 13867 13677 13901
rect 13729 13951 13763 13985
rect 13729 13883 13763 13917
rect 13815 13935 13849 13969
rect 13815 13867 13849 13901
rect 13901 13943 13935 13977
rect 13901 13875 13935 13909
rect 13987 13935 14021 13969
rect 13987 13867 14021 13901
rect 14297 13893 14331 13927
rect 14381 13867 14415 13901
rect 14535 13893 14569 13927
rect 14639 13893 14673 13927
rect 14798 13867 14832 13901
rect 14888 13893 14922 13927
rect 15195 14003 15229 14037
rect 15195 13935 15229 13969
rect 15195 13867 15229 13901
rect 15279 14003 15313 14037
rect 15279 13935 15313 13969
rect 15279 13867 15313 13901
rect 15515 13927 15549 13961
rect 15590 13927 15624 13961
rect 15787 13927 15821 13961
rect 15873 13927 15907 13961
rect 16023 13956 16057 13990
rect 16023 13875 16057 13909
rect 16109 13943 16143 13977
rect 16109 13875 16143 13909
rect 16195 13943 16229 13977
rect 16195 13875 16229 13909
rect 16299 13956 16333 13990
rect 16299 13875 16333 13909
rect 16385 13943 16419 13977
rect 16385 13875 16419 13909
rect 16471 13943 16505 13977
rect 16471 13875 16505 13909
rect 16667 13867 16701 13901
rect 17667 13867 17701 13901
rect 17771 13867 17805 13901
rect 18771 13867 18805 13901
rect 18875 13867 18909 13901
rect 19875 13867 19909 13901
rect 19979 13962 20013 13996
rect 19979 13867 20013 13901
rect 20151 13962 20185 13996
rect 20151 13867 20185 13901
rect 4983 13715 5017 13749
rect 4983 13620 5017 13654
rect 5155 13715 5189 13749
rect 5155 13620 5189 13654
rect 5443 13715 5477 13749
rect 5443 13613 5477 13647
rect 6075 13715 6109 13749
rect 6075 13613 6109 13647
rect 6179 13715 6213 13749
rect 7179 13715 7213 13749
rect 7467 13715 7501 13749
rect 8467 13715 8501 13749
rect 8571 13715 8605 13749
rect 9571 13715 9605 13749
rect 9675 13707 9709 13741
rect 9675 13639 9709 13673
rect 9761 13707 9795 13741
rect 9761 13639 9795 13673
rect 9847 13707 9881 13741
rect 9847 13626 9881 13660
rect 9968 13691 10002 13725
rect 10054 13671 10088 13705
rect 10054 13585 10088 13619
rect 10140 13691 10174 13725
rect 10226 13671 10260 13705
rect 10226 13585 10260 13619
rect 10312 13691 10346 13725
rect 10398 13671 10432 13705
rect 10398 13585 10432 13619
rect 10484 13691 10518 13725
rect 10570 13671 10604 13705
rect 10570 13585 10604 13619
rect 10655 13691 10689 13725
rect 10741 13671 10775 13705
rect 10741 13585 10775 13619
rect 10827 13691 10861 13725
rect 10913 13671 10947 13705
rect 10913 13585 10947 13619
rect 10999 13691 11033 13725
rect 11085 13671 11119 13705
rect 11085 13585 11119 13619
rect 11171 13691 11205 13725
rect 11257 13671 11291 13705
rect 11257 13585 11291 13619
rect 11343 13715 11377 13749
rect 11343 13647 11377 13681
rect 11429 13699 11463 13733
rect 11429 13631 11463 13665
rect 11515 13715 11549 13749
rect 11515 13647 11549 13681
rect 11601 13707 11635 13741
rect 11601 13639 11635 13673
rect 11687 13715 11721 13749
rect 11687 13647 11721 13681
rect 11883 13715 11917 13749
rect 11883 13613 11917 13647
rect 12331 13715 12365 13749
rect 12331 13613 12365 13647
rect 12527 13707 12561 13741
rect 12527 13626 12561 13660
rect 12613 13707 12647 13741
rect 12613 13639 12647 13673
rect 12699 13707 12733 13741
rect 12699 13639 12733 13673
rect 12895 13679 12929 13713
rect 12895 13611 12929 13645
rect 12979 13715 13013 13749
rect 12979 13647 13013 13681
rect 13108 13715 13142 13749
rect 13194 13689 13228 13723
rect 13278 13715 13312 13749
rect 13470 13714 13504 13748
rect 13567 13707 13601 13741
rect 13655 13715 13689 13749
rect 13768 13689 13802 13723
rect 13852 13705 13886 13739
rect 13949 13689 13983 13723
rect 14103 13713 14137 13747
rect 14196 13707 14230 13741
rect 14280 13715 14314 13749
rect 14463 13707 14497 13741
rect 14463 13639 14497 13673
rect 14547 13691 14581 13725
rect 14631 13707 14665 13741
rect 14631 13639 14665 13673
rect 14735 13715 14769 13749
rect 14735 13647 14769 13681
rect 14821 13707 14855 13741
rect 14821 13639 14855 13673
rect 14907 13715 14941 13749
rect 14907 13647 14941 13681
rect 14993 13699 15027 13733
rect 14993 13631 15027 13665
rect 15079 13715 15113 13749
rect 15079 13647 15113 13681
rect 15165 13671 15199 13705
rect 15165 13585 15199 13619
rect 15251 13691 15285 13725
rect 15337 13671 15371 13705
rect 15337 13585 15371 13619
rect 15423 13691 15457 13725
rect 15509 13671 15543 13705
rect 15509 13585 15543 13619
rect 15595 13691 15629 13725
rect 15681 13671 15715 13705
rect 15681 13585 15715 13619
rect 15767 13691 15801 13725
rect 15852 13671 15886 13705
rect 15852 13585 15886 13619
rect 15938 13691 15972 13725
rect 16024 13671 16058 13705
rect 16024 13585 16058 13619
rect 16110 13691 16144 13725
rect 16196 13671 16230 13705
rect 16196 13585 16230 13619
rect 16282 13691 16316 13725
rect 16368 13671 16402 13705
rect 16368 13585 16402 13619
rect 16454 13691 16488 13725
rect 16575 13715 16609 13749
rect 16575 13647 16609 13681
rect 16575 13579 16609 13613
rect 16659 13715 16693 13749
rect 16659 13647 16693 13681
rect 16895 13655 16929 13689
rect 16970 13655 17004 13689
rect 17167 13655 17201 13689
rect 17253 13655 17287 13689
rect 16659 13579 16693 13613
rect 17771 13715 17805 13749
rect 18771 13715 18805 13749
rect 18875 13715 18909 13749
rect 19875 13715 19909 13749
rect 19979 13715 20013 13749
rect 19979 13620 20013 13654
rect 20151 13715 20185 13749
rect 20151 13620 20185 13654
rect 4983 12874 5017 12908
rect 4983 12779 5017 12813
rect 5155 12874 5189 12908
rect 5155 12779 5189 12813
rect 5259 12881 5293 12915
rect 5259 12779 5293 12813
rect 5707 12881 5741 12915
rect 5707 12779 5741 12813
rect 5811 12779 5845 12813
rect 6811 12779 6845 12813
rect 6915 12779 6949 12813
rect 7915 12779 7949 12813
rect 8019 12779 8053 12813
rect 9019 12779 9053 12813
rect 9145 12805 9179 12839
rect 9229 12779 9263 12813
rect 9383 12805 9417 12839
rect 9487 12805 9521 12839
rect 9646 12779 9680 12813
rect 9736 12805 9770 12839
rect 10043 12881 10077 12915
rect 10043 12779 10077 12813
rect 10307 12881 10341 12915
rect 10307 12779 10341 12813
rect 10411 12883 10445 12917
rect 10411 12815 10445 12849
rect 10495 12847 10529 12881
rect 10495 12779 10529 12813
rect 10624 12779 10658 12813
rect 10710 12805 10744 12839
rect 10794 12779 10828 12813
rect 10986 12780 11020 12814
rect 11083 12787 11117 12821
rect 11979 12855 12013 12889
rect 11171 12779 11205 12813
rect 11284 12805 11318 12839
rect 11368 12789 11402 12823
rect 11465 12805 11499 12839
rect 11619 12781 11653 12815
rect 11712 12787 11746 12821
rect 11796 12779 11830 12813
rect 11979 12787 12013 12821
rect 12063 12803 12097 12837
rect 12147 12855 12181 12889
rect 12147 12787 12181 12821
rect 12251 12855 12285 12889
rect 12251 12787 12285 12821
rect 12335 12803 12369 12837
rect 12419 12855 12453 12889
rect 12419 12787 12453 12821
rect 12602 12779 12636 12813
rect 12686 12787 12720 12821
rect 12779 12781 12813 12815
rect 12933 12805 12967 12839
rect 13030 12789 13064 12823
rect 13114 12805 13148 12839
rect 13227 12779 13261 12813
rect 13315 12787 13349 12821
rect 13412 12780 13446 12814
rect 13604 12779 13638 12813
rect 13688 12805 13722 12839
rect 13774 12779 13808 12813
rect 13903 12847 13937 12881
rect 13903 12779 13937 12813
rect 13987 12883 14021 12917
rect 13987 12815 14021 12849
rect 14091 12915 14125 12949
rect 14091 12847 14125 12881
rect 14091 12779 14125 12813
rect 14175 12915 14209 12949
rect 14175 12847 14209 12881
rect 14175 12779 14209 12813
rect 14411 12839 14445 12873
rect 14486 12839 14520 12873
rect 14683 12839 14717 12873
rect 14769 12839 14803 12873
rect 15103 12883 15137 12917
rect 15103 12815 15137 12849
rect 15187 12847 15221 12881
rect 15187 12779 15221 12813
rect 15316 12779 15350 12813
rect 15402 12805 15436 12839
rect 15486 12779 15520 12813
rect 15678 12780 15712 12814
rect 15775 12787 15809 12821
rect 16671 12855 16705 12889
rect 15863 12779 15897 12813
rect 15976 12805 16010 12839
rect 16060 12789 16094 12823
rect 16157 12805 16191 12839
rect 16311 12781 16345 12815
rect 16404 12787 16438 12821
rect 16488 12779 16522 12813
rect 16671 12787 16705 12821
rect 16755 12803 16789 12837
rect 16839 12855 16873 12889
rect 16839 12787 16873 12821
rect 16962 12805 16996 12839
rect 17052 12779 17086 12813
rect 17211 12805 17245 12839
rect 17315 12805 17349 12839
rect 17469 12779 17503 12813
rect 17553 12805 17587 12839
rect 17771 12779 17805 12813
rect 18771 12779 18805 12813
rect 18875 12779 18909 12813
rect 19875 12779 19909 12813
rect 19979 12874 20013 12908
rect 19979 12779 20013 12813
rect 20151 12874 20185 12908
rect 20151 12779 20185 12813
rect 4983 12627 5017 12661
rect 4983 12532 5017 12566
rect 5155 12627 5189 12661
rect 5155 12532 5189 12566
rect 5627 12627 5661 12661
rect 6627 12627 6661 12661
rect 6739 12613 6773 12647
rect 6739 12545 6773 12579
rect 6825 12619 6859 12653
rect 6825 12551 6859 12585
rect 6825 12483 6859 12517
rect 6911 12627 6945 12661
rect 6997 12592 7031 12626
rect 7093 12627 7127 12661
rect 7093 12559 7127 12593
rect 7179 12619 7213 12653
rect 7179 12497 7213 12531
rect 7375 12627 7409 12661
rect 7375 12525 7409 12559
rect 7639 12627 7673 12661
rect 7639 12525 7673 12559
rect 7743 12627 7777 12661
rect 8743 12627 8777 12661
rect 8855 12613 8889 12647
rect 8855 12545 8889 12579
rect 8941 12619 8975 12653
rect 8941 12551 8975 12585
rect 8941 12483 8975 12517
rect 9027 12627 9061 12661
rect 9113 12592 9147 12626
rect 9209 12627 9243 12661
rect 9209 12559 9243 12593
rect 9295 12619 9329 12653
rect 9295 12497 9329 12531
rect 9491 12627 9525 12661
rect 9491 12525 9525 12559
rect 9755 12627 9789 12661
rect 9755 12525 9789 12559
rect 9959 12613 9993 12647
rect 9959 12545 9993 12579
rect 10045 12619 10079 12653
rect 10045 12551 10079 12585
rect 10045 12483 10079 12517
rect 10131 12627 10165 12661
rect 10217 12592 10251 12626
rect 10313 12627 10347 12661
rect 10313 12559 10347 12593
rect 10399 12619 10433 12653
rect 10399 12497 10433 12531
rect 10503 12627 10537 12661
rect 10503 12559 10537 12593
rect 10503 12491 10537 12525
rect 10587 12627 10621 12661
rect 10587 12559 10621 12593
rect 10823 12567 10857 12601
rect 10898 12567 10932 12601
rect 11095 12567 11129 12601
rect 11181 12567 11215 12601
rect 11469 12567 11503 12601
rect 11555 12567 11589 12601
rect 11752 12567 11786 12601
rect 11827 12567 11861 12601
rect 12063 12627 12097 12661
rect 12063 12559 12097 12593
rect 10587 12491 10621 12525
rect 12063 12491 12097 12525
rect 12147 12627 12181 12661
rect 12147 12559 12181 12593
rect 12147 12491 12181 12525
rect 12719 12613 12753 12647
rect 12719 12545 12753 12579
rect 12805 12619 12839 12653
rect 12805 12551 12839 12585
rect 12805 12483 12839 12517
rect 12891 12627 12925 12661
rect 12977 12592 13011 12626
rect 13073 12627 13107 12661
rect 13073 12559 13107 12593
rect 13159 12619 13193 12653
rect 13159 12497 13193 12531
rect 13263 12619 13297 12653
rect 13263 12497 13297 12531
rect 13349 12627 13383 12661
rect 13349 12559 13383 12593
rect 13445 12592 13479 12626
rect 13531 12627 13565 12661
rect 13617 12619 13651 12653
rect 13617 12551 13651 12585
rect 13617 12483 13651 12517
rect 13703 12613 13737 12647
rect 13703 12545 13737 12579
rect 13815 12619 13849 12653
rect 13815 12551 13849 12585
rect 13901 12619 13935 12653
rect 13901 12551 13935 12585
rect 13987 12619 14021 12653
rect 14113 12601 14147 12635
rect 14197 12627 14231 12661
rect 14351 12601 14385 12635
rect 14455 12601 14489 12635
rect 14614 12627 14648 12661
rect 13987 12538 14021 12572
rect 14704 12601 14738 12635
rect 15103 12619 15137 12653
rect 15103 12551 15137 12585
rect 15187 12603 15221 12637
rect 15271 12619 15305 12653
rect 15454 12627 15488 12661
rect 15538 12619 15572 12653
rect 15631 12625 15665 12659
rect 15785 12601 15819 12635
rect 15882 12617 15916 12651
rect 15966 12601 16000 12635
rect 16079 12627 16113 12661
rect 15271 12551 15305 12585
rect 16167 12619 16201 12653
rect 16264 12626 16298 12660
rect 16456 12627 16490 12661
rect 16540 12601 16574 12635
rect 16626 12627 16660 12661
rect 16755 12627 16789 12661
rect 16755 12559 16789 12593
rect 16839 12591 16873 12625
rect 16839 12523 16873 12557
rect 17035 12619 17069 12653
rect 17035 12497 17069 12531
rect 17121 12627 17155 12661
rect 17121 12559 17155 12593
rect 17217 12592 17251 12626
rect 17303 12627 17337 12661
rect 17389 12619 17423 12653
rect 17389 12551 17423 12585
rect 17389 12483 17423 12517
rect 17475 12613 17509 12647
rect 17475 12545 17509 12579
rect 17771 12627 17805 12661
rect 17771 12525 17805 12559
rect 18219 12627 18253 12661
rect 18219 12525 18253 12559
rect 18323 12627 18357 12661
rect 19323 12627 19357 12661
rect 19427 12619 19461 12653
rect 19427 12497 19461 12531
rect 19513 12627 19547 12661
rect 19513 12559 19547 12593
rect 19609 12592 19643 12626
rect 19695 12627 19729 12661
rect 19781 12619 19815 12653
rect 19781 12551 19815 12585
rect 19781 12483 19815 12517
rect 19867 12613 19901 12647
rect 19867 12545 19901 12579
rect 19979 12627 20013 12661
rect 19979 12532 20013 12566
rect 20151 12627 20185 12661
rect 20151 12532 20185 12566
rect 29768 6162 29802 6738
rect 30026 6162 30060 6738
rect 30148 6162 30182 6738
rect 30406 6162 30440 6738
rect 30664 6162 30698 6738
rect 30788 6162 30822 6738
rect 31046 6162 31080 6738
rect 31304 6162 31338 6738
rect 31562 6162 31596 6738
rect 31688 6162 31722 6738
rect 31946 6162 31980 6738
rect 32204 6162 32238 6738
rect 32462 6162 32496 6738
rect 32720 6162 32754 6738
rect 32978 6162 33012 6738
rect 33236 6162 33270 6738
rect 33494 6162 33528 6738
rect 33752 6162 33786 6738
rect 34010 6162 34044 6738
rect 34268 6162 34302 6738
rect 34388 6162 34422 6738
rect 34646 6162 34680 6738
rect 30028 5142 30062 5718
rect 30116 5142 30150 5718
rect 30248 5142 30282 5718
rect 30344 5142 30378 5718
rect 30440 5142 30474 5718
rect 30536 5142 30570 5718
rect 30648 5142 30682 5718
rect 30744 5142 30778 5718
rect 30840 5142 30874 5718
rect 30936 5142 30970 5718
rect 31048 5142 31082 5718
rect 31136 5142 31170 5718
rect 1438 3242 1472 4218
rect 1526 3242 1560 4218
rect 1638 3242 1672 3818
rect 1726 3242 1760 3818
rect 1851 3235 1885 4211
rect 1947 3235 1981 4211
rect 2043 3235 2077 4211
rect 2139 3235 2173 4211
rect 2235 3235 2269 4211
rect 2331 3235 2365 4211
rect 2427 3235 2461 4211
rect 2523 3235 2557 4211
rect 2619 3235 2653 4211
rect 2715 3235 2749 4211
rect 2811 3235 2845 4211
rect 2907 3235 2941 4211
rect 3003 3235 3037 4211
rect 3138 3242 3172 4218
rect 3226 3242 3260 4218
rect 4738 3242 4772 4218
rect 4826 3242 4860 4218
rect 4938 3242 4972 3818
rect 5026 3242 5060 3818
rect 5151 3235 5185 4211
rect 5247 3235 5281 4211
rect 5343 3235 5377 4211
rect 5439 3235 5473 4211
rect 5535 3235 5569 4211
rect 5631 3235 5665 4211
rect 5727 3235 5761 4211
rect 5823 3235 5857 4211
rect 5919 3235 5953 4211
rect 6015 3235 6049 4211
rect 6111 3235 6145 4211
rect 6207 3235 6241 4211
rect 6303 3235 6337 4211
rect 6438 3242 6472 4218
rect 6526 3242 6560 4218
rect 8038 3242 8072 4218
rect 8126 3242 8160 4218
rect 8238 3242 8272 3818
rect 8326 3242 8360 3818
rect 8451 3235 8485 4211
rect 8547 3235 8581 4211
rect 8643 3235 8677 4211
rect 8739 3235 8773 4211
rect 8835 3235 8869 4211
rect 8931 3235 8965 4211
rect 9027 3235 9061 4211
rect 9123 3235 9157 4211
rect 9219 3235 9253 4211
rect 9315 3235 9349 4211
rect 9411 3235 9445 4211
rect 9507 3235 9541 4211
rect 9603 3235 9637 4211
rect 9738 3242 9772 4218
rect 9826 3242 9860 4218
rect 11338 3242 11372 4218
rect 11426 3242 11460 4218
rect 11538 3242 11572 3818
rect 11626 3242 11660 3818
rect 11751 3235 11785 4211
rect 11847 3235 11881 4211
rect 11943 3235 11977 4211
rect 12039 3235 12073 4211
rect 12135 3235 12169 4211
rect 12231 3235 12265 4211
rect 12327 3235 12361 4211
rect 12423 3235 12457 4211
rect 12519 3235 12553 4211
rect 12615 3235 12649 4211
rect 12711 3235 12745 4211
rect 12807 3235 12841 4211
rect 12903 3235 12937 4211
rect 13038 3242 13072 4218
rect 13126 3242 13160 4218
rect 14938 3242 14972 4218
rect 15026 3242 15060 4218
rect 15138 3242 15172 3818
rect 15226 3242 15260 3818
rect 15351 3235 15385 4211
rect 15447 3235 15481 4211
rect 15543 3235 15577 4211
rect 15639 3235 15673 4211
rect 15735 3235 15769 4211
rect 15831 3235 15865 4211
rect 15927 3235 15961 4211
rect 16023 3235 16057 4211
rect 16119 3235 16153 4211
rect 16215 3235 16249 4211
rect 16311 3235 16345 4211
rect 16407 3235 16441 4211
rect 16503 3235 16537 4211
rect 16638 3242 16672 4218
rect 16726 3242 16760 4218
rect 18438 3242 18472 4218
rect 18526 3242 18560 4218
rect 18638 3242 18672 3818
rect 18726 3242 18760 3818
rect 18851 3235 18885 4211
rect 18947 3235 18981 4211
rect 19043 3235 19077 4211
rect 19139 3235 19173 4211
rect 19235 3235 19269 4211
rect 19331 3235 19365 4211
rect 19427 3235 19461 4211
rect 19523 3235 19557 4211
rect 19619 3235 19653 4211
rect 19715 3235 19749 4211
rect 19811 3235 19845 4211
rect 19907 3235 19941 4211
rect 20003 3235 20037 4211
rect 20138 3242 20172 4218
rect 20226 3242 20260 4218
rect 22138 3242 22172 4218
rect 22226 3242 22260 4218
rect 22338 3242 22372 3818
rect 22426 3242 22460 3818
rect 22551 3235 22585 4211
rect 22647 3235 22681 4211
rect 22743 3235 22777 4211
rect 22839 3235 22873 4211
rect 22935 3235 22969 4211
rect 23031 3235 23065 4211
rect 23127 3235 23161 4211
rect 23223 3235 23257 4211
rect 23319 3235 23353 4211
rect 23415 3235 23449 4211
rect 23511 3235 23545 4211
rect 23607 3235 23641 4211
rect 23703 3235 23737 4211
rect 23838 3242 23872 4218
rect 23926 3242 23960 4218
rect 25938 3242 25972 4218
rect 26026 3242 26060 4218
rect 26138 3242 26172 3818
rect 26226 3242 26260 3818
rect 26351 3235 26385 4211
rect 26447 3235 26481 4211
rect 26543 3235 26577 4211
rect 26639 3235 26673 4211
rect 26735 3235 26769 4211
rect 26831 3235 26865 4211
rect 26927 3235 26961 4211
rect 27023 3235 27057 4211
rect 27119 3235 27153 4211
rect 27215 3235 27249 4211
rect 27311 3235 27345 4211
rect 27407 3235 27441 4211
rect 27503 3235 27537 4211
rect 27638 3242 27672 4218
rect 27726 3242 27760 4218
<< psubdiff >>
rect 7277 27297 7311 27344
rect 7277 27239 7311 27263
rect 9853 27297 9887 27344
rect 9853 27239 9887 27263
rect 12429 27297 12463 27344
rect 12429 27239 12463 27263
rect 15005 27297 15039 27344
rect 15005 27239 15039 27263
rect 17581 27297 17615 27344
rect 17581 27239 17615 27263
rect 7277 26465 7311 26489
rect 7277 26384 7311 26431
rect 12429 26465 12463 26489
rect 12429 26384 12463 26431
rect 17581 26465 17615 26489
rect 17581 26384 17615 26431
rect 9853 26209 9887 26256
rect 9853 26151 9887 26175
rect 15005 26209 15039 26256
rect 15005 26151 15039 26175
rect 7277 25377 7311 25401
rect 7277 25296 7311 25343
rect 12429 25377 12463 25401
rect 12429 25296 12463 25343
rect 17581 25377 17615 25401
rect 17581 25296 17615 25343
rect 9853 25121 9887 25168
rect 9853 25063 9887 25087
rect 15005 25121 15039 25168
rect 15005 25063 15039 25087
rect 7277 24289 7311 24313
rect 7277 24208 7311 24255
rect 12429 24289 12463 24313
rect 12429 24208 12463 24255
rect 17581 24289 17615 24313
rect 17581 24208 17615 24255
rect 9853 24033 9887 24080
rect 9853 23975 9887 23999
rect 15005 24033 15039 24080
rect 15005 23975 15039 23999
rect 7277 23201 7311 23225
rect 7277 23120 7311 23167
rect 12429 23201 12463 23225
rect 12429 23120 12463 23167
rect 17581 23201 17615 23225
rect 17581 23120 17615 23167
rect 9853 22945 9887 22992
rect 9853 22887 9887 22911
rect 15005 22945 15039 22992
rect 15005 22887 15039 22911
rect 7277 22113 7311 22137
rect 7277 22032 7311 22079
rect 12429 22113 12463 22137
rect 12429 22032 12463 22079
rect 17581 22113 17615 22137
rect 17581 22032 17615 22079
rect 9853 21857 9887 21904
rect 9853 21799 9887 21823
rect 15005 21857 15039 21904
rect 15005 21799 15039 21823
rect 7277 21025 7311 21049
rect 7277 20944 7311 20991
rect 12429 21025 12463 21049
rect 12429 20944 12463 20991
rect 17581 21025 17615 21049
rect 17581 20944 17615 20991
rect 9853 20769 9887 20816
rect 9853 20711 9887 20735
rect 15005 20769 15039 20816
rect 15005 20711 15039 20735
rect 7277 19937 7311 19961
rect 7277 19856 7311 19903
rect 12429 19937 12463 19961
rect 12429 19856 12463 19903
rect 17581 19937 17615 19961
rect 17581 19856 17615 19903
rect 9853 19681 9887 19728
rect 9853 19623 9887 19647
rect 15005 19681 15039 19728
rect 15005 19623 15039 19647
rect 7277 18849 7311 18873
rect 7277 18768 7311 18815
rect 12429 18849 12463 18873
rect 12429 18768 12463 18815
rect 17581 18849 17615 18873
rect 17581 18768 17615 18815
rect 9853 18593 9887 18640
rect 9853 18535 9887 18559
rect 15005 18593 15039 18640
rect 15005 18535 15039 18559
rect 7277 17761 7311 17785
rect 7277 17680 7311 17727
rect 12429 17761 12463 17785
rect 12429 17680 12463 17727
rect 17581 17761 17615 17785
rect 17581 17680 17615 17727
rect 9853 17505 9887 17552
rect 9853 17447 9887 17471
rect 15005 17505 15039 17552
rect 15005 17447 15039 17471
rect 7277 16673 7311 16697
rect 7277 16592 7311 16639
rect 12429 16673 12463 16697
rect 12429 16592 12463 16639
rect 17581 16673 17615 16697
rect 17581 16592 17615 16639
rect 9853 16417 9887 16464
rect 9853 16359 9887 16383
rect 15005 16417 15039 16464
rect 15005 16359 15039 16383
rect 7277 15585 7311 15609
rect 7277 15504 7311 15551
rect 12429 15585 12463 15609
rect 12429 15504 12463 15551
rect 17581 15585 17615 15609
rect 17581 15504 17615 15551
rect 9853 15329 9887 15376
rect 9853 15271 9887 15295
rect 15005 15329 15039 15376
rect 15005 15271 15039 15295
rect 7277 14497 7311 14521
rect 7277 14416 7311 14463
rect 12429 14497 12463 14521
rect 12429 14416 12463 14463
rect 17581 14497 17615 14521
rect 17581 14416 17615 14463
rect 9853 14241 9887 14288
rect 9853 14183 9887 14207
rect 15005 14241 15039 14288
rect 15005 14183 15039 14207
rect 7277 13409 7311 13433
rect 7277 13328 7311 13375
rect 12429 13409 12463 13433
rect 12429 13328 12463 13375
rect 17581 13409 17615 13433
rect 17581 13328 17615 13375
rect 9853 13153 9887 13200
rect 9853 13095 9887 13119
rect 15005 13153 15039 13200
rect 15005 13095 15039 13119
rect 7277 12321 7311 12345
rect 7277 12240 7311 12287
rect 9853 12321 9887 12345
rect 9853 12240 9887 12287
rect 12429 12321 12463 12345
rect 12429 12240 12463 12287
rect 15005 12321 15039 12345
rect 15005 12240 15039 12287
rect 17581 12321 17615 12345
rect 17581 12240 17615 12287
rect 25716 9190 25812 9224
rect 28176 9190 28272 9224
rect 25716 9128 25750 9190
rect 28238 9128 28272 9190
rect 25716 7050 25750 7112
rect 28238 7050 28272 7112
rect 25716 7016 25812 7050
rect 28176 7016 28272 7050
rect 16886 6850 16982 6884
rect 17120 6850 17216 6884
rect 16886 6788 16920 6850
rect 13286 6290 13382 6324
rect 13520 6290 13616 6324
rect 13286 6228 13320 6290
rect 9986 6010 10082 6044
rect 10220 6010 10316 6044
rect 3386 5966 3482 6000
rect 3620 5966 3716 6000
rect 3386 5904 3420 5966
rect 3682 5904 3716 5966
rect 9986 5948 10020 6010
rect 3386 4710 3420 4772
rect 3682 4710 3716 4772
rect 3386 4676 3482 4710
rect 3620 4676 3716 4710
rect 6686 5870 6782 5904
rect 6920 5870 7016 5904
rect 6686 5808 6720 5870
rect 6982 5808 7016 5870
rect 6686 4710 6720 4772
rect 6982 4710 7016 4772
rect 6686 4676 6782 4710
rect 6920 4676 7016 4710
rect 10282 5948 10316 6010
rect 9986 4710 10020 4772
rect 10282 4710 10316 4772
rect 9986 4676 10082 4710
rect 10220 4676 10316 4710
rect 13582 6228 13616 6290
rect 13286 4710 13320 4772
rect 13582 4710 13616 4772
rect 13286 4676 13382 4710
rect 13520 4676 13616 4710
rect 17182 6788 17216 6850
rect 16886 4710 16920 4772
rect 17182 4710 17216 4772
rect 16886 4676 16982 4710
rect 17120 4676 17216 4710
rect 20086 6850 20182 6884
rect 20638 6850 20734 6884
rect 20086 6788 20120 6850
rect 20700 6788 20734 6850
rect 20086 4710 20120 4772
rect 20700 4710 20734 4772
rect 20086 4676 20182 4710
rect 20638 4676 20734 4710
rect 23186 6850 23282 6884
rect 24374 6850 24470 6884
rect 23186 6788 23220 6850
rect 24436 6788 24470 6850
rect 23186 4710 23220 4772
rect 24436 4710 24470 4772
rect 23186 4676 23282 4710
rect 24374 4676 24470 4710
rect 25686 6850 25782 6884
rect 28146 6850 28242 6884
rect 25686 6788 25720 6850
rect 28208 6788 28242 6850
rect 25686 4710 25720 4772
rect 28208 4710 28242 4772
rect 25686 4676 25782 4710
rect 28146 4676 28242 4710
rect 29560 4810 34800 4830
rect 29560 4770 29660 4810
rect 34700 4790 34800 4810
rect 34700 4770 34740 4790
rect 29560 4750 34740 4770
rect 29560 4110 29580 4750
rect 29620 4110 29640 4750
rect 34720 4130 34740 4750
rect 34780 4130 34800 4790
rect 34720 4110 34800 4130
rect 29560 4090 34800 4110
rect 29560 4050 29660 4090
rect 34720 4050 34800 4090
rect 29560 4030 34800 4050
rect 1280 2900 3410 2930
rect 440 2690 620 2714
rect 440 2486 620 2510
rect 1280 1520 1310 2900
rect 1350 2860 1390 2900
rect 3310 2890 3410 2900
rect 3310 2860 3350 2890
rect 1350 2840 3350 2860
rect 1350 1570 1370 2840
rect 3330 1570 3350 2840
rect 1350 1540 3350 1570
rect 1350 1520 1390 1540
rect 1280 1500 1390 1520
rect 3310 1510 3350 1540
rect 3390 1510 3410 2890
rect 3310 1500 3410 1510
rect 1280 1480 3410 1500
rect 4580 2900 6710 2930
rect 4580 1520 4610 2900
rect 4650 2860 4690 2900
rect 6610 2890 6710 2900
rect 6610 2860 6650 2890
rect 4650 2840 6650 2860
rect 4650 1570 4670 2840
rect 6630 1570 6650 2840
rect 4650 1540 6650 1570
rect 4650 1520 4690 1540
rect 4580 1500 4690 1520
rect 6610 1510 6650 1540
rect 6690 1510 6710 2890
rect 6610 1500 6710 1510
rect 4580 1480 6710 1500
rect 7880 2900 10010 2930
rect 7880 1520 7910 2900
rect 7950 2860 7990 2900
rect 9910 2890 10010 2900
rect 9910 2860 9950 2890
rect 7950 2840 9950 2860
rect 7950 1570 7970 2840
rect 9930 1570 9950 2840
rect 7950 1540 9950 1570
rect 7950 1520 7990 1540
rect 7880 1500 7990 1520
rect 9910 1510 9950 1540
rect 9990 1510 10010 2890
rect 9910 1500 10010 1510
rect 7880 1480 10010 1500
rect 11180 2900 13310 2930
rect 11180 1520 11210 2900
rect 11250 2860 11290 2900
rect 13210 2890 13310 2900
rect 13210 2860 13250 2890
rect 11250 2840 13250 2860
rect 11250 1570 11270 2840
rect 13230 1570 13250 2840
rect 11250 1540 13250 1570
rect 11250 1520 11290 1540
rect 11180 1500 11290 1520
rect 13210 1510 13250 1540
rect 13290 1510 13310 2890
rect 13210 1500 13310 1510
rect 11180 1480 13310 1500
rect 14780 2900 16910 2930
rect 14780 1520 14810 2900
rect 14850 2860 14890 2900
rect 16810 2890 16910 2900
rect 16810 2860 16850 2890
rect 14850 2840 16850 2860
rect 14850 1570 14870 2840
rect 16830 1570 16850 2840
rect 14850 1540 16850 1570
rect 14850 1520 14890 1540
rect 14780 1500 14890 1520
rect 16810 1510 16850 1540
rect 16890 1510 16910 2890
rect 16810 1500 16910 1510
rect 14780 1480 16910 1500
rect 18280 2900 20410 2930
rect 18280 1520 18310 2900
rect 18350 2860 18390 2900
rect 20310 2890 20410 2900
rect 20310 2860 20350 2890
rect 18350 2840 20350 2860
rect 18350 1570 18370 2840
rect 20330 1570 20350 2840
rect 18350 1540 20350 1570
rect 18350 1520 18390 1540
rect 18280 1500 18390 1520
rect 20310 1510 20350 1540
rect 20390 1510 20410 2890
rect 20310 1500 20410 1510
rect 18280 1480 20410 1500
rect 21980 2900 24110 2930
rect 21980 1520 22010 2900
rect 22050 2860 22090 2900
rect 24010 2890 24110 2900
rect 24010 2860 24050 2890
rect 22050 2840 24050 2860
rect 22050 1570 22070 2840
rect 24030 1570 24050 2840
rect 22050 1540 24050 1570
rect 22050 1520 22090 1540
rect 21980 1500 22090 1520
rect 24010 1510 24050 1540
rect 24090 1510 24110 2890
rect 24010 1500 24110 1510
rect 21980 1480 24110 1500
rect 25780 2900 27910 2930
rect 25780 1520 25810 2900
rect 25850 2860 25890 2900
rect 27810 2890 27910 2900
rect 27810 2860 27850 2890
rect 25850 2840 27850 2860
rect 25850 1570 25870 2840
rect 27830 1570 27850 2840
rect 25850 1540 27850 1570
rect 25850 1520 25890 1540
rect 25780 1500 25890 1520
rect 27810 1510 27850 1540
rect 27890 1510 27910 2890
rect 27810 1500 27910 1510
rect 25780 1480 27910 1500
<< nsubdiff >>
rect 7277 27079 7311 27103
rect 7277 26986 7311 27045
rect 7277 26928 7311 26952
rect 9853 27079 9887 27103
rect 9853 26986 9887 27045
rect 9853 26928 9887 26952
rect 12429 27079 12463 27103
rect 12429 26986 12463 27045
rect 12429 26928 12463 26952
rect 15005 27079 15039 27103
rect 15005 26986 15039 27045
rect 15005 26928 15039 26952
rect 17581 27079 17615 27103
rect 17581 26986 17615 27045
rect 17581 26928 17615 26952
rect 7277 26776 7311 26800
rect 7277 26683 7311 26742
rect 7277 26625 7311 26649
rect 12429 26776 12463 26800
rect 12429 26683 12463 26742
rect 12429 26625 12463 26649
rect 17581 26776 17615 26800
rect 17581 26683 17615 26742
rect 17581 26625 17615 26649
rect 9853 25991 9887 26015
rect 9853 25898 9887 25957
rect 9853 25840 9887 25864
rect 15005 25991 15039 26015
rect 15005 25898 15039 25957
rect 15005 25840 15039 25864
rect 7277 25688 7311 25712
rect 7277 25595 7311 25654
rect 7277 25537 7311 25561
rect 12429 25688 12463 25712
rect 12429 25595 12463 25654
rect 12429 25537 12463 25561
rect 17581 25688 17615 25712
rect 17581 25595 17615 25654
rect 17581 25537 17615 25561
rect 9853 24903 9887 24927
rect 9853 24810 9887 24869
rect 9853 24752 9887 24776
rect 15005 24903 15039 24927
rect 15005 24810 15039 24869
rect 15005 24752 15039 24776
rect 7277 24600 7311 24624
rect 7277 24507 7311 24566
rect 7277 24449 7311 24473
rect 12429 24600 12463 24624
rect 12429 24507 12463 24566
rect 12429 24449 12463 24473
rect 17581 24600 17615 24624
rect 17581 24507 17615 24566
rect 17581 24449 17615 24473
rect 9853 23815 9887 23839
rect 9853 23722 9887 23781
rect 9853 23664 9887 23688
rect 15005 23815 15039 23839
rect 15005 23722 15039 23781
rect 15005 23664 15039 23688
rect 7277 23512 7311 23536
rect 7277 23419 7311 23478
rect 7277 23361 7311 23385
rect 12429 23512 12463 23536
rect 12429 23419 12463 23478
rect 12429 23361 12463 23385
rect 17581 23512 17615 23536
rect 17581 23419 17615 23478
rect 17581 23361 17615 23385
rect 9853 22727 9887 22751
rect 9853 22634 9887 22693
rect 9853 22576 9887 22600
rect 15005 22727 15039 22751
rect 15005 22634 15039 22693
rect 15005 22576 15039 22600
rect 7277 22424 7311 22448
rect 7277 22331 7311 22390
rect 7277 22273 7311 22297
rect 12429 22424 12463 22448
rect 12429 22331 12463 22390
rect 12429 22273 12463 22297
rect 17581 22424 17615 22448
rect 17581 22331 17615 22390
rect 17581 22273 17615 22297
rect 9853 21639 9887 21663
rect 9853 21546 9887 21605
rect 9853 21488 9887 21512
rect 15005 21639 15039 21663
rect 15005 21546 15039 21605
rect 15005 21488 15039 21512
rect 7277 21336 7311 21360
rect 7277 21243 7311 21302
rect 7277 21185 7311 21209
rect 12429 21336 12463 21360
rect 12429 21243 12463 21302
rect 12429 21185 12463 21209
rect 17581 21336 17615 21360
rect 17581 21243 17615 21302
rect 17581 21185 17615 21209
rect 9853 20551 9887 20575
rect 9853 20458 9887 20517
rect 9853 20400 9887 20424
rect 15005 20551 15039 20575
rect 15005 20458 15039 20517
rect 15005 20400 15039 20424
rect 7277 20248 7311 20272
rect 7277 20155 7311 20214
rect 7277 20097 7311 20121
rect 12429 20248 12463 20272
rect 12429 20155 12463 20214
rect 12429 20097 12463 20121
rect 17581 20248 17615 20272
rect 17581 20155 17615 20214
rect 17581 20097 17615 20121
rect 9853 19463 9887 19487
rect 9853 19370 9887 19429
rect 9853 19312 9887 19336
rect 15005 19463 15039 19487
rect 15005 19370 15039 19429
rect 15005 19312 15039 19336
rect 7277 19160 7311 19184
rect 7277 19067 7311 19126
rect 7277 19009 7311 19033
rect 12429 19160 12463 19184
rect 12429 19067 12463 19126
rect 12429 19009 12463 19033
rect 17581 19160 17615 19184
rect 17581 19067 17615 19126
rect 17581 19009 17615 19033
rect 9853 18375 9887 18399
rect 9853 18282 9887 18341
rect 9853 18224 9887 18248
rect 15005 18375 15039 18399
rect 15005 18282 15039 18341
rect 15005 18224 15039 18248
rect 7277 18072 7311 18096
rect 7277 17979 7311 18038
rect 7277 17921 7311 17945
rect 12429 18072 12463 18096
rect 12429 17979 12463 18038
rect 12429 17921 12463 17945
rect 17581 18072 17615 18096
rect 17581 17979 17615 18038
rect 17581 17921 17615 17945
rect 9853 17287 9887 17311
rect 9853 17194 9887 17253
rect 9853 17136 9887 17160
rect 15005 17287 15039 17311
rect 15005 17194 15039 17253
rect 15005 17136 15039 17160
rect 7277 16984 7311 17008
rect 7277 16891 7311 16950
rect 7277 16833 7311 16857
rect 12429 16984 12463 17008
rect 12429 16891 12463 16950
rect 12429 16833 12463 16857
rect 17581 16984 17615 17008
rect 17581 16891 17615 16950
rect 17581 16833 17615 16857
rect 9853 16199 9887 16223
rect 9853 16106 9887 16165
rect 9853 16048 9887 16072
rect 15005 16199 15039 16223
rect 15005 16106 15039 16165
rect 15005 16048 15039 16072
rect 7277 15896 7311 15920
rect 7277 15803 7311 15862
rect 7277 15745 7311 15769
rect 12429 15896 12463 15920
rect 12429 15803 12463 15862
rect 12429 15745 12463 15769
rect 17581 15896 17615 15920
rect 17581 15803 17615 15862
rect 17581 15745 17615 15769
rect 9853 15111 9887 15135
rect 9853 15018 9887 15077
rect 9853 14960 9887 14984
rect 15005 15111 15039 15135
rect 15005 15018 15039 15077
rect 15005 14960 15039 14984
rect 7277 14808 7311 14832
rect 7277 14715 7311 14774
rect 7277 14657 7311 14681
rect 12429 14808 12463 14832
rect 12429 14715 12463 14774
rect 12429 14657 12463 14681
rect 17581 14808 17615 14832
rect 17581 14715 17615 14774
rect 17581 14657 17615 14681
rect 9853 14023 9887 14047
rect 9853 13930 9887 13989
rect 9853 13872 9887 13896
rect 15005 14023 15039 14047
rect 15005 13930 15039 13989
rect 15005 13872 15039 13896
rect 7277 13720 7311 13744
rect 7277 13627 7311 13686
rect 7277 13569 7311 13593
rect 12429 13720 12463 13744
rect 12429 13627 12463 13686
rect 12429 13569 12463 13593
rect 17581 13720 17615 13744
rect 17581 13627 17615 13686
rect 17581 13569 17615 13593
rect 9853 12935 9887 12959
rect 9853 12842 9887 12901
rect 9853 12784 9887 12808
rect 15005 12935 15039 12959
rect 15005 12842 15039 12901
rect 15005 12784 15039 12808
rect 7277 12632 7311 12656
rect 7277 12539 7311 12598
rect 7277 12481 7311 12505
rect 9853 12632 9887 12656
rect 9853 12539 9887 12598
rect 9853 12481 9887 12505
rect 12429 12632 12463 12656
rect 12429 12539 12463 12598
rect 12429 12481 12463 12505
rect 15005 12632 15039 12656
rect 15005 12539 15039 12598
rect 15005 12481 15039 12505
rect 17581 12632 17615 12656
rect 17581 12539 17615 12598
rect 17581 12481 17615 12505
rect 29580 7050 34840 7070
rect 29580 7010 29680 7050
rect 34760 7010 34840 7050
rect 29580 6990 34840 7010
rect 29580 4970 29600 6990
rect 29640 4990 29660 6990
rect 34760 6970 34840 6990
rect 34760 5030 34780 6970
rect 34820 5030 34840 6970
rect 34760 4990 34840 5030
rect 29640 4970 34840 4990
rect 29580 4930 29680 4970
rect 34780 4930 34840 4970
rect 29580 4910 34840 4930
rect 1290 4460 3410 4480
rect 1290 4440 1390 4460
rect 1290 3040 1310 4440
rect 1350 4420 1390 4440
rect 3310 4440 3410 4460
rect 3310 4420 3350 4440
rect 1350 4400 3350 4420
rect 1350 3100 1370 4400
rect 1350 3080 1390 3100
rect 3330 3080 3350 4400
rect 1350 3060 3350 3080
rect 1350 3040 1390 3060
rect 1290 3020 1390 3040
rect 3310 3040 3350 3060
rect 3390 3040 3410 4440
rect 3310 3020 3410 3040
rect 1290 3000 3410 3020
rect 4590 4460 6710 4480
rect 4590 4440 4690 4460
rect 4590 3040 4610 4440
rect 4650 4420 4690 4440
rect 6610 4440 6710 4460
rect 6610 4420 6650 4440
rect 4650 4400 6650 4420
rect 4650 3100 4670 4400
rect 4650 3080 4690 3100
rect 6630 3080 6650 4400
rect 4650 3060 6650 3080
rect 4650 3040 4690 3060
rect 4590 3020 4690 3040
rect 6610 3040 6650 3060
rect 6690 3040 6710 4440
rect 6610 3020 6710 3040
rect 4590 3000 6710 3020
rect 7890 4460 10010 4480
rect 7890 4440 7990 4460
rect 7890 3040 7910 4440
rect 7950 4420 7990 4440
rect 9910 4440 10010 4460
rect 9910 4420 9950 4440
rect 7950 4400 9950 4420
rect 7950 3100 7970 4400
rect 7950 3080 7990 3100
rect 9930 3080 9950 4400
rect 7950 3060 9950 3080
rect 7950 3040 7990 3060
rect 7890 3020 7990 3040
rect 9910 3040 9950 3060
rect 9990 3040 10010 4440
rect 9910 3020 10010 3040
rect 7890 3000 10010 3020
rect 11190 4460 13310 4480
rect 11190 4440 11290 4460
rect 11190 3040 11210 4440
rect 11250 4420 11290 4440
rect 13210 4440 13310 4460
rect 13210 4420 13250 4440
rect 11250 4400 13250 4420
rect 11250 3100 11270 4400
rect 11250 3080 11290 3100
rect 13230 3080 13250 4400
rect 11250 3060 13250 3080
rect 11250 3040 11290 3060
rect 11190 3020 11290 3040
rect 13210 3040 13250 3060
rect 13290 3040 13310 4440
rect 13210 3020 13310 3040
rect 11190 3000 13310 3020
rect 14790 4460 16910 4480
rect 14790 4440 14890 4460
rect 14790 3040 14810 4440
rect 14850 4420 14890 4440
rect 16810 4440 16910 4460
rect 16810 4420 16850 4440
rect 14850 4400 16850 4420
rect 14850 3100 14870 4400
rect 14850 3080 14890 3100
rect 16830 3080 16850 4400
rect 14850 3060 16850 3080
rect 14850 3040 14890 3060
rect 14790 3020 14890 3040
rect 16810 3040 16850 3060
rect 16890 3040 16910 4440
rect 16810 3020 16910 3040
rect 14790 3000 16910 3020
rect 18290 4460 20410 4480
rect 18290 4440 18390 4460
rect 18290 3040 18310 4440
rect 18350 4420 18390 4440
rect 20310 4440 20410 4460
rect 20310 4420 20350 4440
rect 18350 4400 20350 4420
rect 18350 3100 18370 4400
rect 18350 3080 18390 3100
rect 20330 3080 20350 4400
rect 18350 3060 20350 3080
rect 18350 3040 18390 3060
rect 18290 3020 18390 3040
rect 20310 3040 20350 3060
rect 20390 3040 20410 4440
rect 20310 3020 20410 3040
rect 18290 3000 20410 3020
rect 21990 4460 24110 4480
rect 21990 4440 22090 4460
rect 21990 3040 22010 4440
rect 22050 4420 22090 4440
rect 24010 4440 24110 4460
rect 24010 4420 24050 4440
rect 22050 4400 24050 4420
rect 22050 3100 22070 4400
rect 22050 3080 22090 3100
rect 24030 3080 24050 4400
rect 22050 3060 24050 3080
rect 22050 3040 22090 3060
rect 21990 3020 22090 3040
rect 24010 3040 24050 3060
rect 24090 3040 24110 4440
rect 24010 3020 24110 3040
rect 21990 3000 24110 3020
rect 25790 4460 27910 4480
rect 25790 4440 25890 4460
rect 25790 3040 25810 4440
rect 25850 4420 25890 4440
rect 27810 4440 27910 4460
rect 27810 4420 27850 4440
rect 25850 4400 27850 4420
rect 25850 3100 25870 4400
rect 25850 3080 25890 3100
rect 27830 3080 27850 4400
rect 25850 3060 27850 3080
rect 25850 3040 25890 3060
rect 25790 3020 25890 3040
rect 27810 3040 27850 3060
rect 27890 3040 27910 4440
rect 27810 3020 27910 3040
rect 25790 3000 27910 3020
<< psubdiffcont >>
rect 7277 27263 7311 27297
rect 9853 27263 9887 27297
rect 12429 27263 12463 27297
rect 15005 27263 15039 27297
rect 17581 27263 17615 27297
rect 7277 26431 7311 26465
rect 12429 26431 12463 26465
rect 17581 26431 17615 26465
rect 9853 26175 9887 26209
rect 15005 26175 15039 26209
rect 7277 25343 7311 25377
rect 12429 25343 12463 25377
rect 17581 25343 17615 25377
rect 9853 25087 9887 25121
rect 15005 25087 15039 25121
rect 7277 24255 7311 24289
rect 12429 24255 12463 24289
rect 17581 24255 17615 24289
rect 9853 23999 9887 24033
rect 15005 23999 15039 24033
rect 7277 23167 7311 23201
rect 12429 23167 12463 23201
rect 17581 23167 17615 23201
rect 9853 22911 9887 22945
rect 15005 22911 15039 22945
rect 7277 22079 7311 22113
rect 12429 22079 12463 22113
rect 17581 22079 17615 22113
rect 9853 21823 9887 21857
rect 15005 21823 15039 21857
rect 7277 20991 7311 21025
rect 12429 20991 12463 21025
rect 17581 20991 17615 21025
rect 9853 20735 9887 20769
rect 15005 20735 15039 20769
rect 7277 19903 7311 19937
rect 12429 19903 12463 19937
rect 17581 19903 17615 19937
rect 9853 19647 9887 19681
rect 15005 19647 15039 19681
rect 7277 18815 7311 18849
rect 12429 18815 12463 18849
rect 17581 18815 17615 18849
rect 9853 18559 9887 18593
rect 15005 18559 15039 18593
rect 7277 17727 7311 17761
rect 12429 17727 12463 17761
rect 17581 17727 17615 17761
rect 9853 17471 9887 17505
rect 15005 17471 15039 17505
rect 7277 16639 7311 16673
rect 12429 16639 12463 16673
rect 17581 16639 17615 16673
rect 9853 16383 9887 16417
rect 15005 16383 15039 16417
rect 7277 15551 7311 15585
rect 12429 15551 12463 15585
rect 17581 15551 17615 15585
rect 9853 15295 9887 15329
rect 15005 15295 15039 15329
rect 7277 14463 7311 14497
rect 12429 14463 12463 14497
rect 17581 14463 17615 14497
rect 9853 14207 9887 14241
rect 15005 14207 15039 14241
rect 7277 13375 7311 13409
rect 12429 13375 12463 13409
rect 17581 13375 17615 13409
rect 9853 13119 9887 13153
rect 15005 13119 15039 13153
rect 7277 12287 7311 12321
rect 9853 12287 9887 12321
rect 12429 12287 12463 12321
rect 15005 12287 15039 12321
rect 17581 12287 17615 12321
rect 25812 9190 28176 9224
rect 25716 7112 25750 9128
rect 28238 7112 28272 9128
rect 25812 7016 28176 7050
rect 16982 6850 17120 6884
rect 13382 6290 13520 6324
rect 10082 6010 10220 6044
rect 3482 5966 3620 6000
rect 3386 4772 3420 5904
rect 3682 4772 3716 5904
rect 3482 4676 3620 4710
rect 6782 5870 6920 5904
rect 6686 4772 6720 5808
rect 6982 4772 7016 5808
rect 6782 4676 6920 4710
rect 9986 4772 10020 5948
rect 10282 4772 10316 5948
rect 10082 4676 10220 4710
rect 13286 4772 13320 6228
rect 13582 4772 13616 6228
rect 13382 4676 13520 4710
rect 16886 4772 16920 6788
rect 17182 4772 17216 6788
rect 16982 4676 17120 4710
rect 20182 6850 20638 6884
rect 20086 4772 20120 6788
rect 20700 4772 20734 6788
rect 20182 4676 20638 4710
rect 23282 6850 24374 6884
rect 23186 4772 23220 6788
rect 24436 4772 24470 6788
rect 23282 4676 24374 4710
rect 25782 6850 28146 6884
rect 25686 4772 25720 6788
rect 28208 4772 28242 6788
rect 25782 4676 28146 4710
rect 29660 4770 34700 4810
rect 29580 4110 29620 4750
rect 34740 4130 34780 4790
rect 29660 4050 34720 4090
rect 440 2510 620 2690
rect 1310 1520 1350 2900
rect 1390 2860 3310 2900
rect 1390 1500 3310 1540
rect 3350 1510 3390 2890
rect 4610 1520 4650 2900
rect 4690 2860 6610 2900
rect 4690 1500 6610 1540
rect 6650 1510 6690 2890
rect 7910 1520 7950 2900
rect 7990 2860 9910 2900
rect 7990 1500 9910 1540
rect 9950 1510 9990 2890
rect 11210 1520 11250 2900
rect 11290 2860 13210 2900
rect 11290 1500 13210 1540
rect 13250 1510 13290 2890
rect 14810 1520 14850 2900
rect 14890 2860 16810 2900
rect 14890 1500 16810 1540
rect 16850 1510 16890 2890
rect 18310 1520 18350 2900
rect 18390 2860 20310 2900
rect 18390 1500 20310 1540
rect 20350 1510 20390 2890
rect 22010 1520 22050 2900
rect 22090 2860 24010 2900
rect 22090 1500 24010 1540
rect 24050 1510 24090 2890
rect 25810 1520 25850 2900
rect 25890 2860 27810 2900
rect 25890 1500 27810 1540
rect 27850 1510 27890 2890
<< nsubdiffcont >>
rect 7277 27045 7311 27079
rect 7277 26952 7311 26986
rect 9853 27045 9887 27079
rect 9853 26952 9887 26986
rect 12429 27045 12463 27079
rect 12429 26952 12463 26986
rect 15005 27045 15039 27079
rect 15005 26952 15039 26986
rect 17581 27045 17615 27079
rect 17581 26952 17615 26986
rect 7277 26742 7311 26776
rect 7277 26649 7311 26683
rect 12429 26742 12463 26776
rect 12429 26649 12463 26683
rect 17581 26742 17615 26776
rect 17581 26649 17615 26683
rect 9853 25957 9887 25991
rect 9853 25864 9887 25898
rect 15005 25957 15039 25991
rect 15005 25864 15039 25898
rect 7277 25654 7311 25688
rect 7277 25561 7311 25595
rect 12429 25654 12463 25688
rect 12429 25561 12463 25595
rect 17581 25654 17615 25688
rect 17581 25561 17615 25595
rect 9853 24869 9887 24903
rect 9853 24776 9887 24810
rect 15005 24869 15039 24903
rect 15005 24776 15039 24810
rect 7277 24566 7311 24600
rect 7277 24473 7311 24507
rect 12429 24566 12463 24600
rect 12429 24473 12463 24507
rect 17581 24566 17615 24600
rect 17581 24473 17615 24507
rect 9853 23781 9887 23815
rect 9853 23688 9887 23722
rect 15005 23781 15039 23815
rect 15005 23688 15039 23722
rect 7277 23478 7311 23512
rect 7277 23385 7311 23419
rect 12429 23478 12463 23512
rect 12429 23385 12463 23419
rect 17581 23478 17615 23512
rect 17581 23385 17615 23419
rect 9853 22693 9887 22727
rect 9853 22600 9887 22634
rect 15005 22693 15039 22727
rect 15005 22600 15039 22634
rect 7277 22390 7311 22424
rect 7277 22297 7311 22331
rect 12429 22390 12463 22424
rect 12429 22297 12463 22331
rect 17581 22390 17615 22424
rect 17581 22297 17615 22331
rect 9853 21605 9887 21639
rect 9853 21512 9887 21546
rect 15005 21605 15039 21639
rect 15005 21512 15039 21546
rect 7277 21302 7311 21336
rect 7277 21209 7311 21243
rect 12429 21302 12463 21336
rect 12429 21209 12463 21243
rect 17581 21302 17615 21336
rect 17581 21209 17615 21243
rect 9853 20517 9887 20551
rect 9853 20424 9887 20458
rect 15005 20517 15039 20551
rect 15005 20424 15039 20458
rect 7277 20214 7311 20248
rect 7277 20121 7311 20155
rect 12429 20214 12463 20248
rect 12429 20121 12463 20155
rect 17581 20214 17615 20248
rect 17581 20121 17615 20155
rect 9853 19429 9887 19463
rect 9853 19336 9887 19370
rect 15005 19429 15039 19463
rect 15005 19336 15039 19370
rect 7277 19126 7311 19160
rect 7277 19033 7311 19067
rect 12429 19126 12463 19160
rect 12429 19033 12463 19067
rect 17581 19126 17615 19160
rect 17581 19033 17615 19067
rect 9853 18341 9887 18375
rect 9853 18248 9887 18282
rect 15005 18341 15039 18375
rect 15005 18248 15039 18282
rect 7277 18038 7311 18072
rect 7277 17945 7311 17979
rect 12429 18038 12463 18072
rect 12429 17945 12463 17979
rect 17581 18038 17615 18072
rect 17581 17945 17615 17979
rect 9853 17253 9887 17287
rect 9853 17160 9887 17194
rect 15005 17253 15039 17287
rect 15005 17160 15039 17194
rect 7277 16950 7311 16984
rect 7277 16857 7311 16891
rect 12429 16950 12463 16984
rect 12429 16857 12463 16891
rect 17581 16950 17615 16984
rect 17581 16857 17615 16891
rect 9853 16165 9887 16199
rect 9853 16072 9887 16106
rect 15005 16165 15039 16199
rect 15005 16072 15039 16106
rect 7277 15862 7311 15896
rect 7277 15769 7311 15803
rect 12429 15862 12463 15896
rect 12429 15769 12463 15803
rect 17581 15862 17615 15896
rect 17581 15769 17615 15803
rect 9853 15077 9887 15111
rect 9853 14984 9887 15018
rect 15005 15077 15039 15111
rect 15005 14984 15039 15018
rect 7277 14774 7311 14808
rect 7277 14681 7311 14715
rect 12429 14774 12463 14808
rect 12429 14681 12463 14715
rect 17581 14774 17615 14808
rect 17581 14681 17615 14715
rect 9853 13989 9887 14023
rect 9853 13896 9887 13930
rect 15005 13989 15039 14023
rect 15005 13896 15039 13930
rect 7277 13686 7311 13720
rect 7277 13593 7311 13627
rect 12429 13686 12463 13720
rect 12429 13593 12463 13627
rect 17581 13686 17615 13720
rect 17581 13593 17615 13627
rect 9853 12901 9887 12935
rect 9853 12808 9887 12842
rect 15005 12901 15039 12935
rect 15005 12808 15039 12842
rect 7277 12598 7311 12632
rect 7277 12505 7311 12539
rect 9853 12598 9887 12632
rect 9853 12505 9887 12539
rect 12429 12598 12463 12632
rect 12429 12505 12463 12539
rect 15005 12598 15039 12632
rect 15005 12505 15039 12539
rect 17581 12598 17615 12632
rect 17581 12505 17615 12539
rect 29680 7010 34760 7050
rect 29600 4970 29640 6990
rect 34780 5030 34820 6970
rect 29680 4930 34780 4970
rect 1310 3040 1350 4440
rect 1390 4420 3310 4460
rect 1390 3020 3310 3060
rect 3350 3040 3390 4440
rect 4610 3040 4650 4440
rect 4690 4420 6610 4460
rect 4690 3020 6610 3060
rect 6650 3040 6690 4440
rect 7910 3040 7950 4440
rect 7990 4420 9910 4460
rect 7990 3020 9910 3060
rect 9950 3040 9990 4440
rect 11210 3040 11250 4440
rect 11290 4420 13210 4460
rect 11290 3020 13210 3060
rect 13250 3040 13290 4440
rect 14810 3040 14850 4440
rect 14890 4420 16810 4460
rect 14890 3020 16810 3060
rect 16850 3040 16890 4440
rect 18310 3040 18350 4440
rect 18390 4420 20310 4460
rect 18390 3020 20310 3060
rect 20350 3040 20390 4440
rect 22010 3040 22050 4440
rect 22090 4420 24010 4460
rect 22090 3020 24010 3060
rect 24050 3040 24090 4440
rect 25810 3040 25850 4440
rect 25890 4420 27810 4460
rect 25890 3020 27810 3060
rect 27850 3040 27890 4440
<< poly >>
rect 5027 27361 5145 27387
rect 5303 27361 5421 27387
rect 5587 27361 5617 27387
rect 5673 27361 5703 27387
rect 5759 27361 5789 27387
rect 5845 27361 5875 27387
rect 5942 27361 5972 27387
rect 6223 27361 7169 27387
rect 7419 27361 7537 27387
rect 7695 27361 8641 27387
rect 8799 27361 9745 27387
rect 10179 27361 10209 27387
rect 10267 27361 10297 27387
rect 10639 27361 11217 27387
rect 11375 27361 12321 27387
rect 12571 27361 12689 27387
rect 12847 27361 13793 27387
rect 13951 27361 14897 27387
rect 15147 27361 15265 27387
rect 15423 27361 16369 27387
rect 16527 27361 17473 27387
rect 17815 27361 18393 27387
rect 18559 27361 18589 27387
rect 18645 27361 18675 27387
rect 18731 27361 18761 27387
rect 18817 27361 18847 27387
rect 18914 27361 18944 27387
rect 19287 27361 19865 27387
rect 20023 27361 20141 27387
rect 5027 27225 5145 27251
rect 5107 27223 5145 27225
rect 5303 27225 5421 27251
rect 5303 27223 5341 27225
rect 5107 27207 5173 27223
rect 4999 27167 5065 27183
rect 4999 27133 5015 27167
rect 5049 27133 5065 27167
rect 5107 27173 5123 27207
rect 5157 27173 5173 27207
rect 5107 27157 5173 27173
rect 5275 27207 5341 27223
rect 5275 27173 5291 27207
rect 5325 27173 5341 27207
rect 5587 27204 5617 27277
rect 5673 27204 5703 27277
rect 5759 27204 5789 27277
rect 5845 27204 5875 27277
rect 5942 27209 5972 27277
rect 6223 27225 7169 27251
rect 7419 27225 7537 27251
rect 7695 27225 8641 27251
rect 8799 27225 9745 27251
rect 10179 27242 10209 27257
rect 5587 27198 5875 27204
rect 5587 27193 5876 27198
rect 5275 27157 5341 27173
rect 5383 27167 5449 27183
rect 5587 27171 5651 27193
rect 4999 27117 5065 27133
rect 5027 27115 5065 27117
rect 5383 27133 5399 27167
rect 5433 27133 5449 27167
rect 5383 27117 5449 27133
rect 5588 27159 5651 27171
rect 5685 27159 5719 27193
rect 5753 27159 5787 27193
rect 5821 27159 5876 27193
rect 5588 27149 5876 27159
rect 5383 27115 5421 27117
rect 5027 27085 5145 27115
rect 5303 27085 5421 27115
rect 5588 27111 5618 27149
rect 5674 27111 5704 27149
rect 5760 27111 5790 27149
rect 5846 27111 5876 27149
rect 5923 27193 5983 27209
rect 5923 27159 5933 27193
rect 5967 27159 5983 27193
rect 5923 27143 5983 27159
rect 6223 27203 6677 27225
rect 7419 27223 7457 27225
rect 6223 27169 6499 27203
rect 6533 27169 6677 27203
rect 7391 27207 7457 27223
rect 6223 27153 6677 27169
rect 6719 27167 7169 27183
rect 5942 27111 5972 27143
rect 6719 27133 6863 27167
rect 6897 27133 7169 27167
rect 7391 27173 7407 27207
rect 7441 27173 7457 27207
rect 7695 27203 8149 27225
rect 7391 27157 7457 27173
rect 7499 27167 7565 27183
rect 6719 27111 7169 27133
rect 7499 27133 7515 27167
rect 7549 27133 7565 27167
rect 7695 27169 7971 27203
rect 8005 27169 8149 27203
rect 8799 27203 9253 27225
rect 10173 27218 10209 27242
rect 10173 27209 10203 27218
rect 7695 27153 8149 27169
rect 8191 27167 8641 27183
rect 7499 27117 7565 27133
rect 8191 27133 8335 27167
rect 8369 27133 8641 27167
rect 8799 27169 9075 27203
rect 9109 27169 9253 27203
rect 10127 27193 10203 27209
rect 10267 27196 10297 27257
rect 10639 27225 11217 27251
rect 11375 27225 12321 27251
rect 12571 27225 12689 27251
rect 12847 27225 13793 27251
rect 13951 27225 14897 27251
rect 15147 27225 15265 27251
rect 15423 27225 16369 27251
rect 16527 27225 17473 27251
rect 17815 27225 18393 27251
rect 10639 27203 10911 27225
rect 8799 27153 9253 27169
rect 9295 27167 9745 27183
rect 7499 27115 7537 27117
rect 6223 27085 7169 27111
rect 7419 27085 7537 27115
rect 8191 27111 8641 27133
rect 9295 27133 9439 27167
rect 9473 27133 9745 27167
rect 10127 27159 10137 27193
rect 10171 27159 10203 27193
rect 10127 27143 10203 27159
rect 9295 27111 9745 27133
rect 7695 27085 8641 27111
rect 8799 27085 9745 27111
rect 10173 27108 10203 27143
rect 10245 27180 10299 27196
rect 10245 27146 10255 27180
rect 10289 27146 10299 27180
rect 10639 27169 10655 27203
rect 10689 27169 10758 27203
rect 10792 27169 10861 27203
rect 10895 27169 10911 27203
rect 11375 27203 11829 27225
rect 12571 27223 12609 27225
rect 10639 27153 10911 27169
rect 10953 27167 11217 27183
rect 10245 27130 10299 27146
rect 10953 27133 10969 27167
rect 11003 27133 11068 27167
rect 11102 27133 11167 27167
rect 11201 27133 11217 27167
rect 11375 27169 11651 27203
rect 11685 27169 11829 27203
rect 12543 27207 12609 27223
rect 11375 27153 11829 27169
rect 11871 27167 12321 27183
rect 10173 27084 10209 27108
rect 10179 27069 10209 27084
rect 10267 27069 10297 27130
rect 10953 27111 11217 27133
rect 11871 27133 12015 27167
rect 12049 27133 12321 27167
rect 12543 27173 12559 27207
rect 12593 27173 12609 27207
rect 12847 27203 13301 27225
rect 12543 27157 12609 27173
rect 12651 27167 12717 27183
rect 11871 27111 12321 27133
rect 12651 27133 12667 27167
rect 12701 27133 12717 27167
rect 12847 27169 13123 27203
rect 13157 27169 13301 27203
rect 13951 27203 14405 27225
rect 15147 27223 15185 27225
rect 12847 27153 13301 27169
rect 13343 27167 13793 27183
rect 12651 27117 12717 27133
rect 13343 27133 13487 27167
rect 13521 27133 13793 27167
rect 13951 27169 14227 27203
rect 14261 27169 14405 27203
rect 15119 27207 15185 27223
rect 13951 27153 14405 27169
rect 14447 27167 14897 27183
rect 12651 27115 12689 27117
rect 10639 27085 11217 27111
rect 11375 27085 12321 27111
rect 12571 27085 12689 27115
rect 13343 27111 13793 27133
rect 14447 27133 14591 27167
rect 14625 27133 14897 27167
rect 15119 27173 15135 27207
rect 15169 27173 15185 27207
rect 15423 27203 15877 27225
rect 15119 27157 15185 27173
rect 15227 27167 15293 27183
rect 14447 27111 14897 27133
rect 15227 27133 15243 27167
rect 15277 27133 15293 27167
rect 15423 27169 15699 27203
rect 15733 27169 15877 27203
rect 16527 27203 16981 27225
rect 15423 27153 15877 27169
rect 15919 27167 16369 27183
rect 15227 27117 15293 27133
rect 15919 27133 16063 27167
rect 16097 27133 16369 27167
rect 16527 27169 16803 27203
rect 16837 27169 16981 27203
rect 17815 27203 18087 27225
rect 16527 27153 16981 27169
rect 17023 27167 17473 27183
rect 15227 27115 15265 27117
rect 12847 27085 13793 27111
rect 13951 27085 14897 27111
rect 15147 27085 15265 27115
rect 15919 27111 16369 27133
rect 17023 27133 17167 27167
rect 17201 27133 17473 27167
rect 17815 27169 17831 27203
rect 17865 27169 17934 27203
rect 17968 27169 18037 27203
rect 18071 27169 18087 27203
rect 18559 27204 18589 27277
rect 18645 27204 18675 27277
rect 18731 27204 18761 27277
rect 18817 27204 18847 27277
rect 18914 27209 18944 27277
rect 19287 27225 19865 27251
rect 20023 27225 20141 27251
rect 18559 27198 18847 27204
rect 18559 27193 18848 27198
rect 17815 27153 18087 27169
rect 18129 27167 18393 27183
rect 18559 27171 18623 27193
rect 17023 27111 17473 27133
rect 18129 27133 18145 27167
rect 18179 27133 18244 27167
rect 18278 27133 18343 27167
rect 18377 27133 18393 27167
rect 18129 27111 18393 27133
rect 18560 27159 18623 27171
rect 18657 27159 18691 27193
rect 18725 27159 18759 27193
rect 18793 27159 18848 27193
rect 18560 27149 18848 27159
rect 18560 27111 18590 27149
rect 18646 27111 18676 27149
rect 18732 27111 18762 27149
rect 18818 27111 18848 27149
rect 18895 27193 18955 27209
rect 18895 27159 18905 27193
rect 18939 27159 18955 27193
rect 18895 27143 18955 27159
rect 19287 27203 19559 27225
rect 20023 27223 20061 27225
rect 19287 27169 19303 27203
rect 19337 27169 19406 27203
rect 19440 27169 19509 27203
rect 19543 27169 19559 27203
rect 19995 27207 20061 27223
rect 19287 27153 19559 27169
rect 19601 27167 19865 27183
rect 18914 27111 18944 27143
rect 19601 27133 19617 27167
rect 19651 27133 19716 27167
rect 19750 27133 19815 27167
rect 19849 27133 19865 27167
rect 19995 27173 20011 27207
rect 20045 27173 20061 27207
rect 19995 27157 20061 27173
rect 20103 27167 20169 27183
rect 19601 27111 19865 27133
rect 20103 27133 20119 27167
rect 20153 27133 20169 27167
rect 20103 27117 20169 27133
rect 20103 27115 20141 27117
rect 15423 27085 16369 27111
rect 16527 27085 17473 27111
rect 17815 27085 18393 27111
rect 19287 27085 19865 27111
rect 20023 27085 20141 27115
rect 5027 26885 5145 26911
rect 5303 26885 5421 26911
rect 5588 26885 5618 26911
rect 5674 26885 5704 26911
rect 5760 26885 5790 26911
rect 5846 26885 5876 26911
rect 5942 26885 5972 26911
rect 6223 26885 7169 26911
rect 7419 26885 7537 26911
rect 7695 26885 8641 26911
rect 8799 26885 9745 26911
rect 10179 26885 10209 26911
rect 10267 26885 10297 26911
rect 10639 26885 11217 26911
rect 11375 26885 12321 26911
rect 12571 26885 12689 26911
rect 12847 26885 13793 26911
rect 13951 26885 14897 26911
rect 15147 26885 15265 26911
rect 15423 26885 16369 26911
rect 16527 26885 17473 26911
rect 17815 26885 18393 26911
rect 18560 26885 18590 26911
rect 18646 26885 18676 26911
rect 18732 26885 18762 26911
rect 18818 26885 18848 26911
rect 18914 26885 18944 26911
rect 19287 26885 19865 26911
rect 20023 26885 20141 26911
rect 5027 26817 5145 26843
rect 5487 26817 6065 26843
rect 6223 26817 7169 26843
rect 7511 26817 7905 26843
rect 8063 26817 9009 26843
rect 9167 26817 10113 26843
rect 10271 26817 11217 26843
rect 11375 26817 12321 26843
rect 12663 26817 13057 26843
rect 13215 26817 14161 26843
rect 14319 26817 15265 26843
rect 15423 26817 16369 26843
rect 16527 26817 17473 26843
rect 17815 26817 18761 26843
rect 18919 26817 19865 26843
rect 20023 26817 20141 26843
rect 5027 26613 5145 26643
rect 5487 26617 6065 26643
rect 6223 26617 7169 26643
rect 7511 26617 7905 26643
rect 8063 26617 9009 26643
rect 9167 26617 10113 26643
rect 10271 26617 11217 26643
rect 11375 26617 12321 26643
rect 12663 26617 13057 26643
rect 13215 26617 14161 26643
rect 14319 26617 15265 26643
rect 15423 26617 16369 26643
rect 16527 26617 17473 26643
rect 17815 26617 18761 26643
rect 18919 26617 19865 26643
rect 5027 26611 5065 26613
rect 4999 26595 5065 26611
rect 4999 26561 5015 26595
rect 5049 26561 5065 26595
rect 5801 26595 6065 26617
rect 4999 26545 5065 26561
rect 5107 26555 5173 26571
rect 5107 26521 5123 26555
rect 5157 26521 5173 26555
rect 5107 26505 5173 26521
rect 5487 26559 5759 26575
rect 5487 26525 5503 26559
rect 5537 26525 5606 26559
rect 5640 26525 5709 26559
rect 5743 26525 5759 26559
rect 5801 26561 5817 26595
rect 5851 26561 5916 26595
rect 5950 26561 6015 26595
rect 6049 26561 6065 26595
rect 6719 26595 7169 26617
rect 5801 26545 6065 26561
rect 6223 26559 6677 26575
rect 5107 26503 5145 26505
rect 5027 26477 5145 26503
rect 5487 26503 5759 26525
rect 6223 26525 6499 26559
rect 6533 26525 6677 26559
rect 6719 26561 6863 26595
rect 6897 26561 7169 26595
rect 7729 26595 7905 26617
rect 6719 26545 7169 26561
rect 7511 26559 7687 26575
rect 6223 26503 6677 26525
rect 7511 26525 7527 26559
rect 7561 26525 7637 26559
rect 7671 26525 7687 26559
rect 7729 26561 7745 26595
rect 7779 26561 7855 26595
rect 7889 26561 7905 26595
rect 8559 26595 9009 26617
rect 7729 26545 7905 26561
rect 8063 26559 8517 26575
rect 7511 26503 7687 26525
rect 8063 26525 8339 26559
rect 8373 26525 8517 26559
rect 8559 26561 8703 26595
rect 8737 26561 9009 26595
rect 9663 26595 10113 26617
rect 8559 26545 9009 26561
rect 9167 26559 9621 26575
rect 8063 26503 8517 26525
rect 9167 26525 9443 26559
rect 9477 26525 9621 26559
rect 9663 26561 9807 26595
rect 9841 26561 10113 26595
rect 10767 26595 11217 26617
rect 9663 26545 10113 26561
rect 10271 26559 10725 26575
rect 9167 26503 9621 26525
rect 10271 26525 10547 26559
rect 10581 26525 10725 26559
rect 10767 26561 10911 26595
rect 10945 26561 11217 26595
rect 11871 26595 12321 26617
rect 10767 26545 11217 26561
rect 11375 26559 11829 26575
rect 10271 26503 10725 26525
rect 11375 26525 11651 26559
rect 11685 26525 11829 26559
rect 11871 26561 12015 26595
rect 12049 26561 12321 26595
rect 12881 26595 13057 26617
rect 11871 26545 12321 26561
rect 12663 26559 12839 26575
rect 11375 26503 11829 26525
rect 12663 26525 12679 26559
rect 12713 26525 12789 26559
rect 12823 26525 12839 26559
rect 12881 26561 12897 26595
rect 12931 26561 13007 26595
rect 13041 26561 13057 26595
rect 13711 26595 14161 26617
rect 12881 26545 13057 26561
rect 13215 26559 13669 26575
rect 12663 26503 12839 26525
rect 13215 26525 13491 26559
rect 13525 26525 13669 26559
rect 13711 26561 13855 26595
rect 13889 26561 14161 26595
rect 14815 26595 15265 26617
rect 13711 26545 14161 26561
rect 14319 26559 14773 26575
rect 13215 26503 13669 26525
rect 14319 26525 14595 26559
rect 14629 26525 14773 26559
rect 14815 26561 14959 26595
rect 14993 26561 15265 26595
rect 15919 26595 16369 26617
rect 14815 26545 15265 26561
rect 15423 26559 15877 26575
rect 14319 26503 14773 26525
rect 15423 26525 15699 26559
rect 15733 26525 15877 26559
rect 15919 26561 16063 26595
rect 16097 26561 16369 26595
rect 17023 26595 17473 26617
rect 15919 26545 16369 26561
rect 16527 26559 16981 26575
rect 15423 26503 15877 26525
rect 16527 26525 16803 26559
rect 16837 26525 16981 26559
rect 17023 26561 17167 26595
rect 17201 26561 17473 26595
rect 18311 26595 18761 26617
rect 17023 26545 17473 26561
rect 17815 26559 18269 26575
rect 16527 26503 16981 26525
rect 17815 26525 18091 26559
rect 18125 26525 18269 26559
rect 18311 26561 18455 26595
rect 18489 26561 18761 26595
rect 19415 26595 19865 26617
rect 20023 26613 20141 26643
rect 18311 26545 18761 26561
rect 18919 26559 19373 26575
rect 17815 26503 18269 26525
rect 18919 26525 19195 26559
rect 19229 26525 19373 26559
rect 19415 26561 19559 26595
rect 19593 26561 19865 26595
rect 20103 26611 20141 26613
rect 20103 26595 20169 26611
rect 19415 26545 19865 26561
rect 19995 26555 20061 26571
rect 18919 26503 19373 26525
rect 19995 26521 20011 26555
rect 20045 26521 20061 26555
rect 20103 26561 20119 26595
rect 20153 26561 20169 26595
rect 20103 26545 20169 26561
rect 19995 26505 20061 26521
rect 20023 26503 20061 26505
rect 5487 26477 6065 26503
rect 6223 26477 7169 26503
rect 7511 26477 7905 26503
rect 8063 26477 9009 26503
rect 9167 26477 10113 26503
rect 10271 26477 11217 26503
rect 11375 26477 12321 26503
rect 12663 26477 13057 26503
rect 13215 26477 14161 26503
rect 14319 26477 15265 26503
rect 15423 26477 16369 26503
rect 16527 26477 17473 26503
rect 17815 26477 18761 26503
rect 18919 26477 19865 26503
rect 20023 26477 20141 26503
rect 5027 26341 5145 26367
rect 5487 26341 6065 26367
rect 6223 26341 7169 26367
rect 7511 26341 7905 26367
rect 8063 26341 9009 26367
rect 9167 26341 10113 26367
rect 10271 26341 11217 26367
rect 11375 26341 12321 26367
rect 12663 26341 13057 26367
rect 13215 26341 14161 26367
rect 14319 26341 15265 26367
rect 15423 26341 16369 26367
rect 16527 26341 17473 26367
rect 17815 26341 18761 26367
rect 18919 26341 19865 26367
rect 20023 26341 20141 26367
rect 5027 26273 5145 26299
rect 5487 26273 6433 26299
rect 6591 26273 7537 26299
rect 7695 26273 8641 26299
rect 8799 26273 9745 26299
rect 10087 26273 10481 26299
rect 10639 26273 11585 26299
rect 11743 26273 12689 26299
rect 12847 26273 13793 26299
rect 13951 26273 14897 26299
rect 15239 26273 15449 26299
rect 15607 26273 16553 26299
rect 16711 26273 17657 26299
rect 17815 26273 18761 26299
rect 18919 26273 19865 26299
rect 20023 26273 20141 26299
rect 5027 26137 5145 26163
rect 5107 26135 5145 26137
rect 5487 26137 6433 26163
rect 6591 26137 7537 26163
rect 7695 26137 8641 26163
rect 8799 26137 9745 26163
rect 10087 26137 10481 26163
rect 10639 26137 11585 26163
rect 11743 26137 12689 26163
rect 12847 26137 13793 26163
rect 13951 26137 14897 26163
rect 15239 26137 15449 26163
rect 15607 26137 16553 26163
rect 16711 26137 17657 26163
rect 17815 26137 18761 26163
rect 18919 26137 19865 26163
rect 20023 26137 20141 26163
rect 5107 26119 5173 26135
rect 4999 26079 5065 26095
rect 4999 26045 5015 26079
rect 5049 26045 5065 26079
rect 5107 26085 5123 26119
rect 5157 26085 5173 26119
rect 5107 26069 5173 26085
rect 5487 26115 5941 26137
rect 5487 26081 5763 26115
rect 5797 26081 5941 26115
rect 6591 26115 7045 26137
rect 5487 26065 5941 26081
rect 5983 26079 6433 26095
rect 4999 26029 5065 26045
rect 5027 26027 5065 26029
rect 5983 26045 6127 26079
rect 6161 26045 6433 26079
rect 6591 26081 6867 26115
rect 6901 26081 7045 26115
rect 7695 26115 8149 26137
rect 6591 26065 7045 26081
rect 7087 26079 7537 26095
rect 5027 25997 5145 26027
rect 5983 26023 6433 26045
rect 7087 26045 7231 26079
rect 7265 26045 7537 26079
rect 7695 26081 7971 26115
rect 8005 26081 8149 26115
rect 8799 26115 9253 26137
rect 7695 26065 8149 26081
rect 8191 26079 8641 26095
rect 7087 26023 7537 26045
rect 8191 26045 8335 26079
rect 8369 26045 8641 26079
rect 8799 26081 9075 26115
rect 9109 26081 9253 26115
rect 10087 26115 10263 26137
rect 8799 26065 9253 26081
rect 9295 26079 9745 26095
rect 8191 26023 8641 26045
rect 9295 26045 9439 26079
rect 9473 26045 9745 26079
rect 10087 26081 10103 26115
rect 10137 26081 10213 26115
rect 10247 26081 10263 26115
rect 10639 26115 11093 26137
rect 10087 26065 10263 26081
rect 10305 26079 10481 26095
rect 9295 26023 9745 26045
rect 10305 26045 10321 26079
rect 10355 26045 10431 26079
rect 10465 26045 10481 26079
rect 10639 26081 10915 26115
rect 10949 26081 11093 26115
rect 11743 26115 12197 26137
rect 10639 26065 11093 26081
rect 11135 26079 11585 26095
rect 10305 26023 10481 26045
rect 11135 26045 11279 26079
rect 11313 26045 11585 26079
rect 11743 26081 12019 26115
rect 12053 26081 12197 26115
rect 12847 26115 13301 26137
rect 11743 26065 12197 26081
rect 12239 26079 12689 26095
rect 11135 26023 11585 26045
rect 12239 26045 12383 26079
rect 12417 26045 12689 26079
rect 12847 26081 13123 26115
rect 13157 26081 13301 26115
rect 13951 26115 14405 26137
rect 15239 26131 15323 26137
rect 12847 26065 13301 26081
rect 13343 26079 13793 26095
rect 12239 26023 12689 26045
rect 13343 26045 13487 26079
rect 13521 26045 13793 26079
rect 13951 26081 14227 26115
rect 14261 26081 14405 26115
rect 15181 26115 15323 26131
rect 13951 26065 14405 26081
rect 14447 26079 14897 26095
rect 13343 26023 13793 26045
rect 14447 26045 14591 26079
rect 14625 26045 14897 26079
rect 15181 26081 15197 26115
rect 15231 26081 15323 26115
rect 15607 26115 16061 26137
rect 15181 26065 15323 26081
rect 15365 26079 15507 26095
rect 14447 26023 14897 26045
rect 15365 26045 15457 26079
rect 15491 26045 15507 26079
rect 15607 26081 15883 26115
rect 15917 26081 16061 26115
rect 16711 26115 17165 26137
rect 15607 26065 16061 26081
rect 16103 26079 16553 26095
rect 15365 26029 15507 26045
rect 16103 26045 16247 26079
rect 16281 26045 16553 26079
rect 16711 26081 16987 26115
rect 17021 26081 17165 26115
rect 17815 26115 18269 26137
rect 16711 26065 17165 26081
rect 17207 26079 17657 26095
rect 15365 26023 15449 26029
rect 16103 26023 16553 26045
rect 17207 26045 17351 26079
rect 17385 26045 17657 26079
rect 17815 26081 18091 26115
rect 18125 26081 18269 26115
rect 18919 26115 19373 26137
rect 20023 26135 20061 26137
rect 17815 26065 18269 26081
rect 18311 26079 18761 26095
rect 17207 26023 17657 26045
rect 18311 26045 18455 26079
rect 18489 26045 18761 26079
rect 18919 26081 19195 26115
rect 19229 26081 19373 26115
rect 19995 26119 20061 26135
rect 18919 26065 19373 26081
rect 19415 26079 19865 26095
rect 18311 26023 18761 26045
rect 19415 26045 19559 26079
rect 19593 26045 19865 26079
rect 19995 26085 20011 26119
rect 20045 26085 20061 26119
rect 19995 26069 20061 26085
rect 20103 26079 20169 26095
rect 19415 26023 19865 26045
rect 20103 26045 20119 26079
rect 20153 26045 20169 26079
rect 20103 26029 20169 26045
rect 20103 26027 20141 26029
rect 5487 25997 6433 26023
rect 6591 25997 7537 26023
rect 7695 25997 8641 26023
rect 8799 25997 9745 26023
rect 10087 25997 10481 26023
rect 10639 25997 11585 26023
rect 11743 25997 12689 26023
rect 12847 25997 13793 26023
rect 13951 25997 14897 26023
rect 15239 25997 15449 26023
rect 15607 25997 16553 26023
rect 16711 25997 17657 26023
rect 17815 25997 18761 26023
rect 18919 25997 19865 26023
rect 20023 25997 20141 26027
rect 5027 25797 5145 25823
rect 5487 25797 6433 25823
rect 6591 25797 7537 25823
rect 7695 25797 8641 25823
rect 8799 25797 9745 25823
rect 10087 25797 10481 25823
rect 10639 25797 11585 25823
rect 11743 25797 12689 25823
rect 12847 25797 13793 25823
rect 13951 25797 14897 25823
rect 15239 25797 15449 25823
rect 15607 25797 16553 25823
rect 16711 25797 17657 25823
rect 17815 25797 18761 25823
rect 18919 25797 19865 25823
rect 20023 25797 20141 25823
rect 5027 25729 5145 25755
rect 5487 25729 6065 25755
rect 6223 25729 7169 25755
rect 7511 25729 7905 25755
rect 8063 25729 9009 25755
rect 9167 25729 10113 25755
rect 10271 25729 11217 25755
rect 11375 25729 12321 25755
rect 12663 25729 13057 25755
rect 13215 25729 14161 25755
rect 14319 25729 15265 25755
rect 15423 25729 16369 25755
rect 16527 25729 17473 25755
rect 17815 25729 18761 25755
rect 18919 25729 19865 25755
rect 20023 25729 20141 25755
rect 5027 25525 5145 25555
rect 5487 25529 6065 25555
rect 6223 25529 7169 25555
rect 7511 25529 7905 25555
rect 8063 25529 9009 25555
rect 9167 25529 10113 25555
rect 10271 25529 11217 25555
rect 11375 25529 12321 25555
rect 12663 25529 13057 25555
rect 13215 25529 14161 25555
rect 14319 25529 15265 25555
rect 15423 25529 16369 25555
rect 16527 25529 17473 25555
rect 17815 25529 18761 25555
rect 18919 25529 19865 25555
rect 5027 25523 5065 25525
rect 4999 25507 5065 25523
rect 4999 25473 5015 25507
rect 5049 25473 5065 25507
rect 5801 25507 6065 25529
rect 4999 25457 5065 25473
rect 5107 25467 5173 25483
rect 5107 25433 5123 25467
rect 5157 25433 5173 25467
rect 5107 25417 5173 25433
rect 5487 25471 5759 25487
rect 5487 25437 5503 25471
rect 5537 25437 5606 25471
rect 5640 25437 5709 25471
rect 5743 25437 5759 25471
rect 5801 25473 5817 25507
rect 5851 25473 5916 25507
rect 5950 25473 6015 25507
rect 6049 25473 6065 25507
rect 6719 25507 7169 25529
rect 5801 25457 6065 25473
rect 6223 25471 6677 25487
rect 5107 25415 5145 25417
rect 5027 25389 5145 25415
rect 5487 25415 5759 25437
rect 6223 25437 6499 25471
rect 6533 25437 6677 25471
rect 6719 25473 6863 25507
rect 6897 25473 7169 25507
rect 7729 25507 7905 25529
rect 6719 25457 7169 25473
rect 7511 25471 7687 25487
rect 6223 25415 6677 25437
rect 7511 25437 7527 25471
rect 7561 25437 7637 25471
rect 7671 25437 7687 25471
rect 7729 25473 7745 25507
rect 7779 25473 7855 25507
rect 7889 25473 7905 25507
rect 8559 25507 9009 25529
rect 7729 25457 7905 25473
rect 8063 25471 8517 25487
rect 7511 25415 7687 25437
rect 8063 25437 8339 25471
rect 8373 25437 8517 25471
rect 8559 25473 8703 25507
rect 8737 25473 9009 25507
rect 9663 25507 10113 25529
rect 8559 25457 9009 25473
rect 9167 25471 9621 25487
rect 8063 25415 8517 25437
rect 9167 25437 9443 25471
rect 9477 25437 9621 25471
rect 9663 25473 9807 25507
rect 9841 25473 10113 25507
rect 10767 25507 11217 25529
rect 9663 25457 10113 25473
rect 10271 25471 10725 25487
rect 9167 25415 9621 25437
rect 10271 25437 10547 25471
rect 10581 25437 10725 25471
rect 10767 25473 10911 25507
rect 10945 25473 11217 25507
rect 11871 25507 12321 25529
rect 10767 25457 11217 25473
rect 11375 25471 11829 25487
rect 10271 25415 10725 25437
rect 11375 25437 11651 25471
rect 11685 25437 11829 25471
rect 11871 25473 12015 25507
rect 12049 25473 12321 25507
rect 12881 25507 13057 25529
rect 11871 25457 12321 25473
rect 12663 25471 12839 25487
rect 11375 25415 11829 25437
rect 12663 25437 12679 25471
rect 12713 25437 12789 25471
rect 12823 25437 12839 25471
rect 12881 25473 12897 25507
rect 12931 25473 13007 25507
rect 13041 25473 13057 25507
rect 13711 25507 14161 25529
rect 12881 25457 13057 25473
rect 13215 25471 13669 25487
rect 12663 25415 12839 25437
rect 13215 25437 13491 25471
rect 13525 25437 13669 25471
rect 13711 25473 13855 25507
rect 13889 25473 14161 25507
rect 14815 25507 15265 25529
rect 13711 25457 14161 25473
rect 14319 25471 14773 25487
rect 13215 25415 13669 25437
rect 14319 25437 14595 25471
rect 14629 25437 14773 25471
rect 14815 25473 14959 25507
rect 14993 25473 15265 25507
rect 15919 25507 16369 25529
rect 14815 25457 15265 25473
rect 15423 25471 15877 25487
rect 14319 25415 14773 25437
rect 15423 25437 15699 25471
rect 15733 25437 15877 25471
rect 15919 25473 16063 25507
rect 16097 25473 16369 25507
rect 17023 25507 17473 25529
rect 15919 25457 16369 25473
rect 16527 25471 16981 25487
rect 15423 25415 15877 25437
rect 16527 25437 16803 25471
rect 16837 25437 16981 25471
rect 17023 25473 17167 25507
rect 17201 25473 17473 25507
rect 18311 25507 18761 25529
rect 17023 25457 17473 25473
rect 17815 25471 18269 25487
rect 16527 25415 16981 25437
rect 17815 25437 18091 25471
rect 18125 25437 18269 25471
rect 18311 25473 18455 25507
rect 18489 25473 18761 25507
rect 19415 25507 19865 25529
rect 20023 25525 20141 25555
rect 18311 25457 18761 25473
rect 18919 25471 19373 25487
rect 17815 25415 18269 25437
rect 18919 25437 19195 25471
rect 19229 25437 19373 25471
rect 19415 25473 19559 25507
rect 19593 25473 19865 25507
rect 20103 25523 20141 25525
rect 20103 25507 20169 25523
rect 19415 25457 19865 25473
rect 19995 25467 20061 25483
rect 18919 25415 19373 25437
rect 19995 25433 20011 25467
rect 20045 25433 20061 25467
rect 20103 25473 20119 25507
rect 20153 25473 20169 25507
rect 20103 25457 20169 25473
rect 19995 25417 20061 25433
rect 20023 25415 20061 25417
rect 5487 25389 6065 25415
rect 6223 25389 7169 25415
rect 7511 25389 7905 25415
rect 8063 25389 9009 25415
rect 9167 25389 10113 25415
rect 10271 25389 11217 25415
rect 11375 25389 12321 25415
rect 12663 25389 13057 25415
rect 13215 25389 14161 25415
rect 14319 25389 15265 25415
rect 15423 25389 16369 25415
rect 16527 25389 17473 25415
rect 17815 25389 18761 25415
rect 18919 25389 19865 25415
rect 20023 25389 20141 25415
rect 5027 25253 5145 25279
rect 5487 25253 6065 25279
rect 6223 25253 7169 25279
rect 7511 25253 7905 25279
rect 8063 25253 9009 25279
rect 9167 25253 10113 25279
rect 10271 25253 11217 25279
rect 11375 25253 12321 25279
rect 12663 25253 13057 25279
rect 13215 25253 14161 25279
rect 14319 25253 15265 25279
rect 15423 25253 16369 25279
rect 16527 25253 17473 25279
rect 17815 25253 18761 25279
rect 18919 25253 19865 25279
rect 20023 25253 20141 25279
rect 5027 25185 5145 25211
rect 5487 25185 6433 25211
rect 6591 25185 7537 25211
rect 7695 25185 8641 25211
rect 8799 25185 9745 25211
rect 10087 25185 10481 25211
rect 10639 25185 11585 25211
rect 11743 25185 12689 25211
rect 12847 25185 13793 25211
rect 13951 25185 14897 25211
rect 15239 25185 15449 25211
rect 15607 25185 16553 25211
rect 16711 25185 17657 25211
rect 17815 25185 18761 25211
rect 18919 25185 19865 25211
rect 20023 25185 20141 25211
rect 5027 25049 5145 25075
rect 5107 25047 5145 25049
rect 5487 25049 6433 25075
rect 6591 25049 7537 25075
rect 7695 25049 8641 25075
rect 8799 25049 9745 25075
rect 10087 25049 10481 25075
rect 10639 25049 11585 25075
rect 11743 25049 12689 25075
rect 12847 25049 13793 25075
rect 13951 25049 14897 25075
rect 15239 25049 15449 25075
rect 15607 25049 16553 25075
rect 16711 25049 17657 25075
rect 17815 25049 18761 25075
rect 18919 25049 19865 25075
rect 20023 25049 20141 25075
rect 5107 25031 5173 25047
rect 4999 24991 5065 25007
rect 4999 24957 5015 24991
rect 5049 24957 5065 24991
rect 5107 24997 5123 25031
rect 5157 24997 5173 25031
rect 5107 24981 5173 24997
rect 5487 25027 5941 25049
rect 5487 24993 5763 25027
rect 5797 24993 5941 25027
rect 6591 25027 7045 25049
rect 5487 24977 5941 24993
rect 5983 24991 6433 25007
rect 4999 24941 5065 24957
rect 5027 24939 5065 24941
rect 5983 24957 6127 24991
rect 6161 24957 6433 24991
rect 6591 24993 6867 25027
rect 6901 24993 7045 25027
rect 7695 25027 8149 25049
rect 6591 24977 7045 24993
rect 7087 24991 7537 25007
rect 5027 24909 5145 24939
rect 5983 24935 6433 24957
rect 7087 24957 7231 24991
rect 7265 24957 7537 24991
rect 7695 24993 7971 25027
rect 8005 24993 8149 25027
rect 8799 25027 9253 25049
rect 7695 24977 8149 24993
rect 8191 24991 8641 25007
rect 7087 24935 7537 24957
rect 8191 24957 8335 24991
rect 8369 24957 8641 24991
rect 8799 24993 9075 25027
rect 9109 24993 9253 25027
rect 10087 25027 10263 25049
rect 8799 24977 9253 24993
rect 9295 24991 9745 25007
rect 8191 24935 8641 24957
rect 9295 24957 9439 24991
rect 9473 24957 9745 24991
rect 10087 24993 10103 25027
rect 10137 24993 10213 25027
rect 10247 24993 10263 25027
rect 10639 25027 11093 25049
rect 10087 24977 10263 24993
rect 10305 24991 10481 25007
rect 9295 24935 9745 24957
rect 10305 24957 10321 24991
rect 10355 24957 10431 24991
rect 10465 24957 10481 24991
rect 10639 24993 10915 25027
rect 10949 24993 11093 25027
rect 11743 25027 12197 25049
rect 10639 24977 11093 24993
rect 11135 24991 11585 25007
rect 10305 24935 10481 24957
rect 11135 24957 11279 24991
rect 11313 24957 11585 24991
rect 11743 24993 12019 25027
rect 12053 24993 12197 25027
rect 12847 25027 13301 25049
rect 11743 24977 12197 24993
rect 12239 24991 12689 25007
rect 11135 24935 11585 24957
rect 12239 24957 12383 24991
rect 12417 24957 12689 24991
rect 12847 24993 13123 25027
rect 13157 24993 13301 25027
rect 13951 25027 14405 25049
rect 15239 25043 15323 25049
rect 12847 24977 13301 24993
rect 13343 24991 13793 25007
rect 12239 24935 12689 24957
rect 13343 24957 13487 24991
rect 13521 24957 13793 24991
rect 13951 24993 14227 25027
rect 14261 24993 14405 25027
rect 15181 25027 15323 25043
rect 13951 24977 14405 24993
rect 14447 24991 14897 25007
rect 13343 24935 13793 24957
rect 14447 24957 14591 24991
rect 14625 24957 14897 24991
rect 15181 24993 15197 25027
rect 15231 24993 15323 25027
rect 15607 25027 16061 25049
rect 15181 24977 15323 24993
rect 15365 24991 15507 25007
rect 14447 24935 14897 24957
rect 15365 24957 15457 24991
rect 15491 24957 15507 24991
rect 15607 24993 15883 25027
rect 15917 24993 16061 25027
rect 16711 25027 17165 25049
rect 15607 24977 16061 24993
rect 16103 24991 16553 25007
rect 15365 24941 15507 24957
rect 16103 24957 16247 24991
rect 16281 24957 16553 24991
rect 16711 24993 16987 25027
rect 17021 24993 17165 25027
rect 17815 25027 18269 25049
rect 16711 24977 17165 24993
rect 17207 24991 17657 25007
rect 15365 24935 15449 24941
rect 16103 24935 16553 24957
rect 17207 24957 17351 24991
rect 17385 24957 17657 24991
rect 17815 24993 18091 25027
rect 18125 24993 18269 25027
rect 18919 25027 19373 25049
rect 20023 25047 20061 25049
rect 17815 24977 18269 24993
rect 18311 24991 18761 25007
rect 17207 24935 17657 24957
rect 18311 24957 18455 24991
rect 18489 24957 18761 24991
rect 18919 24993 19195 25027
rect 19229 24993 19373 25027
rect 19995 25031 20061 25047
rect 18919 24977 19373 24993
rect 19415 24991 19865 25007
rect 18311 24935 18761 24957
rect 19415 24957 19559 24991
rect 19593 24957 19865 24991
rect 19995 24997 20011 25031
rect 20045 24997 20061 25031
rect 19995 24981 20061 24997
rect 20103 24991 20169 25007
rect 19415 24935 19865 24957
rect 20103 24957 20119 24991
rect 20153 24957 20169 24991
rect 20103 24941 20169 24957
rect 20103 24939 20141 24941
rect 5487 24909 6433 24935
rect 6591 24909 7537 24935
rect 7695 24909 8641 24935
rect 8799 24909 9745 24935
rect 10087 24909 10481 24935
rect 10639 24909 11585 24935
rect 11743 24909 12689 24935
rect 12847 24909 13793 24935
rect 13951 24909 14897 24935
rect 15239 24909 15449 24935
rect 15607 24909 16553 24935
rect 16711 24909 17657 24935
rect 17815 24909 18761 24935
rect 18919 24909 19865 24935
rect 20023 24909 20141 24939
rect 5027 24709 5145 24735
rect 5487 24709 6433 24735
rect 6591 24709 7537 24735
rect 7695 24709 8641 24735
rect 8799 24709 9745 24735
rect 10087 24709 10481 24735
rect 10639 24709 11585 24735
rect 11743 24709 12689 24735
rect 12847 24709 13793 24735
rect 13951 24709 14897 24735
rect 15239 24709 15449 24735
rect 15607 24709 16553 24735
rect 16711 24709 17657 24735
rect 17815 24709 18761 24735
rect 18919 24709 19865 24735
rect 20023 24709 20141 24735
rect 5027 24641 5145 24667
rect 5487 24641 6065 24667
rect 6223 24641 7169 24667
rect 7511 24641 7905 24667
rect 8063 24641 9009 24667
rect 9167 24641 10113 24667
rect 10271 24641 11217 24667
rect 11375 24641 12321 24667
rect 12663 24641 13057 24667
rect 13215 24641 14161 24667
rect 14319 24641 15265 24667
rect 15423 24641 16369 24667
rect 16527 24641 17473 24667
rect 17815 24641 18761 24667
rect 18919 24641 19865 24667
rect 20023 24641 20141 24667
rect 5027 24437 5145 24467
rect 5487 24441 6065 24467
rect 6223 24441 7169 24467
rect 7511 24441 7905 24467
rect 8063 24441 9009 24467
rect 9167 24441 10113 24467
rect 10271 24441 11217 24467
rect 11375 24441 12321 24467
rect 12663 24441 13057 24467
rect 13215 24441 14161 24467
rect 14319 24441 15265 24467
rect 15423 24441 16369 24467
rect 16527 24441 17473 24467
rect 17815 24441 18761 24467
rect 18919 24441 19865 24467
rect 5027 24435 5065 24437
rect 4999 24419 5065 24435
rect 4999 24385 5015 24419
rect 5049 24385 5065 24419
rect 5801 24419 6065 24441
rect 4999 24369 5065 24385
rect 5107 24379 5173 24395
rect 5107 24345 5123 24379
rect 5157 24345 5173 24379
rect 5107 24329 5173 24345
rect 5487 24383 5759 24399
rect 5487 24349 5503 24383
rect 5537 24349 5606 24383
rect 5640 24349 5709 24383
rect 5743 24349 5759 24383
rect 5801 24385 5817 24419
rect 5851 24385 5916 24419
rect 5950 24385 6015 24419
rect 6049 24385 6065 24419
rect 6719 24419 7169 24441
rect 5801 24369 6065 24385
rect 6223 24383 6677 24399
rect 5107 24327 5145 24329
rect 5027 24301 5145 24327
rect 5487 24327 5759 24349
rect 6223 24349 6499 24383
rect 6533 24349 6677 24383
rect 6719 24385 6863 24419
rect 6897 24385 7169 24419
rect 7729 24419 7905 24441
rect 6719 24369 7169 24385
rect 7511 24383 7687 24399
rect 6223 24327 6677 24349
rect 7511 24349 7527 24383
rect 7561 24349 7637 24383
rect 7671 24349 7687 24383
rect 7729 24385 7745 24419
rect 7779 24385 7855 24419
rect 7889 24385 7905 24419
rect 8559 24419 9009 24441
rect 7729 24369 7905 24385
rect 8063 24383 8517 24399
rect 7511 24327 7687 24349
rect 8063 24349 8339 24383
rect 8373 24349 8517 24383
rect 8559 24385 8703 24419
rect 8737 24385 9009 24419
rect 9663 24419 10113 24441
rect 8559 24369 9009 24385
rect 9167 24383 9621 24399
rect 8063 24327 8517 24349
rect 9167 24349 9443 24383
rect 9477 24349 9621 24383
rect 9663 24385 9807 24419
rect 9841 24385 10113 24419
rect 10767 24419 11217 24441
rect 9663 24369 10113 24385
rect 10271 24383 10725 24399
rect 9167 24327 9621 24349
rect 10271 24349 10547 24383
rect 10581 24349 10725 24383
rect 10767 24385 10911 24419
rect 10945 24385 11217 24419
rect 11871 24419 12321 24441
rect 10767 24369 11217 24385
rect 11375 24383 11829 24399
rect 10271 24327 10725 24349
rect 11375 24349 11651 24383
rect 11685 24349 11829 24383
rect 11871 24385 12015 24419
rect 12049 24385 12321 24419
rect 12881 24419 13057 24441
rect 11871 24369 12321 24385
rect 12663 24383 12839 24399
rect 11375 24327 11829 24349
rect 12663 24349 12679 24383
rect 12713 24349 12789 24383
rect 12823 24349 12839 24383
rect 12881 24385 12897 24419
rect 12931 24385 13007 24419
rect 13041 24385 13057 24419
rect 13711 24419 14161 24441
rect 12881 24369 13057 24385
rect 13215 24383 13669 24399
rect 12663 24327 12839 24349
rect 13215 24349 13491 24383
rect 13525 24349 13669 24383
rect 13711 24385 13855 24419
rect 13889 24385 14161 24419
rect 14815 24419 15265 24441
rect 13711 24369 14161 24385
rect 14319 24383 14773 24399
rect 13215 24327 13669 24349
rect 14319 24349 14595 24383
rect 14629 24349 14773 24383
rect 14815 24385 14959 24419
rect 14993 24385 15265 24419
rect 15919 24419 16369 24441
rect 14815 24369 15265 24385
rect 15423 24383 15877 24399
rect 14319 24327 14773 24349
rect 15423 24349 15699 24383
rect 15733 24349 15877 24383
rect 15919 24385 16063 24419
rect 16097 24385 16369 24419
rect 17023 24419 17473 24441
rect 15919 24369 16369 24385
rect 16527 24383 16981 24399
rect 15423 24327 15877 24349
rect 16527 24349 16803 24383
rect 16837 24349 16981 24383
rect 17023 24385 17167 24419
rect 17201 24385 17473 24419
rect 18311 24419 18761 24441
rect 17023 24369 17473 24385
rect 17815 24383 18269 24399
rect 16527 24327 16981 24349
rect 17815 24349 18091 24383
rect 18125 24349 18269 24383
rect 18311 24385 18455 24419
rect 18489 24385 18761 24419
rect 19415 24419 19865 24441
rect 20023 24437 20141 24467
rect 18311 24369 18761 24385
rect 18919 24383 19373 24399
rect 17815 24327 18269 24349
rect 18919 24349 19195 24383
rect 19229 24349 19373 24383
rect 19415 24385 19559 24419
rect 19593 24385 19865 24419
rect 20103 24435 20141 24437
rect 20103 24419 20169 24435
rect 19415 24369 19865 24385
rect 19995 24379 20061 24395
rect 18919 24327 19373 24349
rect 19995 24345 20011 24379
rect 20045 24345 20061 24379
rect 20103 24385 20119 24419
rect 20153 24385 20169 24419
rect 20103 24369 20169 24385
rect 19995 24329 20061 24345
rect 20023 24327 20061 24329
rect 5487 24301 6065 24327
rect 6223 24301 7169 24327
rect 7511 24301 7905 24327
rect 8063 24301 9009 24327
rect 9167 24301 10113 24327
rect 10271 24301 11217 24327
rect 11375 24301 12321 24327
rect 12663 24301 13057 24327
rect 13215 24301 14161 24327
rect 14319 24301 15265 24327
rect 15423 24301 16369 24327
rect 16527 24301 17473 24327
rect 17815 24301 18761 24327
rect 18919 24301 19865 24327
rect 20023 24301 20141 24327
rect 5027 24165 5145 24191
rect 5487 24165 6065 24191
rect 6223 24165 7169 24191
rect 7511 24165 7905 24191
rect 8063 24165 9009 24191
rect 9167 24165 10113 24191
rect 10271 24165 11217 24191
rect 11375 24165 12321 24191
rect 12663 24165 13057 24191
rect 13215 24165 14161 24191
rect 14319 24165 15265 24191
rect 15423 24165 16369 24191
rect 16527 24165 17473 24191
rect 17815 24165 18761 24191
rect 18919 24165 19865 24191
rect 20023 24165 20141 24191
rect 5027 24097 5145 24123
rect 5487 24097 6433 24123
rect 6591 24097 7537 24123
rect 7695 24097 8641 24123
rect 8799 24097 9745 24123
rect 10087 24097 10481 24123
rect 10639 24097 11585 24123
rect 11743 24097 12689 24123
rect 12847 24097 13793 24123
rect 13951 24097 14897 24123
rect 15239 24097 15449 24123
rect 15607 24097 16553 24123
rect 16711 24097 17657 24123
rect 17815 24097 18761 24123
rect 18919 24097 19865 24123
rect 20023 24097 20141 24123
rect 5027 23961 5145 23987
rect 5107 23959 5145 23961
rect 5487 23961 6433 23987
rect 6591 23961 7537 23987
rect 7695 23961 8641 23987
rect 8799 23961 9745 23987
rect 10087 23961 10481 23987
rect 10639 23961 11585 23987
rect 11743 23961 12689 23987
rect 12847 23961 13793 23987
rect 13951 23961 14897 23987
rect 15239 23961 15449 23987
rect 15607 23961 16553 23987
rect 16711 23961 17657 23987
rect 17815 23961 18761 23987
rect 18919 23961 19865 23987
rect 20023 23961 20141 23987
rect 5107 23943 5173 23959
rect 4999 23903 5065 23919
rect 4999 23869 5015 23903
rect 5049 23869 5065 23903
rect 5107 23909 5123 23943
rect 5157 23909 5173 23943
rect 5107 23893 5173 23909
rect 5487 23939 5941 23961
rect 5487 23905 5763 23939
rect 5797 23905 5941 23939
rect 6591 23939 7045 23961
rect 5487 23889 5941 23905
rect 5983 23903 6433 23919
rect 4999 23853 5065 23869
rect 5027 23851 5065 23853
rect 5983 23869 6127 23903
rect 6161 23869 6433 23903
rect 6591 23905 6867 23939
rect 6901 23905 7045 23939
rect 7695 23939 8149 23961
rect 6591 23889 7045 23905
rect 7087 23903 7537 23919
rect 5027 23821 5145 23851
rect 5983 23847 6433 23869
rect 7087 23869 7231 23903
rect 7265 23869 7537 23903
rect 7695 23905 7971 23939
rect 8005 23905 8149 23939
rect 8799 23939 9253 23961
rect 7695 23889 8149 23905
rect 8191 23903 8641 23919
rect 7087 23847 7537 23869
rect 8191 23869 8335 23903
rect 8369 23869 8641 23903
rect 8799 23905 9075 23939
rect 9109 23905 9253 23939
rect 10087 23939 10263 23961
rect 8799 23889 9253 23905
rect 9295 23903 9745 23919
rect 8191 23847 8641 23869
rect 9295 23869 9439 23903
rect 9473 23869 9745 23903
rect 10087 23905 10103 23939
rect 10137 23905 10213 23939
rect 10247 23905 10263 23939
rect 10639 23939 11093 23961
rect 10087 23889 10263 23905
rect 10305 23903 10481 23919
rect 9295 23847 9745 23869
rect 10305 23869 10321 23903
rect 10355 23869 10431 23903
rect 10465 23869 10481 23903
rect 10639 23905 10915 23939
rect 10949 23905 11093 23939
rect 11743 23939 12197 23961
rect 10639 23889 11093 23905
rect 11135 23903 11585 23919
rect 10305 23847 10481 23869
rect 11135 23869 11279 23903
rect 11313 23869 11585 23903
rect 11743 23905 12019 23939
rect 12053 23905 12197 23939
rect 12847 23939 13301 23961
rect 11743 23889 12197 23905
rect 12239 23903 12689 23919
rect 11135 23847 11585 23869
rect 12239 23869 12383 23903
rect 12417 23869 12689 23903
rect 12847 23905 13123 23939
rect 13157 23905 13301 23939
rect 13951 23939 14405 23961
rect 15239 23955 15323 23961
rect 12847 23889 13301 23905
rect 13343 23903 13793 23919
rect 12239 23847 12689 23869
rect 13343 23869 13487 23903
rect 13521 23869 13793 23903
rect 13951 23905 14227 23939
rect 14261 23905 14405 23939
rect 15181 23939 15323 23955
rect 13951 23889 14405 23905
rect 14447 23903 14897 23919
rect 13343 23847 13793 23869
rect 14447 23869 14591 23903
rect 14625 23869 14897 23903
rect 15181 23905 15197 23939
rect 15231 23905 15323 23939
rect 15607 23939 16061 23961
rect 15181 23889 15323 23905
rect 15365 23903 15507 23919
rect 14447 23847 14897 23869
rect 15365 23869 15457 23903
rect 15491 23869 15507 23903
rect 15607 23905 15883 23939
rect 15917 23905 16061 23939
rect 16711 23939 17165 23961
rect 15607 23889 16061 23905
rect 16103 23903 16553 23919
rect 15365 23853 15507 23869
rect 16103 23869 16247 23903
rect 16281 23869 16553 23903
rect 16711 23905 16987 23939
rect 17021 23905 17165 23939
rect 17815 23939 18269 23961
rect 16711 23889 17165 23905
rect 17207 23903 17657 23919
rect 15365 23847 15449 23853
rect 16103 23847 16553 23869
rect 17207 23869 17351 23903
rect 17385 23869 17657 23903
rect 17815 23905 18091 23939
rect 18125 23905 18269 23939
rect 18919 23939 19373 23961
rect 20023 23959 20061 23961
rect 17815 23889 18269 23905
rect 18311 23903 18761 23919
rect 17207 23847 17657 23869
rect 18311 23869 18455 23903
rect 18489 23869 18761 23903
rect 18919 23905 19195 23939
rect 19229 23905 19373 23939
rect 19995 23943 20061 23959
rect 18919 23889 19373 23905
rect 19415 23903 19865 23919
rect 18311 23847 18761 23869
rect 19415 23869 19559 23903
rect 19593 23869 19865 23903
rect 19995 23909 20011 23943
rect 20045 23909 20061 23943
rect 19995 23893 20061 23909
rect 20103 23903 20169 23919
rect 19415 23847 19865 23869
rect 20103 23869 20119 23903
rect 20153 23869 20169 23903
rect 20103 23853 20169 23869
rect 20103 23851 20141 23853
rect 5487 23821 6433 23847
rect 6591 23821 7537 23847
rect 7695 23821 8641 23847
rect 8799 23821 9745 23847
rect 10087 23821 10481 23847
rect 10639 23821 11585 23847
rect 11743 23821 12689 23847
rect 12847 23821 13793 23847
rect 13951 23821 14897 23847
rect 15239 23821 15449 23847
rect 15607 23821 16553 23847
rect 16711 23821 17657 23847
rect 17815 23821 18761 23847
rect 18919 23821 19865 23847
rect 20023 23821 20141 23851
rect 5027 23621 5145 23647
rect 5487 23621 6433 23647
rect 6591 23621 7537 23647
rect 7695 23621 8641 23647
rect 8799 23621 9745 23647
rect 10087 23621 10481 23647
rect 10639 23621 11585 23647
rect 11743 23621 12689 23647
rect 12847 23621 13793 23647
rect 13951 23621 14897 23647
rect 15239 23621 15449 23647
rect 15607 23621 16553 23647
rect 16711 23621 17657 23647
rect 17815 23621 18761 23647
rect 18919 23621 19865 23647
rect 20023 23621 20141 23647
rect 5027 23553 5145 23579
rect 5487 23553 6065 23579
rect 6223 23553 7169 23579
rect 7511 23553 7905 23579
rect 8063 23553 9009 23579
rect 9167 23553 10113 23579
rect 10271 23553 11217 23579
rect 11375 23553 12321 23579
rect 12663 23553 13057 23579
rect 13215 23553 14161 23579
rect 14319 23553 15265 23579
rect 15423 23553 16369 23579
rect 16527 23553 17473 23579
rect 17815 23553 18761 23579
rect 18919 23553 19865 23579
rect 20023 23553 20141 23579
rect 5027 23349 5145 23379
rect 5487 23353 6065 23379
rect 6223 23353 7169 23379
rect 7511 23353 7905 23379
rect 8063 23353 9009 23379
rect 9167 23353 10113 23379
rect 10271 23353 11217 23379
rect 11375 23353 12321 23379
rect 12663 23353 13057 23379
rect 13215 23353 14161 23379
rect 14319 23353 15265 23379
rect 15423 23353 16369 23379
rect 16527 23353 17473 23379
rect 17815 23353 18761 23379
rect 18919 23353 19865 23379
rect 5027 23347 5065 23349
rect 4999 23331 5065 23347
rect 4999 23297 5015 23331
rect 5049 23297 5065 23331
rect 5801 23331 6065 23353
rect 4999 23281 5065 23297
rect 5107 23291 5173 23307
rect 5107 23257 5123 23291
rect 5157 23257 5173 23291
rect 5107 23241 5173 23257
rect 5487 23295 5759 23311
rect 5487 23261 5503 23295
rect 5537 23261 5606 23295
rect 5640 23261 5709 23295
rect 5743 23261 5759 23295
rect 5801 23297 5817 23331
rect 5851 23297 5916 23331
rect 5950 23297 6015 23331
rect 6049 23297 6065 23331
rect 6719 23331 7169 23353
rect 5801 23281 6065 23297
rect 6223 23295 6677 23311
rect 5107 23239 5145 23241
rect 5027 23213 5145 23239
rect 5487 23239 5759 23261
rect 6223 23261 6499 23295
rect 6533 23261 6677 23295
rect 6719 23297 6863 23331
rect 6897 23297 7169 23331
rect 7729 23331 7905 23353
rect 6719 23281 7169 23297
rect 7511 23295 7687 23311
rect 6223 23239 6677 23261
rect 7511 23261 7527 23295
rect 7561 23261 7637 23295
rect 7671 23261 7687 23295
rect 7729 23297 7745 23331
rect 7779 23297 7855 23331
rect 7889 23297 7905 23331
rect 8559 23331 9009 23353
rect 7729 23281 7905 23297
rect 8063 23295 8517 23311
rect 7511 23239 7687 23261
rect 8063 23261 8339 23295
rect 8373 23261 8517 23295
rect 8559 23297 8703 23331
rect 8737 23297 9009 23331
rect 9663 23331 10113 23353
rect 8559 23281 9009 23297
rect 9167 23295 9621 23311
rect 8063 23239 8517 23261
rect 9167 23261 9443 23295
rect 9477 23261 9621 23295
rect 9663 23297 9807 23331
rect 9841 23297 10113 23331
rect 10767 23331 11217 23353
rect 9663 23281 10113 23297
rect 10271 23295 10725 23311
rect 9167 23239 9621 23261
rect 10271 23261 10547 23295
rect 10581 23261 10725 23295
rect 10767 23297 10911 23331
rect 10945 23297 11217 23331
rect 11871 23331 12321 23353
rect 10767 23281 11217 23297
rect 11375 23295 11829 23311
rect 10271 23239 10725 23261
rect 11375 23261 11651 23295
rect 11685 23261 11829 23295
rect 11871 23297 12015 23331
rect 12049 23297 12321 23331
rect 12881 23331 13057 23353
rect 11871 23281 12321 23297
rect 12663 23295 12839 23311
rect 11375 23239 11829 23261
rect 12663 23261 12679 23295
rect 12713 23261 12789 23295
rect 12823 23261 12839 23295
rect 12881 23297 12897 23331
rect 12931 23297 13007 23331
rect 13041 23297 13057 23331
rect 13711 23331 14161 23353
rect 12881 23281 13057 23297
rect 13215 23295 13669 23311
rect 12663 23239 12839 23261
rect 13215 23261 13491 23295
rect 13525 23261 13669 23295
rect 13711 23297 13855 23331
rect 13889 23297 14161 23331
rect 14815 23331 15265 23353
rect 13711 23281 14161 23297
rect 14319 23295 14773 23311
rect 13215 23239 13669 23261
rect 14319 23261 14595 23295
rect 14629 23261 14773 23295
rect 14815 23297 14959 23331
rect 14993 23297 15265 23331
rect 15919 23331 16369 23353
rect 14815 23281 15265 23297
rect 15423 23295 15877 23311
rect 14319 23239 14773 23261
rect 15423 23261 15699 23295
rect 15733 23261 15877 23295
rect 15919 23297 16063 23331
rect 16097 23297 16369 23331
rect 17023 23331 17473 23353
rect 15919 23281 16369 23297
rect 16527 23295 16981 23311
rect 15423 23239 15877 23261
rect 16527 23261 16803 23295
rect 16837 23261 16981 23295
rect 17023 23297 17167 23331
rect 17201 23297 17473 23331
rect 18311 23331 18761 23353
rect 17023 23281 17473 23297
rect 17815 23295 18269 23311
rect 16527 23239 16981 23261
rect 17815 23261 18091 23295
rect 18125 23261 18269 23295
rect 18311 23297 18455 23331
rect 18489 23297 18761 23331
rect 19415 23331 19865 23353
rect 20023 23349 20141 23379
rect 18311 23281 18761 23297
rect 18919 23295 19373 23311
rect 17815 23239 18269 23261
rect 18919 23261 19195 23295
rect 19229 23261 19373 23295
rect 19415 23297 19559 23331
rect 19593 23297 19865 23331
rect 20103 23347 20141 23349
rect 20103 23331 20169 23347
rect 19415 23281 19865 23297
rect 19995 23291 20061 23307
rect 18919 23239 19373 23261
rect 19995 23257 20011 23291
rect 20045 23257 20061 23291
rect 20103 23297 20119 23331
rect 20153 23297 20169 23331
rect 20103 23281 20169 23297
rect 19995 23241 20061 23257
rect 20023 23239 20061 23241
rect 5487 23213 6065 23239
rect 6223 23213 7169 23239
rect 7511 23213 7905 23239
rect 8063 23213 9009 23239
rect 9167 23213 10113 23239
rect 10271 23213 11217 23239
rect 11375 23213 12321 23239
rect 12663 23213 13057 23239
rect 13215 23213 14161 23239
rect 14319 23213 15265 23239
rect 15423 23213 16369 23239
rect 16527 23213 17473 23239
rect 17815 23213 18761 23239
rect 18919 23213 19865 23239
rect 20023 23213 20141 23239
rect 5027 23077 5145 23103
rect 5487 23077 6065 23103
rect 6223 23077 7169 23103
rect 7511 23077 7905 23103
rect 8063 23077 9009 23103
rect 9167 23077 10113 23103
rect 10271 23077 11217 23103
rect 11375 23077 12321 23103
rect 12663 23077 13057 23103
rect 13215 23077 14161 23103
rect 14319 23077 15265 23103
rect 15423 23077 16369 23103
rect 16527 23077 17473 23103
rect 17815 23077 18761 23103
rect 18919 23077 19865 23103
rect 20023 23077 20141 23103
rect 5027 23009 5145 23035
rect 5487 23009 6433 23035
rect 6591 23009 7537 23035
rect 7695 23009 8641 23035
rect 8799 23009 9745 23035
rect 10087 23009 10481 23035
rect 10639 23009 11585 23035
rect 11743 23009 12689 23035
rect 12847 23009 13793 23035
rect 13951 23009 14897 23035
rect 15239 23009 15449 23035
rect 15607 23009 16553 23035
rect 16711 23009 17657 23035
rect 17815 23009 18761 23035
rect 18919 23009 19865 23035
rect 20023 23009 20141 23035
rect 5027 22873 5145 22899
rect 5107 22871 5145 22873
rect 5487 22873 6433 22899
rect 6591 22873 7537 22899
rect 7695 22873 8641 22899
rect 8799 22873 9745 22899
rect 10087 22873 10481 22899
rect 10639 22873 11585 22899
rect 11743 22873 12689 22899
rect 12847 22873 13793 22899
rect 13951 22873 14897 22899
rect 15239 22873 15449 22899
rect 15607 22873 16553 22899
rect 16711 22873 17657 22899
rect 17815 22873 18761 22899
rect 18919 22873 19865 22899
rect 20023 22873 20141 22899
rect 5107 22855 5173 22871
rect 4999 22815 5065 22831
rect 4999 22781 5015 22815
rect 5049 22781 5065 22815
rect 5107 22821 5123 22855
rect 5157 22821 5173 22855
rect 5107 22805 5173 22821
rect 5487 22851 5941 22873
rect 5487 22817 5763 22851
rect 5797 22817 5941 22851
rect 6591 22851 7045 22873
rect 5487 22801 5941 22817
rect 5983 22815 6433 22831
rect 4999 22765 5065 22781
rect 5027 22763 5065 22765
rect 5983 22781 6127 22815
rect 6161 22781 6433 22815
rect 6591 22817 6867 22851
rect 6901 22817 7045 22851
rect 7695 22851 8149 22873
rect 6591 22801 7045 22817
rect 7087 22815 7537 22831
rect 5027 22733 5145 22763
rect 5983 22759 6433 22781
rect 7087 22781 7231 22815
rect 7265 22781 7537 22815
rect 7695 22817 7971 22851
rect 8005 22817 8149 22851
rect 8799 22851 9253 22873
rect 7695 22801 8149 22817
rect 8191 22815 8641 22831
rect 7087 22759 7537 22781
rect 8191 22781 8335 22815
rect 8369 22781 8641 22815
rect 8799 22817 9075 22851
rect 9109 22817 9253 22851
rect 10087 22851 10263 22873
rect 8799 22801 9253 22817
rect 9295 22815 9745 22831
rect 8191 22759 8641 22781
rect 9295 22781 9439 22815
rect 9473 22781 9745 22815
rect 10087 22817 10103 22851
rect 10137 22817 10213 22851
rect 10247 22817 10263 22851
rect 10639 22851 11093 22873
rect 10087 22801 10263 22817
rect 10305 22815 10481 22831
rect 9295 22759 9745 22781
rect 10305 22781 10321 22815
rect 10355 22781 10431 22815
rect 10465 22781 10481 22815
rect 10639 22817 10915 22851
rect 10949 22817 11093 22851
rect 11743 22851 12197 22873
rect 10639 22801 11093 22817
rect 11135 22815 11585 22831
rect 10305 22759 10481 22781
rect 11135 22781 11279 22815
rect 11313 22781 11585 22815
rect 11743 22817 12019 22851
rect 12053 22817 12197 22851
rect 12847 22851 13301 22873
rect 11743 22801 12197 22817
rect 12239 22815 12689 22831
rect 11135 22759 11585 22781
rect 12239 22781 12383 22815
rect 12417 22781 12689 22815
rect 12847 22817 13123 22851
rect 13157 22817 13301 22851
rect 13951 22851 14405 22873
rect 15239 22867 15323 22873
rect 12847 22801 13301 22817
rect 13343 22815 13793 22831
rect 12239 22759 12689 22781
rect 13343 22781 13487 22815
rect 13521 22781 13793 22815
rect 13951 22817 14227 22851
rect 14261 22817 14405 22851
rect 15181 22851 15323 22867
rect 13951 22801 14405 22817
rect 14447 22815 14897 22831
rect 13343 22759 13793 22781
rect 14447 22781 14591 22815
rect 14625 22781 14897 22815
rect 15181 22817 15197 22851
rect 15231 22817 15323 22851
rect 15607 22851 16061 22873
rect 15181 22801 15323 22817
rect 15365 22815 15507 22831
rect 14447 22759 14897 22781
rect 15365 22781 15457 22815
rect 15491 22781 15507 22815
rect 15607 22817 15883 22851
rect 15917 22817 16061 22851
rect 16711 22851 17165 22873
rect 15607 22801 16061 22817
rect 16103 22815 16553 22831
rect 15365 22765 15507 22781
rect 16103 22781 16247 22815
rect 16281 22781 16553 22815
rect 16711 22817 16987 22851
rect 17021 22817 17165 22851
rect 17815 22851 18269 22873
rect 16711 22801 17165 22817
rect 17207 22815 17657 22831
rect 15365 22759 15449 22765
rect 16103 22759 16553 22781
rect 17207 22781 17351 22815
rect 17385 22781 17657 22815
rect 17815 22817 18091 22851
rect 18125 22817 18269 22851
rect 18919 22851 19373 22873
rect 20023 22871 20061 22873
rect 17815 22801 18269 22817
rect 18311 22815 18761 22831
rect 17207 22759 17657 22781
rect 18311 22781 18455 22815
rect 18489 22781 18761 22815
rect 18919 22817 19195 22851
rect 19229 22817 19373 22851
rect 19995 22855 20061 22871
rect 18919 22801 19373 22817
rect 19415 22815 19865 22831
rect 18311 22759 18761 22781
rect 19415 22781 19559 22815
rect 19593 22781 19865 22815
rect 19995 22821 20011 22855
rect 20045 22821 20061 22855
rect 19995 22805 20061 22821
rect 20103 22815 20169 22831
rect 19415 22759 19865 22781
rect 20103 22781 20119 22815
rect 20153 22781 20169 22815
rect 20103 22765 20169 22781
rect 20103 22763 20141 22765
rect 5487 22733 6433 22759
rect 6591 22733 7537 22759
rect 7695 22733 8641 22759
rect 8799 22733 9745 22759
rect 10087 22733 10481 22759
rect 10639 22733 11585 22759
rect 11743 22733 12689 22759
rect 12847 22733 13793 22759
rect 13951 22733 14897 22759
rect 15239 22733 15449 22759
rect 15607 22733 16553 22759
rect 16711 22733 17657 22759
rect 17815 22733 18761 22759
rect 18919 22733 19865 22759
rect 20023 22733 20141 22763
rect 5027 22533 5145 22559
rect 5487 22533 6433 22559
rect 6591 22533 7537 22559
rect 7695 22533 8641 22559
rect 8799 22533 9745 22559
rect 10087 22533 10481 22559
rect 10639 22533 11585 22559
rect 11743 22533 12689 22559
rect 12847 22533 13793 22559
rect 13951 22533 14897 22559
rect 15239 22533 15449 22559
rect 15607 22533 16553 22559
rect 16711 22533 17657 22559
rect 17815 22533 18761 22559
rect 18919 22533 19865 22559
rect 20023 22533 20141 22559
rect 5027 22465 5145 22491
rect 5487 22465 6065 22491
rect 6223 22465 7169 22491
rect 7511 22465 7905 22491
rect 8063 22465 9009 22491
rect 9167 22465 10113 22491
rect 10271 22465 11217 22491
rect 11375 22465 12321 22491
rect 12663 22465 13057 22491
rect 13215 22465 14161 22491
rect 14319 22465 15265 22491
rect 15423 22465 16369 22491
rect 16527 22465 17473 22491
rect 17815 22465 18761 22491
rect 18919 22465 19865 22491
rect 20023 22465 20141 22491
rect 5027 22261 5145 22291
rect 5487 22265 6065 22291
rect 6223 22265 7169 22291
rect 7511 22265 7905 22291
rect 8063 22265 9009 22291
rect 9167 22265 10113 22291
rect 10271 22265 11217 22291
rect 11375 22265 12321 22291
rect 12663 22265 13057 22291
rect 13215 22265 14161 22291
rect 14319 22265 15265 22291
rect 15423 22265 16369 22291
rect 16527 22265 17473 22291
rect 17815 22265 18761 22291
rect 18919 22265 19865 22291
rect 5027 22259 5065 22261
rect 4999 22243 5065 22259
rect 4999 22209 5015 22243
rect 5049 22209 5065 22243
rect 5801 22243 6065 22265
rect 4999 22193 5065 22209
rect 5107 22203 5173 22219
rect 5107 22169 5123 22203
rect 5157 22169 5173 22203
rect 5107 22153 5173 22169
rect 5487 22207 5759 22223
rect 5487 22173 5503 22207
rect 5537 22173 5606 22207
rect 5640 22173 5709 22207
rect 5743 22173 5759 22207
rect 5801 22209 5817 22243
rect 5851 22209 5916 22243
rect 5950 22209 6015 22243
rect 6049 22209 6065 22243
rect 6719 22243 7169 22265
rect 5801 22193 6065 22209
rect 6223 22207 6677 22223
rect 5107 22151 5145 22153
rect 5027 22125 5145 22151
rect 5487 22151 5759 22173
rect 6223 22173 6499 22207
rect 6533 22173 6677 22207
rect 6719 22209 6863 22243
rect 6897 22209 7169 22243
rect 7729 22243 7905 22265
rect 6719 22193 7169 22209
rect 7511 22207 7687 22223
rect 6223 22151 6677 22173
rect 7511 22173 7527 22207
rect 7561 22173 7637 22207
rect 7671 22173 7687 22207
rect 7729 22209 7745 22243
rect 7779 22209 7855 22243
rect 7889 22209 7905 22243
rect 8559 22243 9009 22265
rect 7729 22193 7905 22209
rect 8063 22207 8517 22223
rect 7511 22151 7687 22173
rect 8063 22173 8339 22207
rect 8373 22173 8517 22207
rect 8559 22209 8703 22243
rect 8737 22209 9009 22243
rect 9663 22243 10113 22265
rect 8559 22193 9009 22209
rect 9167 22207 9621 22223
rect 8063 22151 8517 22173
rect 9167 22173 9443 22207
rect 9477 22173 9621 22207
rect 9663 22209 9807 22243
rect 9841 22209 10113 22243
rect 10767 22243 11217 22265
rect 9663 22193 10113 22209
rect 10271 22207 10725 22223
rect 9167 22151 9621 22173
rect 10271 22173 10547 22207
rect 10581 22173 10725 22207
rect 10767 22209 10911 22243
rect 10945 22209 11217 22243
rect 11871 22243 12321 22265
rect 10767 22193 11217 22209
rect 11375 22207 11829 22223
rect 10271 22151 10725 22173
rect 11375 22173 11651 22207
rect 11685 22173 11829 22207
rect 11871 22209 12015 22243
rect 12049 22209 12321 22243
rect 12881 22243 13057 22265
rect 11871 22193 12321 22209
rect 12663 22207 12839 22223
rect 11375 22151 11829 22173
rect 12663 22173 12679 22207
rect 12713 22173 12789 22207
rect 12823 22173 12839 22207
rect 12881 22209 12897 22243
rect 12931 22209 13007 22243
rect 13041 22209 13057 22243
rect 13711 22243 14161 22265
rect 12881 22193 13057 22209
rect 13215 22207 13669 22223
rect 12663 22151 12839 22173
rect 13215 22173 13491 22207
rect 13525 22173 13669 22207
rect 13711 22209 13855 22243
rect 13889 22209 14161 22243
rect 14815 22243 15265 22265
rect 13711 22193 14161 22209
rect 14319 22207 14773 22223
rect 13215 22151 13669 22173
rect 14319 22173 14595 22207
rect 14629 22173 14773 22207
rect 14815 22209 14959 22243
rect 14993 22209 15265 22243
rect 15919 22243 16369 22265
rect 14815 22193 15265 22209
rect 15423 22207 15877 22223
rect 14319 22151 14773 22173
rect 15423 22173 15699 22207
rect 15733 22173 15877 22207
rect 15919 22209 16063 22243
rect 16097 22209 16369 22243
rect 17023 22243 17473 22265
rect 15919 22193 16369 22209
rect 16527 22207 16981 22223
rect 15423 22151 15877 22173
rect 16527 22173 16803 22207
rect 16837 22173 16981 22207
rect 17023 22209 17167 22243
rect 17201 22209 17473 22243
rect 18311 22243 18761 22265
rect 17023 22193 17473 22209
rect 17815 22207 18269 22223
rect 16527 22151 16981 22173
rect 17815 22173 18091 22207
rect 18125 22173 18269 22207
rect 18311 22209 18455 22243
rect 18489 22209 18761 22243
rect 19415 22243 19865 22265
rect 20023 22261 20141 22291
rect 18311 22193 18761 22209
rect 18919 22207 19373 22223
rect 17815 22151 18269 22173
rect 18919 22173 19195 22207
rect 19229 22173 19373 22207
rect 19415 22209 19559 22243
rect 19593 22209 19865 22243
rect 20103 22259 20141 22261
rect 20103 22243 20169 22259
rect 19415 22193 19865 22209
rect 19995 22203 20061 22219
rect 18919 22151 19373 22173
rect 19995 22169 20011 22203
rect 20045 22169 20061 22203
rect 20103 22209 20119 22243
rect 20153 22209 20169 22243
rect 20103 22193 20169 22209
rect 19995 22153 20061 22169
rect 20023 22151 20061 22153
rect 5487 22125 6065 22151
rect 6223 22125 7169 22151
rect 7511 22125 7905 22151
rect 8063 22125 9009 22151
rect 9167 22125 10113 22151
rect 10271 22125 11217 22151
rect 11375 22125 12321 22151
rect 12663 22125 13057 22151
rect 13215 22125 14161 22151
rect 14319 22125 15265 22151
rect 15423 22125 16369 22151
rect 16527 22125 17473 22151
rect 17815 22125 18761 22151
rect 18919 22125 19865 22151
rect 20023 22125 20141 22151
rect 5027 21989 5145 22015
rect 5487 21989 6065 22015
rect 6223 21989 7169 22015
rect 7511 21989 7905 22015
rect 8063 21989 9009 22015
rect 9167 21989 10113 22015
rect 10271 21989 11217 22015
rect 11375 21989 12321 22015
rect 12663 21989 13057 22015
rect 13215 21989 14161 22015
rect 14319 21989 15265 22015
rect 15423 21989 16369 22015
rect 16527 21989 17473 22015
rect 17815 21989 18761 22015
rect 18919 21989 19865 22015
rect 20023 21989 20141 22015
rect 5027 21921 5145 21947
rect 5487 21921 6433 21947
rect 6591 21921 7537 21947
rect 7695 21921 8641 21947
rect 8799 21921 9745 21947
rect 10087 21921 10481 21947
rect 10639 21921 11585 21947
rect 11743 21921 12689 21947
rect 12847 21921 13793 21947
rect 13951 21921 14897 21947
rect 15239 21921 15449 21947
rect 15607 21921 16553 21947
rect 16711 21921 17657 21947
rect 17815 21921 18761 21947
rect 18919 21921 19865 21947
rect 20023 21921 20141 21947
rect 5027 21785 5145 21811
rect 5107 21783 5145 21785
rect 5487 21785 6433 21811
rect 6591 21785 7537 21811
rect 7695 21785 8641 21811
rect 8799 21785 9745 21811
rect 10087 21785 10481 21811
rect 10639 21785 11585 21811
rect 11743 21785 12689 21811
rect 12847 21785 13793 21811
rect 13951 21785 14897 21811
rect 15239 21785 15449 21811
rect 15607 21785 16553 21811
rect 16711 21785 17657 21811
rect 17815 21785 18761 21811
rect 18919 21785 19865 21811
rect 20023 21785 20141 21811
rect 5107 21767 5173 21783
rect 4999 21727 5065 21743
rect 4999 21693 5015 21727
rect 5049 21693 5065 21727
rect 5107 21733 5123 21767
rect 5157 21733 5173 21767
rect 5107 21717 5173 21733
rect 5487 21763 5941 21785
rect 5487 21729 5763 21763
rect 5797 21729 5941 21763
rect 6591 21763 7045 21785
rect 5487 21713 5941 21729
rect 5983 21727 6433 21743
rect 4999 21677 5065 21693
rect 5027 21675 5065 21677
rect 5983 21693 6127 21727
rect 6161 21693 6433 21727
rect 6591 21729 6867 21763
rect 6901 21729 7045 21763
rect 7695 21763 8149 21785
rect 6591 21713 7045 21729
rect 7087 21727 7537 21743
rect 5027 21645 5145 21675
rect 5983 21671 6433 21693
rect 7087 21693 7231 21727
rect 7265 21693 7537 21727
rect 7695 21729 7971 21763
rect 8005 21729 8149 21763
rect 8799 21763 9253 21785
rect 7695 21713 8149 21729
rect 8191 21727 8641 21743
rect 7087 21671 7537 21693
rect 8191 21693 8335 21727
rect 8369 21693 8641 21727
rect 8799 21729 9075 21763
rect 9109 21729 9253 21763
rect 10087 21763 10263 21785
rect 8799 21713 9253 21729
rect 9295 21727 9745 21743
rect 8191 21671 8641 21693
rect 9295 21693 9439 21727
rect 9473 21693 9745 21727
rect 10087 21729 10103 21763
rect 10137 21729 10213 21763
rect 10247 21729 10263 21763
rect 10639 21763 11093 21785
rect 10087 21713 10263 21729
rect 10305 21727 10481 21743
rect 9295 21671 9745 21693
rect 10305 21693 10321 21727
rect 10355 21693 10431 21727
rect 10465 21693 10481 21727
rect 10639 21729 10915 21763
rect 10949 21729 11093 21763
rect 11743 21763 12197 21785
rect 10639 21713 11093 21729
rect 11135 21727 11585 21743
rect 10305 21671 10481 21693
rect 11135 21693 11279 21727
rect 11313 21693 11585 21727
rect 11743 21729 12019 21763
rect 12053 21729 12197 21763
rect 12847 21763 13301 21785
rect 11743 21713 12197 21729
rect 12239 21727 12689 21743
rect 11135 21671 11585 21693
rect 12239 21693 12383 21727
rect 12417 21693 12689 21727
rect 12847 21729 13123 21763
rect 13157 21729 13301 21763
rect 13951 21763 14405 21785
rect 15239 21779 15323 21785
rect 12847 21713 13301 21729
rect 13343 21727 13793 21743
rect 12239 21671 12689 21693
rect 13343 21693 13487 21727
rect 13521 21693 13793 21727
rect 13951 21729 14227 21763
rect 14261 21729 14405 21763
rect 15181 21763 15323 21779
rect 13951 21713 14405 21729
rect 14447 21727 14897 21743
rect 13343 21671 13793 21693
rect 14447 21693 14591 21727
rect 14625 21693 14897 21727
rect 15181 21729 15197 21763
rect 15231 21729 15323 21763
rect 15607 21763 16061 21785
rect 15181 21713 15323 21729
rect 15365 21727 15507 21743
rect 14447 21671 14897 21693
rect 15365 21693 15457 21727
rect 15491 21693 15507 21727
rect 15607 21729 15883 21763
rect 15917 21729 16061 21763
rect 16711 21763 17165 21785
rect 15607 21713 16061 21729
rect 16103 21727 16553 21743
rect 15365 21677 15507 21693
rect 16103 21693 16247 21727
rect 16281 21693 16553 21727
rect 16711 21729 16987 21763
rect 17021 21729 17165 21763
rect 17815 21763 18269 21785
rect 16711 21713 17165 21729
rect 17207 21727 17657 21743
rect 15365 21671 15449 21677
rect 16103 21671 16553 21693
rect 17207 21693 17351 21727
rect 17385 21693 17657 21727
rect 17815 21729 18091 21763
rect 18125 21729 18269 21763
rect 18919 21763 19373 21785
rect 20023 21783 20061 21785
rect 17815 21713 18269 21729
rect 18311 21727 18761 21743
rect 17207 21671 17657 21693
rect 18311 21693 18455 21727
rect 18489 21693 18761 21727
rect 18919 21729 19195 21763
rect 19229 21729 19373 21763
rect 19995 21767 20061 21783
rect 18919 21713 19373 21729
rect 19415 21727 19865 21743
rect 18311 21671 18761 21693
rect 19415 21693 19559 21727
rect 19593 21693 19865 21727
rect 19995 21733 20011 21767
rect 20045 21733 20061 21767
rect 19995 21717 20061 21733
rect 20103 21727 20169 21743
rect 19415 21671 19865 21693
rect 20103 21693 20119 21727
rect 20153 21693 20169 21727
rect 20103 21677 20169 21693
rect 20103 21675 20141 21677
rect 5487 21645 6433 21671
rect 6591 21645 7537 21671
rect 7695 21645 8641 21671
rect 8799 21645 9745 21671
rect 10087 21645 10481 21671
rect 10639 21645 11585 21671
rect 11743 21645 12689 21671
rect 12847 21645 13793 21671
rect 13951 21645 14897 21671
rect 15239 21645 15449 21671
rect 15607 21645 16553 21671
rect 16711 21645 17657 21671
rect 17815 21645 18761 21671
rect 18919 21645 19865 21671
rect 20023 21645 20141 21675
rect 5027 21445 5145 21471
rect 5487 21445 6433 21471
rect 6591 21445 7537 21471
rect 7695 21445 8641 21471
rect 8799 21445 9745 21471
rect 10087 21445 10481 21471
rect 10639 21445 11585 21471
rect 11743 21445 12689 21471
rect 12847 21445 13793 21471
rect 13951 21445 14897 21471
rect 15239 21445 15449 21471
rect 15607 21445 16553 21471
rect 16711 21445 17657 21471
rect 17815 21445 18761 21471
rect 18919 21445 19865 21471
rect 20023 21445 20141 21471
rect 5027 21377 5145 21403
rect 5487 21377 6065 21403
rect 6223 21377 7169 21403
rect 7511 21377 7905 21403
rect 8063 21377 9009 21403
rect 9167 21377 10113 21403
rect 10271 21377 11217 21403
rect 11375 21377 12321 21403
rect 12663 21377 13057 21403
rect 13215 21377 14161 21403
rect 14319 21377 15265 21403
rect 15423 21377 16369 21403
rect 16527 21377 17473 21403
rect 17815 21377 18761 21403
rect 18919 21377 19865 21403
rect 20023 21377 20141 21403
rect 5027 21173 5145 21203
rect 5487 21177 6065 21203
rect 6223 21177 7169 21203
rect 7511 21177 7905 21203
rect 8063 21177 9009 21203
rect 9167 21177 10113 21203
rect 10271 21177 11217 21203
rect 11375 21177 12321 21203
rect 12663 21177 13057 21203
rect 13215 21177 14161 21203
rect 14319 21177 15265 21203
rect 15423 21177 16369 21203
rect 16527 21177 17473 21203
rect 17815 21177 18761 21203
rect 18919 21177 19865 21203
rect 5027 21171 5065 21173
rect 4999 21155 5065 21171
rect 4999 21121 5015 21155
rect 5049 21121 5065 21155
rect 5801 21155 6065 21177
rect 4999 21105 5065 21121
rect 5107 21115 5173 21131
rect 5107 21081 5123 21115
rect 5157 21081 5173 21115
rect 5107 21065 5173 21081
rect 5487 21119 5759 21135
rect 5487 21085 5503 21119
rect 5537 21085 5606 21119
rect 5640 21085 5709 21119
rect 5743 21085 5759 21119
rect 5801 21121 5817 21155
rect 5851 21121 5916 21155
rect 5950 21121 6015 21155
rect 6049 21121 6065 21155
rect 6719 21155 7169 21177
rect 5801 21105 6065 21121
rect 6223 21119 6677 21135
rect 5107 21063 5145 21065
rect 5027 21037 5145 21063
rect 5487 21063 5759 21085
rect 6223 21085 6499 21119
rect 6533 21085 6677 21119
rect 6719 21121 6863 21155
rect 6897 21121 7169 21155
rect 7729 21155 7905 21177
rect 6719 21105 7169 21121
rect 7511 21119 7687 21135
rect 6223 21063 6677 21085
rect 7511 21085 7527 21119
rect 7561 21085 7637 21119
rect 7671 21085 7687 21119
rect 7729 21121 7745 21155
rect 7779 21121 7855 21155
rect 7889 21121 7905 21155
rect 8559 21155 9009 21177
rect 7729 21105 7905 21121
rect 8063 21119 8517 21135
rect 7511 21063 7687 21085
rect 8063 21085 8339 21119
rect 8373 21085 8517 21119
rect 8559 21121 8703 21155
rect 8737 21121 9009 21155
rect 9663 21155 10113 21177
rect 8559 21105 9009 21121
rect 9167 21119 9621 21135
rect 8063 21063 8517 21085
rect 9167 21085 9443 21119
rect 9477 21085 9621 21119
rect 9663 21121 9807 21155
rect 9841 21121 10113 21155
rect 10767 21155 11217 21177
rect 9663 21105 10113 21121
rect 10271 21119 10725 21135
rect 9167 21063 9621 21085
rect 10271 21085 10547 21119
rect 10581 21085 10725 21119
rect 10767 21121 10911 21155
rect 10945 21121 11217 21155
rect 11871 21155 12321 21177
rect 10767 21105 11217 21121
rect 11375 21119 11829 21135
rect 10271 21063 10725 21085
rect 11375 21085 11651 21119
rect 11685 21085 11829 21119
rect 11871 21121 12015 21155
rect 12049 21121 12321 21155
rect 12881 21155 13057 21177
rect 11871 21105 12321 21121
rect 12663 21119 12839 21135
rect 11375 21063 11829 21085
rect 12663 21085 12679 21119
rect 12713 21085 12789 21119
rect 12823 21085 12839 21119
rect 12881 21121 12897 21155
rect 12931 21121 13007 21155
rect 13041 21121 13057 21155
rect 13711 21155 14161 21177
rect 12881 21105 13057 21121
rect 13215 21119 13669 21135
rect 12663 21063 12839 21085
rect 13215 21085 13491 21119
rect 13525 21085 13669 21119
rect 13711 21121 13855 21155
rect 13889 21121 14161 21155
rect 14815 21155 15265 21177
rect 13711 21105 14161 21121
rect 14319 21119 14773 21135
rect 13215 21063 13669 21085
rect 14319 21085 14595 21119
rect 14629 21085 14773 21119
rect 14815 21121 14959 21155
rect 14993 21121 15265 21155
rect 15919 21155 16369 21177
rect 14815 21105 15265 21121
rect 15423 21119 15877 21135
rect 14319 21063 14773 21085
rect 15423 21085 15699 21119
rect 15733 21085 15877 21119
rect 15919 21121 16063 21155
rect 16097 21121 16369 21155
rect 17023 21155 17473 21177
rect 15919 21105 16369 21121
rect 16527 21119 16981 21135
rect 15423 21063 15877 21085
rect 16527 21085 16803 21119
rect 16837 21085 16981 21119
rect 17023 21121 17167 21155
rect 17201 21121 17473 21155
rect 18311 21155 18761 21177
rect 17023 21105 17473 21121
rect 17815 21119 18269 21135
rect 16527 21063 16981 21085
rect 17815 21085 18091 21119
rect 18125 21085 18269 21119
rect 18311 21121 18455 21155
rect 18489 21121 18761 21155
rect 19415 21155 19865 21177
rect 20023 21173 20141 21203
rect 18311 21105 18761 21121
rect 18919 21119 19373 21135
rect 17815 21063 18269 21085
rect 18919 21085 19195 21119
rect 19229 21085 19373 21119
rect 19415 21121 19559 21155
rect 19593 21121 19865 21155
rect 20103 21171 20141 21173
rect 20103 21155 20169 21171
rect 19415 21105 19865 21121
rect 19995 21115 20061 21131
rect 18919 21063 19373 21085
rect 19995 21081 20011 21115
rect 20045 21081 20061 21115
rect 20103 21121 20119 21155
rect 20153 21121 20169 21155
rect 20103 21105 20169 21121
rect 19995 21065 20061 21081
rect 20023 21063 20061 21065
rect 5487 21037 6065 21063
rect 6223 21037 7169 21063
rect 7511 21037 7905 21063
rect 8063 21037 9009 21063
rect 9167 21037 10113 21063
rect 10271 21037 11217 21063
rect 11375 21037 12321 21063
rect 12663 21037 13057 21063
rect 13215 21037 14161 21063
rect 14319 21037 15265 21063
rect 15423 21037 16369 21063
rect 16527 21037 17473 21063
rect 17815 21037 18761 21063
rect 18919 21037 19865 21063
rect 20023 21037 20141 21063
rect 5027 20901 5145 20927
rect 5487 20901 6065 20927
rect 6223 20901 7169 20927
rect 7511 20901 7905 20927
rect 8063 20901 9009 20927
rect 9167 20901 10113 20927
rect 10271 20901 11217 20927
rect 11375 20901 12321 20927
rect 12663 20901 13057 20927
rect 13215 20901 14161 20927
rect 14319 20901 15265 20927
rect 15423 20901 16369 20927
rect 16527 20901 17473 20927
rect 17815 20901 18761 20927
rect 18919 20901 19865 20927
rect 20023 20901 20141 20927
rect 5027 20833 5145 20859
rect 5487 20833 6433 20859
rect 6591 20833 7537 20859
rect 7695 20833 8641 20859
rect 8799 20833 9745 20859
rect 10087 20833 10481 20859
rect 10639 20833 11585 20859
rect 11743 20833 12689 20859
rect 12847 20833 13793 20859
rect 13951 20833 14897 20859
rect 15239 20833 15449 20859
rect 15607 20833 16553 20859
rect 16711 20833 17657 20859
rect 17815 20833 18761 20859
rect 18919 20833 19865 20859
rect 20023 20833 20141 20859
rect 5027 20697 5145 20723
rect 5107 20695 5145 20697
rect 5487 20697 6433 20723
rect 6591 20697 7537 20723
rect 7695 20697 8641 20723
rect 8799 20697 9745 20723
rect 10087 20697 10481 20723
rect 10639 20697 11585 20723
rect 11743 20697 12689 20723
rect 12847 20697 13793 20723
rect 13951 20697 14897 20723
rect 15239 20697 15449 20723
rect 15607 20697 16553 20723
rect 16711 20697 17657 20723
rect 17815 20697 18761 20723
rect 18919 20697 19865 20723
rect 20023 20697 20141 20723
rect 5107 20679 5173 20695
rect 4999 20639 5065 20655
rect 4999 20605 5015 20639
rect 5049 20605 5065 20639
rect 5107 20645 5123 20679
rect 5157 20645 5173 20679
rect 5107 20629 5173 20645
rect 5487 20675 5941 20697
rect 5487 20641 5763 20675
rect 5797 20641 5941 20675
rect 6591 20675 7045 20697
rect 5487 20625 5941 20641
rect 5983 20639 6433 20655
rect 4999 20589 5065 20605
rect 5027 20587 5065 20589
rect 5983 20605 6127 20639
rect 6161 20605 6433 20639
rect 6591 20641 6867 20675
rect 6901 20641 7045 20675
rect 7695 20675 8149 20697
rect 6591 20625 7045 20641
rect 7087 20639 7537 20655
rect 5027 20557 5145 20587
rect 5983 20583 6433 20605
rect 7087 20605 7231 20639
rect 7265 20605 7537 20639
rect 7695 20641 7971 20675
rect 8005 20641 8149 20675
rect 8799 20675 9253 20697
rect 7695 20625 8149 20641
rect 8191 20639 8641 20655
rect 7087 20583 7537 20605
rect 8191 20605 8335 20639
rect 8369 20605 8641 20639
rect 8799 20641 9075 20675
rect 9109 20641 9253 20675
rect 10087 20675 10263 20697
rect 8799 20625 9253 20641
rect 9295 20639 9745 20655
rect 8191 20583 8641 20605
rect 9295 20605 9439 20639
rect 9473 20605 9745 20639
rect 10087 20641 10103 20675
rect 10137 20641 10213 20675
rect 10247 20641 10263 20675
rect 10639 20675 11093 20697
rect 10087 20625 10263 20641
rect 10305 20639 10481 20655
rect 9295 20583 9745 20605
rect 10305 20605 10321 20639
rect 10355 20605 10431 20639
rect 10465 20605 10481 20639
rect 10639 20641 10915 20675
rect 10949 20641 11093 20675
rect 11743 20675 12197 20697
rect 10639 20625 11093 20641
rect 11135 20639 11585 20655
rect 10305 20583 10481 20605
rect 11135 20605 11279 20639
rect 11313 20605 11585 20639
rect 11743 20641 12019 20675
rect 12053 20641 12197 20675
rect 12847 20675 13301 20697
rect 11743 20625 12197 20641
rect 12239 20639 12689 20655
rect 11135 20583 11585 20605
rect 12239 20605 12383 20639
rect 12417 20605 12689 20639
rect 12847 20641 13123 20675
rect 13157 20641 13301 20675
rect 13951 20675 14405 20697
rect 15239 20691 15323 20697
rect 12847 20625 13301 20641
rect 13343 20639 13793 20655
rect 12239 20583 12689 20605
rect 13343 20605 13487 20639
rect 13521 20605 13793 20639
rect 13951 20641 14227 20675
rect 14261 20641 14405 20675
rect 15181 20675 15323 20691
rect 13951 20625 14405 20641
rect 14447 20639 14897 20655
rect 13343 20583 13793 20605
rect 14447 20605 14591 20639
rect 14625 20605 14897 20639
rect 15181 20641 15197 20675
rect 15231 20641 15323 20675
rect 15607 20675 16061 20697
rect 15181 20625 15323 20641
rect 15365 20639 15507 20655
rect 14447 20583 14897 20605
rect 15365 20605 15457 20639
rect 15491 20605 15507 20639
rect 15607 20641 15883 20675
rect 15917 20641 16061 20675
rect 16711 20675 17165 20697
rect 15607 20625 16061 20641
rect 16103 20639 16553 20655
rect 15365 20589 15507 20605
rect 16103 20605 16247 20639
rect 16281 20605 16553 20639
rect 16711 20641 16987 20675
rect 17021 20641 17165 20675
rect 17815 20675 18269 20697
rect 16711 20625 17165 20641
rect 17207 20639 17657 20655
rect 15365 20583 15449 20589
rect 16103 20583 16553 20605
rect 17207 20605 17351 20639
rect 17385 20605 17657 20639
rect 17815 20641 18091 20675
rect 18125 20641 18269 20675
rect 18919 20675 19373 20697
rect 20023 20695 20061 20697
rect 17815 20625 18269 20641
rect 18311 20639 18761 20655
rect 17207 20583 17657 20605
rect 18311 20605 18455 20639
rect 18489 20605 18761 20639
rect 18919 20641 19195 20675
rect 19229 20641 19373 20675
rect 19995 20679 20061 20695
rect 18919 20625 19373 20641
rect 19415 20639 19865 20655
rect 18311 20583 18761 20605
rect 19415 20605 19559 20639
rect 19593 20605 19865 20639
rect 19995 20645 20011 20679
rect 20045 20645 20061 20679
rect 19995 20629 20061 20645
rect 20103 20639 20169 20655
rect 19415 20583 19865 20605
rect 20103 20605 20119 20639
rect 20153 20605 20169 20639
rect 20103 20589 20169 20605
rect 20103 20587 20141 20589
rect 5487 20557 6433 20583
rect 6591 20557 7537 20583
rect 7695 20557 8641 20583
rect 8799 20557 9745 20583
rect 10087 20557 10481 20583
rect 10639 20557 11585 20583
rect 11743 20557 12689 20583
rect 12847 20557 13793 20583
rect 13951 20557 14897 20583
rect 15239 20557 15449 20583
rect 15607 20557 16553 20583
rect 16711 20557 17657 20583
rect 17815 20557 18761 20583
rect 18919 20557 19865 20583
rect 20023 20557 20141 20587
rect 5027 20357 5145 20383
rect 5487 20357 6433 20383
rect 6591 20357 7537 20383
rect 7695 20357 8641 20383
rect 8799 20357 9745 20383
rect 10087 20357 10481 20383
rect 10639 20357 11585 20383
rect 11743 20357 12689 20383
rect 12847 20357 13793 20383
rect 13951 20357 14897 20383
rect 15239 20357 15449 20383
rect 15607 20357 16553 20383
rect 16711 20357 17657 20383
rect 17815 20357 18761 20383
rect 18919 20357 19865 20383
rect 20023 20357 20141 20383
rect 5027 20289 5145 20315
rect 5487 20289 6065 20315
rect 6223 20289 7169 20315
rect 7511 20289 7905 20315
rect 8063 20289 9009 20315
rect 9167 20289 10113 20315
rect 10271 20289 11217 20315
rect 11375 20289 12321 20315
rect 12663 20289 13057 20315
rect 13215 20289 14161 20315
rect 14319 20289 15265 20315
rect 15423 20289 16369 20315
rect 16527 20289 17473 20315
rect 17815 20289 18761 20315
rect 18919 20289 19865 20315
rect 20023 20289 20141 20315
rect 5027 20085 5145 20115
rect 5487 20089 6065 20115
rect 6223 20089 7169 20115
rect 7511 20089 7905 20115
rect 8063 20089 9009 20115
rect 9167 20089 10113 20115
rect 10271 20089 11217 20115
rect 11375 20089 12321 20115
rect 12663 20089 13057 20115
rect 13215 20089 14161 20115
rect 14319 20089 15265 20115
rect 15423 20089 16369 20115
rect 16527 20089 17473 20115
rect 17815 20089 18761 20115
rect 18919 20089 19865 20115
rect 5027 20083 5065 20085
rect 4999 20067 5065 20083
rect 4999 20033 5015 20067
rect 5049 20033 5065 20067
rect 5801 20067 6065 20089
rect 4999 20017 5065 20033
rect 5107 20027 5173 20043
rect 5107 19993 5123 20027
rect 5157 19993 5173 20027
rect 5107 19977 5173 19993
rect 5487 20031 5759 20047
rect 5487 19997 5503 20031
rect 5537 19997 5606 20031
rect 5640 19997 5709 20031
rect 5743 19997 5759 20031
rect 5801 20033 5817 20067
rect 5851 20033 5916 20067
rect 5950 20033 6015 20067
rect 6049 20033 6065 20067
rect 6719 20067 7169 20089
rect 5801 20017 6065 20033
rect 6223 20031 6677 20047
rect 5107 19975 5145 19977
rect 5027 19949 5145 19975
rect 5487 19975 5759 19997
rect 6223 19997 6499 20031
rect 6533 19997 6677 20031
rect 6719 20033 6863 20067
rect 6897 20033 7169 20067
rect 7729 20067 7905 20089
rect 6719 20017 7169 20033
rect 7511 20031 7687 20047
rect 6223 19975 6677 19997
rect 7511 19997 7527 20031
rect 7561 19997 7637 20031
rect 7671 19997 7687 20031
rect 7729 20033 7745 20067
rect 7779 20033 7855 20067
rect 7889 20033 7905 20067
rect 8559 20067 9009 20089
rect 7729 20017 7905 20033
rect 8063 20031 8517 20047
rect 7511 19975 7687 19997
rect 8063 19997 8339 20031
rect 8373 19997 8517 20031
rect 8559 20033 8703 20067
rect 8737 20033 9009 20067
rect 9663 20067 10113 20089
rect 8559 20017 9009 20033
rect 9167 20031 9621 20047
rect 8063 19975 8517 19997
rect 9167 19997 9443 20031
rect 9477 19997 9621 20031
rect 9663 20033 9807 20067
rect 9841 20033 10113 20067
rect 10767 20067 11217 20089
rect 9663 20017 10113 20033
rect 10271 20031 10725 20047
rect 9167 19975 9621 19997
rect 10271 19997 10547 20031
rect 10581 19997 10725 20031
rect 10767 20033 10911 20067
rect 10945 20033 11217 20067
rect 11871 20067 12321 20089
rect 10767 20017 11217 20033
rect 11375 20031 11829 20047
rect 10271 19975 10725 19997
rect 11375 19997 11651 20031
rect 11685 19997 11829 20031
rect 11871 20033 12015 20067
rect 12049 20033 12321 20067
rect 12881 20067 13057 20089
rect 11871 20017 12321 20033
rect 12663 20031 12839 20047
rect 11375 19975 11829 19997
rect 12663 19997 12679 20031
rect 12713 19997 12789 20031
rect 12823 19997 12839 20031
rect 12881 20033 12897 20067
rect 12931 20033 13007 20067
rect 13041 20033 13057 20067
rect 13711 20067 14161 20089
rect 12881 20017 13057 20033
rect 13215 20031 13669 20047
rect 12663 19975 12839 19997
rect 13215 19997 13491 20031
rect 13525 19997 13669 20031
rect 13711 20033 13855 20067
rect 13889 20033 14161 20067
rect 14815 20067 15265 20089
rect 13711 20017 14161 20033
rect 14319 20031 14773 20047
rect 13215 19975 13669 19997
rect 14319 19997 14595 20031
rect 14629 19997 14773 20031
rect 14815 20033 14959 20067
rect 14993 20033 15265 20067
rect 15919 20067 16369 20089
rect 14815 20017 15265 20033
rect 15423 20031 15877 20047
rect 14319 19975 14773 19997
rect 15423 19997 15699 20031
rect 15733 19997 15877 20031
rect 15919 20033 16063 20067
rect 16097 20033 16369 20067
rect 17023 20067 17473 20089
rect 15919 20017 16369 20033
rect 16527 20031 16981 20047
rect 15423 19975 15877 19997
rect 16527 19997 16803 20031
rect 16837 19997 16981 20031
rect 17023 20033 17167 20067
rect 17201 20033 17473 20067
rect 18311 20067 18761 20089
rect 17023 20017 17473 20033
rect 17815 20031 18269 20047
rect 16527 19975 16981 19997
rect 17815 19997 18091 20031
rect 18125 19997 18269 20031
rect 18311 20033 18455 20067
rect 18489 20033 18761 20067
rect 19415 20067 19865 20089
rect 20023 20085 20141 20115
rect 18311 20017 18761 20033
rect 18919 20031 19373 20047
rect 17815 19975 18269 19997
rect 18919 19997 19195 20031
rect 19229 19997 19373 20031
rect 19415 20033 19559 20067
rect 19593 20033 19865 20067
rect 20103 20083 20141 20085
rect 20103 20067 20169 20083
rect 19415 20017 19865 20033
rect 19995 20027 20061 20043
rect 18919 19975 19373 19997
rect 19995 19993 20011 20027
rect 20045 19993 20061 20027
rect 20103 20033 20119 20067
rect 20153 20033 20169 20067
rect 20103 20017 20169 20033
rect 19995 19977 20061 19993
rect 20023 19975 20061 19977
rect 5487 19949 6065 19975
rect 6223 19949 7169 19975
rect 7511 19949 7905 19975
rect 8063 19949 9009 19975
rect 9167 19949 10113 19975
rect 10271 19949 11217 19975
rect 11375 19949 12321 19975
rect 12663 19949 13057 19975
rect 13215 19949 14161 19975
rect 14319 19949 15265 19975
rect 15423 19949 16369 19975
rect 16527 19949 17473 19975
rect 17815 19949 18761 19975
rect 18919 19949 19865 19975
rect 20023 19949 20141 19975
rect 5027 19813 5145 19839
rect 5487 19813 6065 19839
rect 6223 19813 7169 19839
rect 7511 19813 7905 19839
rect 8063 19813 9009 19839
rect 9167 19813 10113 19839
rect 10271 19813 11217 19839
rect 11375 19813 12321 19839
rect 12663 19813 13057 19839
rect 13215 19813 14161 19839
rect 14319 19813 15265 19839
rect 15423 19813 16369 19839
rect 16527 19813 17473 19839
rect 17815 19813 18761 19839
rect 18919 19813 19865 19839
rect 20023 19813 20141 19839
rect 5027 19745 5145 19771
rect 5487 19745 6433 19771
rect 6591 19745 7537 19771
rect 7695 19745 8641 19771
rect 8799 19745 9745 19771
rect 10087 19745 10481 19771
rect 10639 19745 11585 19771
rect 11743 19745 12689 19771
rect 12847 19745 13793 19771
rect 13951 19745 14897 19771
rect 15239 19745 15449 19771
rect 15607 19745 16553 19771
rect 16711 19745 17657 19771
rect 17815 19745 18761 19771
rect 18919 19745 19865 19771
rect 20023 19745 20141 19771
rect 5027 19609 5145 19635
rect 5107 19607 5145 19609
rect 5487 19609 6433 19635
rect 6591 19609 7537 19635
rect 7695 19609 8641 19635
rect 8799 19609 9745 19635
rect 10087 19609 10481 19635
rect 10639 19609 11585 19635
rect 11743 19609 12689 19635
rect 12847 19609 13793 19635
rect 13951 19609 14897 19635
rect 15239 19609 15449 19635
rect 15607 19609 16553 19635
rect 16711 19609 17657 19635
rect 17815 19609 18761 19635
rect 18919 19609 19865 19635
rect 20023 19609 20141 19635
rect 5107 19591 5173 19607
rect 4999 19551 5065 19567
rect 4999 19517 5015 19551
rect 5049 19517 5065 19551
rect 5107 19557 5123 19591
rect 5157 19557 5173 19591
rect 5107 19541 5173 19557
rect 5487 19587 5941 19609
rect 5487 19553 5763 19587
rect 5797 19553 5941 19587
rect 6591 19587 7045 19609
rect 5487 19537 5941 19553
rect 5983 19551 6433 19567
rect 4999 19501 5065 19517
rect 5027 19499 5065 19501
rect 5983 19517 6127 19551
rect 6161 19517 6433 19551
rect 6591 19553 6867 19587
rect 6901 19553 7045 19587
rect 7695 19587 8149 19609
rect 6591 19537 7045 19553
rect 7087 19551 7537 19567
rect 5027 19469 5145 19499
rect 5983 19495 6433 19517
rect 7087 19517 7231 19551
rect 7265 19517 7537 19551
rect 7695 19553 7971 19587
rect 8005 19553 8149 19587
rect 8799 19587 9253 19609
rect 7695 19537 8149 19553
rect 8191 19551 8641 19567
rect 7087 19495 7537 19517
rect 8191 19517 8335 19551
rect 8369 19517 8641 19551
rect 8799 19553 9075 19587
rect 9109 19553 9253 19587
rect 10087 19587 10263 19609
rect 8799 19537 9253 19553
rect 9295 19551 9745 19567
rect 8191 19495 8641 19517
rect 9295 19517 9439 19551
rect 9473 19517 9745 19551
rect 10087 19553 10103 19587
rect 10137 19553 10213 19587
rect 10247 19553 10263 19587
rect 10639 19587 11093 19609
rect 10087 19537 10263 19553
rect 10305 19551 10481 19567
rect 9295 19495 9745 19517
rect 10305 19517 10321 19551
rect 10355 19517 10431 19551
rect 10465 19517 10481 19551
rect 10639 19553 10915 19587
rect 10949 19553 11093 19587
rect 11743 19587 12197 19609
rect 10639 19537 11093 19553
rect 11135 19551 11585 19567
rect 10305 19495 10481 19517
rect 11135 19517 11279 19551
rect 11313 19517 11585 19551
rect 11743 19553 12019 19587
rect 12053 19553 12197 19587
rect 12847 19587 13301 19609
rect 11743 19537 12197 19553
rect 12239 19551 12689 19567
rect 11135 19495 11585 19517
rect 12239 19517 12383 19551
rect 12417 19517 12689 19551
rect 12847 19553 13123 19587
rect 13157 19553 13301 19587
rect 13951 19587 14405 19609
rect 15239 19603 15323 19609
rect 12847 19537 13301 19553
rect 13343 19551 13793 19567
rect 12239 19495 12689 19517
rect 13343 19517 13487 19551
rect 13521 19517 13793 19551
rect 13951 19553 14227 19587
rect 14261 19553 14405 19587
rect 15181 19587 15323 19603
rect 13951 19537 14405 19553
rect 14447 19551 14897 19567
rect 13343 19495 13793 19517
rect 14447 19517 14591 19551
rect 14625 19517 14897 19551
rect 15181 19553 15197 19587
rect 15231 19553 15323 19587
rect 15607 19587 16061 19609
rect 15181 19537 15323 19553
rect 15365 19551 15507 19567
rect 14447 19495 14897 19517
rect 15365 19517 15457 19551
rect 15491 19517 15507 19551
rect 15607 19553 15883 19587
rect 15917 19553 16061 19587
rect 16711 19587 17165 19609
rect 15607 19537 16061 19553
rect 16103 19551 16553 19567
rect 15365 19501 15507 19517
rect 16103 19517 16247 19551
rect 16281 19517 16553 19551
rect 16711 19553 16987 19587
rect 17021 19553 17165 19587
rect 17815 19587 18269 19609
rect 16711 19537 17165 19553
rect 17207 19551 17657 19567
rect 15365 19495 15449 19501
rect 16103 19495 16553 19517
rect 17207 19517 17351 19551
rect 17385 19517 17657 19551
rect 17815 19553 18091 19587
rect 18125 19553 18269 19587
rect 18919 19587 19373 19609
rect 20023 19607 20061 19609
rect 17815 19537 18269 19553
rect 18311 19551 18761 19567
rect 17207 19495 17657 19517
rect 18311 19517 18455 19551
rect 18489 19517 18761 19551
rect 18919 19553 19195 19587
rect 19229 19553 19373 19587
rect 19995 19591 20061 19607
rect 18919 19537 19373 19553
rect 19415 19551 19865 19567
rect 18311 19495 18761 19517
rect 19415 19517 19559 19551
rect 19593 19517 19865 19551
rect 19995 19557 20011 19591
rect 20045 19557 20061 19591
rect 19995 19541 20061 19557
rect 20103 19551 20169 19567
rect 19415 19495 19865 19517
rect 20103 19517 20119 19551
rect 20153 19517 20169 19551
rect 20103 19501 20169 19517
rect 20103 19499 20141 19501
rect 5487 19469 6433 19495
rect 6591 19469 7537 19495
rect 7695 19469 8641 19495
rect 8799 19469 9745 19495
rect 10087 19469 10481 19495
rect 10639 19469 11585 19495
rect 11743 19469 12689 19495
rect 12847 19469 13793 19495
rect 13951 19469 14897 19495
rect 15239 19469 15449 19495
rect 15607 19469 16553 19495
rect 16711 19469 17657 19495
rect 17815 19469 18761 19495
rect 18919 19469 19865 19495
rect 20023 19469 20141 19499
rect 5027 19269 5145 19295
rect 5487 19269 6433 19295
rect 6591 19269 7537 19295
rect 7695 19269 8641 19295
rect 8799 19269 9745 19295
rect 10087 19269 10481 19295
rect 10639 19269 11585 19295
rect 11743 19269 12689 19295
rect 12847 19269 13793 19295
rect 13951 19269 14897 19295
rect 15239 19269 15449 19295
rect 15607 19269 16553 19295
rect 16711 19269 17657 19295
rect 17815 19269 18761 19295
rect 18919 19269 19865 19295
rect 20023 19269 20141 19295
rect 5027 19201 5145 19227
rect 5487 19201 6065 19227
rect 6223 19201 7169 19227
rect 7511 19201 7905 19227
rect 8063 19201 9009 19227
rect 9167 19201 10113 19227
rect 10271 19201 11217 19227
rect 11375 19201 12321 19227
rect 12663 19201 13057 19227
rect 13215 19201 14161 19227
rect 14319 19201 15265 19227
rect 15423 19201 16369 19227
rect 16527 19201 17473 19227
rect 17815 19201 18761 19227
rect 18919 19201 19865 19227
rect 20023 19201 20141 19227
rect 5027 18997 5145 19027
rect 5487 19001 6065 19027
rect 6223 19001 7169 19027
rect 7511 19001 7905 19027
rect 8063 19001 9009 19027
rect 9167 19001 10113 19027
rect 10271 19001 11217 19027
rect 11375 19001 12321 19027
rect 12663 19001 13057 19027
rect 13215 19001 14161 19027
rect 14319 19001 15265 19027
rect 15423 19001 16369 19027
rect 16527 19001 17473 19027
rect 17815 19001 18761 19027
rect 18919 19001 19865 19027
rect 5027 18995 5065 18997
rect 4999 18979 5065 18995
rect 4999 18945 5015 18979
rect 5049 18945 5065 18979
rect 5801 18979 6065 19001
rect 4999 18929 5065 18945
rect 5107 18939 5173 18955
rect 5107 18905 5123 18939
rect 5157 18905 5173 18939
rect 5107 18889 5173 18905
rect 5487 18943 5759 18959
rect 5487 18909 5503 18943
rect 5537 18909 5606 18943
rect 5640 18909 5709 18943
rect 5743 18909 5759 18943
rect 5801 18945 5817 18979
rect 5851 18945 5916 18979
rect 5950 18945 6015 18979
rect 6049 18945 6065 18979
rect 6719 18979 7169 19001
rect 5801 18929 6065 18945
rect 6223 18943 6677 18959
rect 5107 18887 5145 18889
rect 5027 18861 5145 18887
rect 5487 18887 5759 18909
rect 6223 18909 6499 18943
rect 6533 18909 6677 18943
rect 6719 18945 6863 18979
rect 6897 18945 7169 18979
rect 7729 18979 7905 19001
rect 6719 18929 7169 18945
rect 7511 18943 7687 18959
rect 6223 18887 6677 18909
rect 7511 18909 7527 18943
rect 7561 18909 7637 18943
rect 7671 18909 7687 18943
rect 7729 18945 7745 18979
rect 7779 18945 7855 18979
rect 7889 18945 7905 18979
rect 8559 18979 9009 19001
rect 7729 18929 7905 18945
rect 8063 18943 8517 18959
rect 7511 18887 7687 18909
rect 8063 18909 8339 18943
rect 8373 18909 8517 18943
rect 8559 18945 8703 18979
rect 8737 18945 9009 18979
rect 9663 18979 10113 19001
rect 8559 18929 9009 18945
rect 9167 18943 9621 18959
rect 8063 18887 8517 18909
rect 9167 18909 9443 18943
rect 9477 18909 9621 18943
rect 9663 18945 9807 18979
rect 9841 18945 10113 18979
rect 10767 18979 11217 19001
rect 9663 18929 10113 18945
rect 10271 18943 10725 18959
rect 9167 18887 9621 18909
rect 10271 18909 10547 18943
rect 10581 18909 10725 18943
rect 10767 18945 10911 18979
rect 10945 18945 11217 18979
rect 11871 18979 12321 19001
rect 10767 18929 11217 18945
rect 11375 18943 11829 18959
rect 10271 18887 10725 18909
rect 11375 18909 11651 18943
rect 11685 18909 11829 18943
rect 11871 18945 12015 18979
rect 12049 18945 12321 18979
rect 12881 18979 13057 19001
rect 11871 18929 12321 18945
rect 12663 18943 12839 18959
rect 11375 18887 11829 18909
rect 12663 18909 12679 18943
rect 12713 18909 12789 18943
rect 12823 18909 12839 18943
rect 12881 18945 12897 18979
rect 12931 18945 13007 18979
rect 13041 18945 13057 18979
rect 13711 18979 14161 19001
rect 12881 18929 13057 18945
rect 13215 18943 13669 18959
rect 12663 18887 12839 18909
rect 13215 18909 13491 18943
rect 13525 18909 13669 18943
rect 13711 18945 13855 18979
rect 13889 18945 14161 18979
rect 14815 18979 15265 19001
rect 13711 18929 14161 18945
rect 14319 18943 14773 18959
rect 13215 18887 13669 18909
rect 14319 18909 14595 18943
rect 14629 18909 14773 18943
rect 14815 18945 14959 18979
rect 14993 18945 15265 18979
rect 15919 18979 16369 19001
rect 14815 18929 15265 18945
rect 15423 18943 15877 18959
rect 14319 18887 14773 18909
rect 15423 18909 15699 18943
rect 15733 18909 15877 18943
rect 15919 18945 16063 18979
rect 16097 18945 16369 18979
rect 17023 18979 17473 19001
rect 15919 18929 16369 18945
rect 16527 18943 16981 18959
rect 15423 18887 15877 18909
rect 16527 18909 16803 18943
rect 16837 18909 16981 18943
rect 17023 18945 17167 18979
rect 17201 18945 17473 18979
rect 18311 18979 18761 19001
rect 17023 18929 17473 18945
rect 17815 18943 18269 18959
rect 16527 18887 16981 18909
rect 17815 18909 18091 18943
rect 18125 18909 18269 18943
rect 18311 18945 18455 18979
rect 18489 18945 18761 18979
rect 19415 18979 19865 19001
rect 20023 18997 20141 19027
rect 18311 18929 18761 18945
rect 18919 18943 19373 18959
rect 17815 18887 18269 18909
rect 18919 18909 19195 18943
rect 19229 18909 19373 18943
rect 19415 18945 19559 18979
rect 19593 18945 19865 18979
rect 20103 18995 20141 18997
rect 20103 18979 20169 18995
rect 19415 18929 19865 18945
rect 19995 18939 20061 18955
rect 18919 18887 19373 18909
rect 19995 18905 20011 18939
rect 20045 18905 20061 18939
rect 20103 18945 20119 18979
rect 20153 18945 20169 18979
rect 20103 18929 20169 18945
rect 19995 18889 20061 18905
rect 20023 18887 20061 18889
rect 5487 18861 6065 18887
rect 6223 18861 7169 18887
rect 7511 18861 7905 18887
rect 8063 18861 9009 18887
rect 9167 18861 10113 18887
rect 10271 18861 11217 18887
rect 11375 18861 12321 18887
rect 12663 18861 13057 18887
rect 13215 18861 14161 18887
rect 14319 18861 15265 18887
rect 15423 18861 16369 18887
rect 16527 18861 17473 18887
rect 17815 18861 18761 18887
rect 18919 18861 19865 18887
rect 20023 18861 20141 18887
rect 5027 18725 5145 18751
rect 5487 18725 6065 18751
rect 6223 18725 7169 18751
rect 7511 18725 7905 18751
rect 8063 18725 9009 18751
rect 9167 18725 10113 18751
rect 10271 18725 11217 18751
rect 11375 18725 12321 18751
rect 12663 18725 13057 18751
rect 13215 18725 14161 18751
rect 14319 18725 15265 18751
rect 15423 18725 16369 18751
rect 16527 18725 17473 18751
rect 17815 18725 18761 18751
rect 18919 18725 19865 18751
rect 20023 18725 20141 18751
rect 5027 18657 5145 18683
rect 5487 18657 6433 18683
rect 6591 18657 7537 18683
rect 7695 18657 8641 18683
rect 8799 18657 9745 18683
rect 10087 18657 10481 18683
rect 10639 18657 11585 18683
rect 11743 18657 12689 18683
rect 12847 18657 13793 18683
rect 13951 18657 14897 18683
rect 15239 18657 15449 18683
rect 15607 18657 16553 18683
rect 16711 18657 17657 18683
rect 17815 18657 18761 18683
rect 18919 18657 19865 18683
rect 20023 18657 20141 18683
rect 5027 18521 5145 18547
rect 5107 18519 5145 18521
rect 5487 18521 6433 18547
rect 6591 18521 7537 18547
rect 7695 18521 8641 18547
rect 8799 18521 9745 18547
rect 10087 18521 10481 18547
rect 10639 18521 11585 18547
rect 11743 18521 12689 18547
rect 12847 18521 13793 18547
rect 13951 18521 14897 18547
rect 15239 18521 15449 18547
rect 15607 18521 16553 18547
rect 16711 18521 17657 18547
rect 17815 18521 18761 18547
rect 18919 18521 19865 18547
rect 20023 18521 20141 18547
rect 5107 18503 5173 18519
rect 4999 18463 5065 18479
rect 4999 18429 5015 18463
rect 5049 18429 5065 18463
rect 5107 18469 5123 18503
rect 5157 18469 5173 18503
rect 5107 18453 5173 18469
rect 5487 18499 5941 18521
rect 5487 18465 5763 18499
rect 5797 18465 5941 18499
rect 6591 18499 7045 18521
rect 5487 18449 5941 18465
rect 5983 18463 6433 18479
rect 4999 18413 5065 18429
rect 5027 18411 5065 18413
rect 5983 18429 6127 18463
rect 6161 18429 6433 18463
rect 6591 18465 6867 18499
rect 6901 18465 7045 18499
rect 7695 18499 8149 18521
rect 6591 18449 7045 18465
rect 7087 18463 7537 18479
rect 5027 18381 5145 18411
rect 5983 18407 6433 18429
rect 7087 18429 7231 18463
rect 7265 18429 7537 18463
rect 7695 18465 7971 18499
rect 8005 18465 8149 18499
rect 8799 18499 9253 18521
rect 7695 18449 8149 18465
rect 8191 18463 8641 18479
rect 7087 18407 7537 18429
rect 8191 18429 8335 18463
rect 8369 18429 8641 18463
rect 8799 18465 9075 18499
rect 9109 18465 9253 18499
rect 10087 18499 10263 18521
rect 8799 18449 9253 18465
rect 9295 18463 9745 18479
rect 8191 18407 8641 18429
rect 9295 18429 9439 18463
rect 9473 18429 9745 18463
rect 10087 18465 10103 18499
rect 10137 18465 10213 18499
rect 10247 18465 10263 18499
rect 10639 18499 11093 18521
rect 10087 18449 10263 18465
rect 10305 18463 10481 18479
rect 9295 18407 9745 18429
rect 10305 18429 10321 18463
rect 10355 18429 10431 18463
rect 10465 18429 10481 18463
rect 10639 18465 10915 18499
rect 10949 18465 11093 18499
rect 11743 18499 12197 18521
rect 10639 18449 11093 18465
rect 11135 18463 11585 18479
rect 10305 18407 10481 18429
rect 11135 18429 11279 18463
rect 11313 18429 11585 18463
rect 11743 18465 12019 18499
rect 12053 18465 12197 18499
rect 12847 18499 13301 18521
rect 11743 18449 12197 18465
rect 12239 18463 12689 18479
rect 11135 18407 11585 18429
rect 12239 18429 12383 18463
rect 12417 18429 12689 18463
rect 12847 18465 13123 18499
rect 13157 18465 13301 18499
rect 13951 18499 14405 18521
rect 15239 18515 15323 18521
rect 12847 18449 13301 18465
rect 13343 18463 13793 18479
rect 12239 18407 12689 18429
rect 13343 18429 13487 18463
rect 13521 18429 13793 18463
rect 13951 18465 14227 18499
rect 14261 18465 14405 18499
rect 15181 18499 15323 18515
rect 13951 18449 14405 18465
rect 14447 18463 14897 18479
rect 13343 18407 13793 18429
rect 14447 18429 14591 18463
rect 14625 18429 14897 18463
rect 15181 18465 15197 18499
rect 15231 18465 15323 18499
rect 15607 18499 16061 18521
rect 15181 18449 15323 18465
rect 15365 18463 15507 18479
rect 14447 18407 14897 18429
rect 15365 18429 15457 18463
rect 15491 18429 15507 18463
rect 15607 18465 15883 18499
rect 15917 18465 16061 18499
rect 16711 18499 17165 18521
rect 15607 18449 16061 18465
rect 16103 18463 16553 18479
rect 15365 18413 15507 18429
rect 16103 18429 16247 18463
rect 16281 18429 16553 18463
rect 16711 18465 16987 18499
rect 17021 18465 17165 18499
rect 17815 18499 18269 18521
rect 16711 18449 17165 18465
rect 17207 18463 17657 18479
rect 15365 18407 15449 18413
rect 16103 18407 16553 18429
rect 17207 18429 17351 18463
rect 17385 18429 17657 18463
rect 17815 18465 18091 18499
rect 18125 18465 18269 18499
rect 18919 18499 19373 18521
rect 20023 18519 20061 18521
rect 17815 18449 18269 18465
rect 18311 18463 18761 18479
rect 17207 18407 17657 18429
rect 18311 18429 18455 18463
rect 18489 18429 18761 18463
rect 18919 18465 19195 18499
rect 19229 18465 19373 18499
rect 19995 18503 20061 18519
rect 18919 18449 19373 18465
rect 19415 18463 19865 18479
rect 18311 18407 18761 18429
rect 19415 18429 19559 18463
rect 19593 18429 19865 18463
rect 19995 18469 20011 18503
rect 20045 18469 20061 18503
rect 19995 18453 20061 18469
rect 20103 18463 20169 18479
rect 19415 18407 19865 18429
rect 20103 18429 20119 18463
rect 20153 18429 20169 18463
rect 20103 18413 20169 18429
rect 20103 18411 20141 18413
rect 5487 18381 6433 18407
rect 6591 18381 7537 18407
rect 7695 18381 8641 18407
rect 8799 18381 9745 18407
rect 10087 18381 10481 18407
rect 10639 18381 11585 18407
rect 11743 18381 12689 18407
rect 12847 18381 13793 18407
rect 13951 18381 14897 18407
rect 15239 18381 15449 18407
rect 15607 18381 16553 18407
rect 16711 18381 17657 18407
rect 17815 18381 18761 18407
rect 18919 18381 19865 18407
rect 20023 18381 20141 18411
rect 5027 18181 5145 18207
rect 5487 18181 6433 18207
rect 6591 18181 7537 18207
rect 7695 18181 8641 18207
rect 8799 18181 9745 18207
rect 10087 18181 10481 18207
rect 10639 18181 11585 18207
rect 11743 18181 12689 18207
rect 12847 18181 13793 18207
rect 13951 18181 14897 18207
rect 15239 18181 15449 18207
rect 15607 18181 16553 18207
rect 16711 18181 17657 18207
rect 17815 18181 18761 18207
rect 18919 18181 19865 18207
rect 20023 18181 20141 18207
rect 5027 18113 5145 18139
rect 5487 18113 6065 18139
rect 6223 18113 7169 18139
rect 7511 18113 7905 18139
rect 8063 18113 9009 18139
rect 9167 18113 10113 18139
rect 10271 18113 11217 18139
rect 11375 18113 12321 18139
rect 12663 18113 13057 18139
rect 13215 18113 14161 18139
rect 14319 18113 15265 18139
rect 15423 18113 16369 18139
rect 16527 18113 17473 18139
rect 17815 18113 18761 18139
rect 18919 18113 19865 18139
rect 20023 18113 20141 18139
rect 5027 17909 5145 17939
rect 5487 17913 6065 17939
rect 6223 17913 7169 17939
rect 7511 17913 7905 17939
rect 8063 17913 9009 17939
rect 9167 17913 10113 17939
rect 10271 17913 11217 17939
rect 11375 17913 12321 17939
rect 12663 17913 13057 17939
rect 13215 17913 14161 17939
rect 14319 17913 15265 17939
rect 15423 17913 16369 17939
rect 16527 17913 17473 17939
rect 17815 17913 18761 17939
rect 18919 17913 19865 17939
rect 5027 17907 5065 17909
rect 4999 17891 5065 17907
rect 4999 17857 5015 17891
rect 5049 17857 5065 17891
rect 5801 17891 6065 17913
rect 4999 17841 5065 17857
rect 5107 17851 5173 17867
rect 5107 17817 5123 17851
rect 5157 17817 5173 17851
rect 5107 17801 5173 17817
rect 5487 17855 5759 17871
rect 5487 17821 5503 17855
rect 5537 17821 5606 17855
rect 5640 17821 5709 17855
rect 5743 17821 5759 17855
rect 5801 17857 5817 17891
rect 5851 17857 5916 17891
rect 5950 17857 6015 17891
rect 6049 17857 6065 17891
rect 6719 17891 7169 17913
rect 5801 17841 6065 17857
rect 6223 17855 6677 17871
rect 5107 17799 5145 17801
rect 5027 17773 5145 17799
rect 5487 17799 5759 17821
rect 6223 17821 6499 17855
rect 6533 17821 6677 17855
rect 6719 17857 6863 17891
rect 6897 17857 7169 17891
rect 7729 17891 7905 17913
rect 6719 17841 7169 17857
rect 7511 17855 7687 17871
rect 6223 17799 6677 17821
rect 7511 17821 7527 17855
rect 7561 17821 7637 17855
rect 7671 17821 7687 17855
rect 7729 17857 7745 17891
rect 7779 17857 7855 17891
rect 7889 17857 7905 17891
rect 8559 17891 9009 17913
rect 7729 17841 7905 17857
rect 8063 17855 8517 17871
rect 7511 17799 7687 17821
rect 8063 17821 8339 17855
rect 8373 17821 8517 17855
rect 8559 17857 8703 17891
rect 8737 17857 9009 17891
rect 9663 17891 10113 17913
rect 8559 17841 9009 17857
rect 9167 17855 9621 17871
rect 8063 17799 8517 17821
rect 9167 17821 9443 17855
rect 9477 17821 9621 17855
rect 9663 17857 9807 17891
rect 9841 17857 10113 17891
rect 10767 17891 11217 17913
rect 9663 17841 10113 17857
rect 10271 17855 10725 17871
rect 9167 17799 9621 17821
rect 10271 17821 10547 17855
rect 10581 17821 10725 17855
rect 10767 17857 10911 17891
rect 10945 17857 11217 17891
rect 11871 17891 12321 17913
rect 10767 17841 11217 17857
rect 11375 17855 11829 17871
rect 10271 17799 10725 17821
rect 11375 17821 11651 17855
rect 11685 17821 11829 17855
rect 11871 17857 12015 17891
rect 12049 17857 12321 17891
rect 12881 17891 13057 17913
rect 11871 17841 12321 17857
rect 12663 17855 12839 17871
rect 11375 17799 11829 17821
rect 12663 17821 12679 17855
rect 12713 17821 12789 17855
rect 12823 17821 12839 17855
rect 12881 17857 12897 17891
rect 12931 17857 13007 17891
rect 13041 17857 13057 17891
rect 13711 17891 14161 17913
rect 12881 17841 13057 17857
rect 13215 17855 13669 17871
rect 12663 17799 12839 17821
rect 13215 17821 13491 17855
rect 13525 17821 13669 17855
rect 13711 17857 13855 17891
rect 13889 17857 14161 17891
rect 14815 17891 15265 17913
rect 13711 17841 14161 17857
rect 14319 17855 14773 17871
rect 13215 17799 13669 17821
rect 14319 17821 14595 17855
rect 14629 17821 14773 17855
rect 14815 17857 14959 17891
rect 14993 17857 15265 17891
rect 15919 17891 16369 17913
rect 14815 17841 15265 17857
rect 15423 17855 15877 17871
rect 14319 17799 14773 17821
rect 15423 17821 15699 17855
rect 15733 17821 15877 17855
rect 15919 17857 16063 17891
rect 16097 17857 16369 17891
rect 17023 17891 17473 17913
rect 15919 17841 16369 17857
rect 16527 17855 16981 17871
rect 15423 17799 15877 17821
rect 16527 17821 16803 17855
rect 16837 17821 16981 17855
rect 17023 17857 17167 17891
rect 17201 17857 17473 17891
rect 18311 17891 18761 17913
rect 17023 17841 17473 17857
rect 17815 17855 18269 17871
rect 16527 17799 16981 17821
rect 17815 17821 18091 17855
rect 18125 17821 18269 17855
rect 18311 17857 18455 17891
rect 18489 17857 18761 17891
rect 19415 17891 19865 17913
rect 20023 17909 20141 17939
rect 18311 17841 18761 17857
rect 18919 17855 19373 17871
rect 17815 17799 18269 17821
rect 18919 17821 19195 17855
rect 19229 17821 19373 17855
rect 19415 17857 19559 17891
rect 19593 17857 19865 17891
rect 20103 17907 20141 17909
rect 20103 17891 20169 17907
rect 19415 17841 19865 17857
rect 19995 17851 20061 17867
rect 18919 17799 19373 17821
rect 19995 17817 20011 17851
rect 20045 17817 20061 17851
rect 20103 17857 20119 17891
rect 20153 17857 20169 17891
rect 20103 17841 20169 17857
rect 19995 17801 20061 17817
rect 20023 17799 20061 17801
rect 5487 17773 6065 17799
rect 6223 17773 7169 17799
rect 7511 17773 7905 17799
rect 8063 17773 9009 17799
rect 9167 17773 10113 17799
rect 10271 17773 11217 17799
rect 11375 17773 12321 17799
rect 12663 17773 13057 17799
rect 13215 17773 14161 17799
rect 14319 17773 15265 17799
rect 15423 17773 16369 17799
rect 16527 17773 17473 17799
rect 17815 17773 18761 17799
rect 18919 17773 19865 17799
rect 20023 17773 20141 17799
rect 5027 17637 5145 17663
rect 5487 17637 6065 17663
rect 6223 17637 7169 17663
rect 7511 17637 7905 17663
rect 8063 17637 9009 17663
rect 9167 17637 10113 17663
rect 10271 17637 11217 17663
rect 11375 17637 12321 17663
rect 12663 17637 13057 17663
rect 13215 17637 14161 17663
rect 14319 17637 15265 17663
rect 15423 17637 16369 17663
rect 16527 17637 17473 17663
rect 17815 17637 18761 17663
rect 18919 17637 19865 17663
rect 20023 17637 20141 17663
rect 5027 17569 5145 17595
rect 5487 17569 6433 17595
rect 6591 17569 7537 17595
rect 7695 17569 8641 17595
rect 8799 17569 9745 17595
rect 10087 17569 10481 17595
rect 10639 17569 11585 17595
rect 11743 17569 12689 17595
rect 12847 17569 13793 17595
rect 13951 17569 14897 17595
rect 15239 17569 15449 17595
rect 15607 17569 16553 17595
rect 16711 17569 17657 17595
rect 17815 17569 18761 17595
rect 18919 17569 19865 17595
rect 20023 17569 20141 17595
rect 5027 17433 5145 17459
rect 5107 17431 5145 17433
rect 5487 17433 6433 17459
rect 6591 17433 7537 17459
rect 7695 17433 8641 17459
rect 8799 17433 9745 17459
rect 10087 17433 10481 17459
rect 10639 17433 11585 17459
rect 11743 17433 12689 17459
rect 12847 17433 13793 17459
rect 13951 17433 14897 17459
rect 15239 17433 15449 17459
rect 15607 17433 16553 17459
rect 16711 17433 17657 17459
rect 17815 17433 18761 17459
rect 18919 17433 19865 17459
rect 20023 17433 20141 17459
rect 5107 17415 5173 17431
rect 4999 17375 5065 17391
rect 4999 17341 5015 17375
rect 5049 17341 5065 17375
rect 5107 17381 5123 17415
rect 5157 17381 5173 17415
rect 5107 17365 5173 17381
rect 5487 17411 5941 17433
rect 5487 17377 5763 17411
rect 5797 17377 5941 17411
rect 6591 17411 7045 17433
rect 5487 17361 5941 17377
rect 5983 17375 6433 17391
rect 4999 17325 5065 17341
rect 5027 17323 5065 17325
rect 5983 17341 6127 17375
rect 6161 17341 6433 17375
rect 6591 17377 6867 17411
rect 6901 17377 7045 17411
rect 7695 17411 8149 17433
rect 6591 17361 7045 17377
rect 7087 17375 7537 17391
rect 5027 17293 5145 17323
rect 5983 17319 6433 17341
rect 7087 17341 7231 17375
rect 7265 17341 7537 17375
rect 7695 17377 7971 17411
rect 8005 17377 8149 17411
rect 8799 17411 9253 17433
rect 7695 17361 8149 17377
rect 8191 17375 8641 17391
rect 7087 17319 7537 17341
rect 8191 17341 8335 17375
rect 8369 17341 8641 17375
rect 8799 17377 9075 17411
rect 9109 17377 9253 17411
rect 10087 17411 10263 17433
rect 8799 17361 9253 17377
rect 9295 17375 9745 17391
rect 8191 17319 8641 17341
rect 9295 17341 9439 17375
rect 9473 17341 9745 17375
rect 10087 17377 10103 17411
rect 10137 17377 10213 17411
rect 10247 17377 10263 17411
rect 10639 17411 11093 17433
rect 10087 17361 10263 17377
rect 10305 17375 10481 17391
rect 9295 17319 9745 17341
rect 10305 17341 10321 17375
rect 10355 17341 10431 17375
rect 10465 17341 10481 17375
rect 10639 17377 10915 17411
rect 10949 17377 11093 17411
rect 11743 17411 12197 17433
rect 10639 17361 11093 17377
rect 11135 17375 11585 17391
rect 10305 17319 10481 17341
rect 11135 17341 11279 17375
rect 11313 17341 11585 17375
rect 11743 17377 12019 17411
rect 12053 17377 12197 17411
rect 12847 17411 13301 17433
rect 11743 17361 12197 17377
rect 12239 17375 12689 17391
rect 11135 17319 11585 17341
rect 12239 17341 12383 17375
rect 12417 17341 12689 17375
rect 12847 17377 13123 17411
rect 13157 17377 13301 17411
rect 13951 17411 14405 17433
rect 15239 17427 15323 17433
rect 12847 17361 13301 17377
rect 13343 17375 13793 17391
rect 12239 17319 12689 17341
rect 13343 17341 13487 17375
rect 13521 17341 13793 17375
rect 13951 17377 14227 17411
rect 14261 17377 14405 17411
rect 15181 17411 15323 17427
rect 13951 17361 14405 17377
rect 14447 17375 14897 17391
rect 13343 17319 13793 17341
rect 14447 17341 14591 17375
rect 14625 17341 14897 17375
rect 15181 17377 15197 17411
rect 15231 17377 15323 17411
rect 15607 17411 16061 17433
rect 15181 17361 15323 17377
rect 15365 17375 15507 17391
rect 14447 17319 14897 17341
rect 15365 17341 15457 17375
rect 15491 17341 15507 17375
rect 15607 17377 15883 17411
rect 15917 17377 16061 17411
rect 16711 17411 17165 17433
rect 15607 17361 16061 17377
rect 16103 17375 16553 17391
rect 15365 17325 15507 17341
rect 16103 17341 16247 17375
rect 16281 17341 16553 17375
rect 16711 17377 16987 17411
rect 17021 17377 17165 17411
rect 17815 17411 18269 17433
rect 16711 17361 17165 17377
rect 17207 17375 17657 17391
rect 15365 17319 15449 17325
rect 16103 17319 16553 17341
rect 17207 17341 17351 17375
rect 17385 17341 17657 17375
rect 17815 17377 18091 17411
rect 18125 17377 18269 17411
rect 18919 17411 19373 17433
rect 20023 17431 20061 17433
rect 17815 17361 18269 17377
rect 18311 17375 18761 17391
rect 17207 17319 17657 17341
rect 18311 17341 18455 17375
rect 18489 17341 18761 17375
rect 18919 17377 19195 17411
rect 19229 17377 19373 17411
rect 19995 17415 20061 17431
rect 18919 17361 19373 17377
rect 19415 17375 19865 17391
rect 18311 17319 18761 17341
rect 19415 17341 19559 17375
rect 19593 17341 19865 17375
rect 19995 17381 20011 17415
rect 20045 17381 20061 17415
rect 19995 17365 20061 17381
rect 20103 17375 20169 17391
rect 19415 17319 19865 17341
rect 20103 17341 20119 17375
rect 20153 17341 20169 17375
rect 20103 17325 20169 17341
rect 20103 17323 20141 17325
rect 5487 17293 6433 17319
rect 6591 17293 7537 17319
rect 7695 17293 8641 17319
rect 8799 17293 9745 17319
rect 10087 17293 10481 17319
rect 10639 17293 11585 17319
rect 11743 17293 12689 17319
rect 12847 17293 13793 17319
rect 13951 17293 14897 17319
rect 15239 17293 15449 17319
rect 15607 17293 16553 17319
rect 16711 17293 17657 17319
rect 17815 17293 18761 17319
rect 18919 17293 19865 17319
rect 20023 17293 20141 17323
rect 5027 17093 5145 17119
rect 5487 17093 6433 17119
rect 6591 17093 7537 17119
rect 7695 17093 8641 17119
rect 8799 17093 9745 17119
rect 10087 17093 10481 17119
rect 10639 17093 11585 17119
rect 11743 17093 12689 17119
rect 12847 17093 13793 17119
rect 13951 17093 14897 17119
rect 15239 17093 15449 17119
rect 15607 17093 16553 17119
rect 16711 17093 17657 17119
rect 17815 17093 18761 17119
rect 18919 17093 19865 17119
rect 20023 17093 20141 17119
rect 5027 17025 5145 17051
rect 5487 17025 6065 17051
rect 6223 17025 7169 17051
rect 7511 17025 7905 17051
rect 8063 17025 9009 17051
rect 9167 17025 10113 17051
rect 10271 17025 11217 17051
rect 11375 17025 12321 17051
rect 12663 17025 13057 17051
rect 13215 17025 14161 17051
rect 14319 17025 15265 17051
rect 15423 17025 16369 17051
rect 16527 17025 17473 17051
rect 17815 17025 18761 17051
rect 18919 17025 19865 17051
rect 20023 17025 20141 17051
rect 5027 16821 5145 16851
rect 5487 16825 6065 16851
rect 6223 16825 7169 16851
rect 7511 16825 7905 16851
rect 8063 16825 9009 16851
rect 9167 16825 10113 16851
rect 10271 16825 11217 16851
rect 11375 16825 12321 16851
rect 12663 16825 13057 16851
rect 13215 16825 14161 16851
rect 14319 16825 15265 16851
rect 15423 16825 16369 16851
rect 16527 16825 17473 16851
rect 17815 16825 18761 16851
rect 18919 16825 19865 16851
rect 5027 16819 5065 16821
rect 4999 16803 5065 16819
rect 4999 16769 5015 16803
rect 5049 16769 5065 16803
rect 5801 16803 6065 16825
rect 4999 16753 5065 16769
rect 5107 16763 5173 16779
rect 5107 16729 5123 16763
rect 5157 16729 5173 16763
rect 5107 16713 5173 16729
rect 5487 16767 5759 16783
rect 5487 16733 5503 16767
rect 5537 16733 5606 16767
rect 5640 16733 5709 16767
rect 5743 16733 5759 16767
rect 5801 16769 5817 16803
rect 5851 16769 5916 16803
rect 5950 16769 6015 16803
rect 6049 16769 6065 16803
rect 6719 16803 7169 16825
rect 5801 16753 6065 16769
rect 6223 16767 6677 16783
rect 5107 16711 5145 16713
rect 5027 16685 5145 16711
rect 5487 16711 5759 16733
rect 6223 16733 6499 16767
rect 6533 16733 6677 16767
rect 6719 16769 6863 16803
rect 6897 16769 7169 16803
rect 7729 16803 7905 16825
rect 6719 16753 7169 16769
rect 7511 16767 7687 16783
rect 6223 16711 6677 16733
rect 7511 16733 7527 16767
rect 7561 16733 7637 16767
rect 7671 16733 7687 16767
rect 7729 16769 7745 16803
rect 7779 16769 7855 16803
rect 7889 16769 7905 16803
rect 8559 16803 9009 16825
rect 7729 16753 7905 16769
rect 8063 16767 8517 16783
rect 7511 16711 7687 16733
rect 8063 16733 8339 16767
rect 8373 16733 8517 16767
rect 8559 16769 8703 16803
rect 8737 16769 9009 16803
rect 9663 16803 10113 16825
rect 8559 16753 9009 16769
rect 9167 16767 9621 16783
rect 8063 16711 8517 16733
rect 9167 16733 9443 16767
rect 9477 16733 9621 16767
rect 9663 16769 9807 16803
rect 9841 16769 10113 16803
rect 10767 16803 11217 16825
rect 9663 16753 10113 16769
rect 10271 16767 10725 16783
rect 9167 16711 9621 16733
rect 10271 16733 10547 16767
rect 10581 16733 10725 16767
rect 10767 16769 10911 16803
rect 10945 16769 11217 16803
rect 11871 16803 12321 16825
rect 10767 16753 11217 16769
rect 11375 16767 11829 16783
rect 10271 16711 10725 16733
rect 11375 16733 11651 16767
rect 11685 16733 11829 16767
rect 11871 16769 12015 16803
rect 12049 16769 12321 16803
rect 12881 16803 13057 16825
rect 11871 16753 12321 16769
rect 12663 16767 12839 16783
rect 11375 16711 11829 16733
rect 12663 16733 12679 16767
rect 12713 16733 12789 16767
rect 12823 16733 12839 16767
rect 12881 16769 12897 16803
rect 12931 16769 13007 16803
rect 13041 16769 13057 16803
rect 13711 16803 14161 16825
rect 12881 16753 13057 16769
rect 13215 16767 13669 16783
rect 12663 16711 12839 16733
rect 13215 16733 13491 16767
rect 13525 16733 13669 16767
rect 13711 16769 13855 16803
rect 13889 16769 14161 16803
rect 14815 16803 15265 16825
rect 13711 16753 14161 16769
rect 14319 16767 14773 16783
rect 13215 16711 13669 16733
rect 14319 16733 14595 16767
rect 14629 16733 14773 16767
rect 14815 16769 14959 16803
rect 14993 16769 15265 16803
rect 15919 16803 16369 16825
rect 14815 16753 15265 16769
rect 15423 16767 15877 16783
rect 14319 16711 14773 16733
rect 15423 16733 15699 16767
rect 15733 16733 15877 16767
rect 15919 16769 16063 16803
rect 16097 16769 16369 16803
rect 17023 16803 17473 16825
rect 15919 16753 16369 16769
rect 16527 16767 16981 16783
rect 15423 16711 15877 16733
rect 16527 16733 16803 16767
rect 16837 16733 16981 16767
rect 17023 16769 17167 16803
rect 17201 16769 17473 16803
rect 18311 16803 18761 16825
rect 17023 16753 17473 16769
rect 17815 16767 18269 16783
rect 16527 16711 16981 16733
rect 17815 16733 18091 16767
rect 18125 16733 18269 16767
rect 18311 16769 18455 16803
rect 18489 16769 18761 16803
rect 19415 16803 19865 16825
rect 20023 16821 20141 16851
rect 18311 16753 18761 16769
rect 18919 16767 19373 16783
rect 17815 16711 18269 16733
rect 18919 16733 19195 16767
rect 19229 16733 19373 16767
rect 19415 16769 19559 16803
rect 19593 16769 19865 16803
rect 20103 16819 20141 16821
rect 20103 16803 20169 16819
rect 19415 16753 19865 16769
rect 19995 16763 20061 16779
rect 18919 16711 19373 16733
rect 19995 16729 20011 16763
rect 20045 16729 20061 16763
rect 20103 16769 20119 16803
rect 20153 16769 20169 16803
rect 20103 16753 20169 16769
rect 19995 16713 20061 16729
rect 20023 16711 20061 16713
rect 5487 16685 6065 16711
rect 6223 16685 7169 16711
rect 7511 16685 7905 16711
rect 8063 16685 9009 16711
rect 9167 16685 10113 16711
rect 10271 16685 11217 16711
rect 11375 16685 12321 16711
rect 12663 16685 13057 16711
rect 13215 16685 14161 16711
rect 14319 16685 15265 16711
rect 15423 16685 16369 16711
rect 16527 16685 17473 16711
rect 17815 16685 18761 16711
rect 18919 16685 19865 16711
rect 20023 16685 20141 16711
rect 5027 16549 5145 16575
rect 5487 16549 6065 16575
rect 6223 16549 7169 16575
rect 7511 16549 7905 16575
rect 8063 16549 9009 16575
rect 9167 16549 10113 16575
rect 10271 16549 11217 16575
rect 11375 16549 12321 16575
rect 12663 16549 13057 16575
rect 13215 16549 14161 16575
rect 14319 16549 15265 16575
rect 15423 16549 16369 16575
rect 16527 16549 17473 16575
rect 17815 16549 18761 16575
rect 18919 16549 19865 16575
rect 20023 16549 20141 16575
rect 5027 16481 5145 16507
rect 5487 16481 6433 16507
rect 6591 16481 7537 16507
rect 7695 16481 8641 16507
rect 8799 16481 9745 16507
rect 10087 16481 10481 16507
rect 10639 16481 11585 16507
rect 11743 16481 12689 16507
rect 12847 16481 13793 16507
rect 13951 16481 14897 16507
rect 15239 16481 15449 16507
rect 15607 16481 16553 16507
rect 16711 16481 17657 16507
rect 17815 16481 18761 16507
rect 18919 16481 19865 16507
rect 20023 16481 20141 16507
rect 5027 16345 5145 16371
rect 5107 16343 5145 16345
rect 5487 16345 6433 16371
rect 6591 16345 7537 16371
rect 7695 16345 8641 16371
rect 8799 16345 9745 16371
rect 10087 16345 10481 16371
rect 10639 16345 11585 16371
rect 11743 16345 12689 16371
rect 12847 16345 13793 16371
rect 13951 16345 14897 16371
rect 15239 16345 15449 16371
rect 15607 16345 16553 16371
rect 16711 16345 17657 16371
rect 17815 16345 18761 16371
rect 18919 16345 19865 16371
rect 20023 16345 20141 16371
rect 5107 16327 5173 16343
rect 4999 16287 5065 16303
rect 4999 16253 5015 16287
rect 5049 16253 5065 16287
rect 5107 16293 5123 16327
rect 5157 16293 5173 16327
rect 5107 16277 5173 16293
rect 5487 16323 5941 16345
rect 5487 16289 5763 16323
rect 5797 16289 5941 16323
rect 6591 16323 7045 16345
rect 5487 16273 5941 16289
rect 5983 16287 6433 16303
rect 4999 16237 5065 16253
rect 5027 16235 5065 16237
rect 5983 16253 6127 16287
rect 6161 16253 6433 16287
rect 6591 16289 6867 16323
rect 6901 16289 7045 16323
rect 7695 16323 8149 16345
rect 6591 16273 7045 16289
rect 7087 16287 7537 16303
rect 5027 16205 5145 16235
rect 5983 16231 6433 16253
rect 7087 16253 7231 16287
rect 7265 16253 7537 16287
rect 7695 16289 7971 16323
rect 8005 16289 8149 16323
rect 8799 16323 9253 16345
rect 7695 16273 8149 16289
rect 8191 16287 8641 16303
rect 7087 16231 7537 16253
rect 8191 16253 8335 16287
rect 8369 16253 8641 16287
rect 8799 16289 9075 16323
rect 9109 16289 9253 16323
rect 10087 16323 10263 16345
rect 8799 16273 9253 16289
rect 9295 16287 9745 16303
rect 8191 16231 8641 16253
rect 9295 16253 9439 16287
rect 9473 16253 9745 16287
rect 10087 16289 10103 16323
rect 10137 16289 10213 16323
rect 10247 16289 10263 16323
rect 10639 16323 11093 16345
rect 10087 16273 10263 16289
rect 10305 16287 10481 16303
rect 9295 16231 9745 16253
rect 10305 16253 10321 16287
rect 10355 16253 10431 16287
rect 10465 16253 10481 16287
rect 10639 16289 10915 16323
rect 10949 16289 11093 16323
rect 11743 16323 12197 16345
rect 10639 16273 11093 16289
rect 11135 16287 11585 16303
rect 10305 16231 10481 16253
rect 11135 16253 11279 16287
rect 11313 16253 11585 16287
rect 11743 16289 12019 16323
rect 12053 16289 12197 16323
rect 12847 16323 13301 16345
rect 11743 16273 12197 16289
rect 12239 16287 12689 16303
rect 11135 16231 11585 16253
rect 12239 16253 12383 16287
rect 12417 16253 12689 16287
rect 12847 16289 13123 16323
rect 13157 16289 13301 16323
rect 13951 16323 14405 16345
rect 15239 16339 15323 16345
rect 12847 16273 13301 16289
rect 13343 16287 13793 16303
rect 12239 16231 12689 16253
rect 13343 16253 13487 16287
rect 13521 16253 13793 16287
rect 13951 16289 14227 16323
rect 14261 16289 14405 16323
rect 15181 16323 15323 16339
rect 13951 16273 14405 16289
rect 14447 16287 14897 16303
rect 13343 16231 13793 16253
rect 14447 16253 14591 16287
rect 14625 16253 14897 16287
rect 15181 16289 15197 16323
rect 15231 16289 15323 16323
rect 15607 16323 16061 16345
rect 15181 16273 15323 16289
rect 15365 16287 15507 16303
rect 14447 16231 14897 16253
rect 15365 16253 15457 16287
rect 15491 16253 15507 16287
rect 15607 16289 15883 16323
rect 15917 16289 16061 16323
rect 16711 16323 17165 16345
rect 15607 16273 16061 16289
rect 16103 16287 16553 16303
rect 15365 16237 15507 16253
rect 16103 16253 16247 16287
rect 16281 16253 16553 16287
rect 16711 16289 16987 16323
rect 17021 16289 17165 16323
rect 17815 16323 18269 16345
rect 16711 16273 17165 16289
rect 17207 16287 17657 16303
rect 15365 16231 15449 16237
rect 16103 16231 16553 16253
rect 17207 16253 17351 16287
rect 17385 16253 17657 16287
rect 17815 16289 18091 16323
rect 18125 16289 18269 16323
rect 18919 16323 19373 16345
rect 20023 16343 20061 16345
rect 17815 16273 18269 16289
rect 18311 16287 18761 16303
rect 17207 16231 17657 16253
rect 18311 16253 18455 16287
rect 18489 16253 18761 16287
rect 18919 16289 19195 16323
rect 19229 16289 19373 16323
rect 19995 16327 20061 16343
rect 18919 16273 19373 16289
rect 19415 16287 19865 16303
rect 18311 16231 18761 16253
rect 19415 16253 19559 16287
rect 19593 16253 19865 16287
rect 19995 16293 20011 16327
rect 20045 16293 20061 16327
rect 19995 16277 20061 16293
rect 20103 16287 20169 16303
rect 19415 16231 19865 16253
rect 20103 16253 20119 16287
rect 20153 16253 20169 16287
rect 20103 16237 20169 16253
rect 20103 16235 20141 16237
rect 5487 16205 6433 16231
rect 6591 16205 7537 16231
rect 7695 16205 8641 16231
rect 8799 16205 9745 16231
rect 10087 16205 10481 16231
rect 10639 16205 11585 16231
rect 11743 16205 12689 16231
rect 12847 16205 13793 16231
rect 13951 16205 14897 16231
rect 15239 16205 15449 16231
rect 15607 16205 16553 16231
rect 16711 16205 17657 16231
rect 17815 16205 18761 16231
rect 18919 16205 19865 16231
rect 20023 16205 20141 16235
rect 5027 16005 5145 16031
rect 5487 16005 6433 16031
rect 6591 16005 7537 16031
rect 7695 16005 8641 16031
rect 8799 16005 9745 16031
rect 10087 16005 10481 16031
rect 10639 16005 11585 16031
rect 11743 16005 12689 16031
rect 12847 16005 13793 16031
rect 13951 16005 14897 16031
rect 15239 16005 15449 16031
rect 15607 16005 16553 16031
rect 16711 16005 17657 16031
rect 17815 16005 18761 16031
rect 18919 16005 19865 16031
rect 20023 16005 20141 16031
rect 5027 15937 5145 15963
rect 5487 15937 6065 15963
rect 6223 15937 7169 15963
rect 7511 15937 7905 15963
rect 8063 15937 9009 15963
rect 9167 15937 10113 15963
rect 10271 15937 11217 15963
rect 11375 15937 12321 15963
rect 12663 15937 13057 15963
rect 13215 15937 14161 15963
rect 14319 15937 15265 15963
rect 15423 15937 16369 15963
rect 16527 15937 17473 15963
rect 17815 15937 18761 15963
rect 18919 15937 19865 15963
rect 20023 15937 20141 15963
rect 5027 15733 5145 15763
rect 5487 15737 6065 15763
rect 6223 15737 7169 15763
rect 7511 15737 7905 15763
rect 8063 15737 9009 15763
rect 9167 15737 10113 15763
rect 10271 15737 11217 15763
rect 11375 15737 12321 15763
rect 12663 15737 13057 15763
rect 13215 15737 14161 15763
rect 14319 15737 15265 15763
rect 15423 15737 16369 15763
rect 16527 15737 17473 15763
rect 17815 15737 18761 15763
rect 18919 15737 19865 15763
rect 5027 15731 5065 15733
rect 4999 15715 5065 15731
rect 4999 15681 5015 15715
rect 5049 15681 5065 15715
rect 5801 15715 6065 15737
rect 4999 15665 5065 15681
rect 5107 15675 5173 15691
rect 5107 15641 5123 15675
rect 5157 15641 5173 15675
rect 5107 15625 5173 15641
rect 5487 15679 5759 15695
rect 5487 15645 5503 15679
rect 5537 15645 5606 15679
rect 5640 15645 5709 15679
rect 5743 15645 5759 15679
rect 5801 15681 5817 15715
rect 5851 15681 5916 15715
rect 5950 15681 6015 15715
rect 6049 15681 6065 15715
rect 6719 15715 7169 15737
rect 5801 15665 6065 15681
rect 6223 15679 6677 15695
rect 5107 15623 5145 15625
rect 5027 15597 5145 15623
rect 5487 15623 5759 15645
rect 6223 15645 6499 15679
rect 6533 15645 6677 15679
rect 6719 15681 6863 15715
rect 6897 15681 7169 15715
rect 7729 15715 7905 15737
rect 6719 15665 7169 15681
rect 7511 15679 7687 15695
rect 6223 15623 6677 15645
rect 7511 15645 7527 15679
rect 7561 15645 7637 15679
rect 7671 15645 7687 15679
rect 7729 15681 7745 15715
rect 7779 15681 7855 15715
rect 7889 15681 7905 15715
rect 8559 15715 9009 15737
rect 7729 15665 7905 15681
rect 8063 15679 8517 15695
rect 7511 15623 7687 15645
rect 8063 15645 8339 15679
rect 8373 15645 8517 15679
rect 8559 15681 8703 15715
rect 8737 15681 9009 15715
rect 9663 15715 10113 15737
rect 8559 15665 9009 15681
rect 9167 15679 9621 15695
rect 8063 15623 8517 15645
rect 9167 15645 9443 15679
rect 9477 15645 9621 15679
rect 9663 15681 9807 15715
rect 9841 15681 10113 15715
rect 10767 15715 11217 15737
rect 9663 15665 10113 15681
rect 10271 15679 10725 15695
rect 9167 15623 9621 15645
rect 10271 15645 10547 15679
rect 10581 15645 10725 15679
rect 10767 15681 10911 15715
rect 10945 15681 11217 15715
rect 11871 15715 12321 15737
rect 10767 15665 11217 15681
rect 11375 15679 11829 15695
rect 10271 15623 10725 15645
rect 11375 15645 11651 15679
rect 11685 15645 11829 15679
rect 11871 15681 12015 15715
rect 12049 15681 12321 15715
rect 12881 15715 13057 15737
rect 11871 15665 12321 15681
rect 12663 15679 12839 15695
rect 11375 15623 11829 15645
rect 12663 15645 12679 15679
rect 12713 15645 12789 15679
rect 12823 15645 12839 15679
rect 12881 15681 12897 15715
rect 12931 15681 13007 15715
rect 13041 15681 13057 15715
rect 13711 15715 14161 15737
rect 12881 15665 13057 15681
rect 13215 15679 13669 15695
rect 12663 15623 12839 15645
rect 13215 15645 13491 15679
rect 13525 15645 13669 15679
rect 13711 15681 13855 15715
rect 13889 15681 14161 15715
rect 14815 15715 15265 15737
rect 13711 15665 14161 15681
rect 14319 15679 14773 15695
rect 13215 15623 13669 15645
rect 14319 15645 14595 15679
rect 14629 15645 14773 15679
rect 14815 15681 14959 15715
rect 14993 15681 15265 15715
rect 15919 15715 16369 15737
rect 14815 15665 15265 15681
rect 15423 15679 15877 15695
rect 14319 15623 14773 15645
rect 15423 15645 15699 15679
rect 15733 15645 15877 15679
rect 15919 15681 16063 15715
rect 16097 15681 16369 15715
rect 17023 15715 17473 15737
rect 15919 15665 16369 15681
rect 16527 15679 16981 15695
rect 15423 15623 15877 15645
rect 16527 15645 16803 15679
rect 16837 15645 16981 15679
rect 17023 15681 17167 15715
rect 17201 15681 17473 15715
rect 18311 15715 18761 15737
rect 17023 15665 17473 15681
rect 17815 15679 18269 15695
rect 16527 15623 16981 15645
rect 17815 15645 18091 15679
rect 18125 15645 18269 15679
rect 18311 15681 18455 15715
rect 18489 15681 18761 15715
rect 19415 15715 19865 15737
rect 20023 15733 20141 15763
rect 18311 15665 18761 15681
rect 18919 15679 19373 15695
rect 17815 15623 18269 15645
rect 18919 15645 19195 15679
rect 19229 15645 19373 15679
rect 19415 15681 19559 15715
rect 19593 15681 19865 15715
rect 20103 15731 20141 15733
rect 20103 15715 20169 15731
rect 19415 15665 19865 15681
rect 19995 15675 20061 15691
rect 18919 15623 19373 15645
rect 19995 15641 20011 15675
rect 20045 15641 20061 15675
rect 20103 15681 20119 15715
rect 20153 15681 20169 15715
rect 20103 15665 20169 15681
rect 19995 15625 20061 15641
rect 20023 15623 20061 15625
rect 5487 15597 6065 15623
rect 6223 15597 7169 15623
rect 7511 15597 7905 15623
rect 8063 15597 9009 15623
rect 9167 15597 10113 15623
rect 10271 15597 11217 15623
rect 11375 15597 12321 15623
rect 12663 15597 13057 15623
rect 13215 15597 14161 15623
rect 14319 15597 15265 15623
rect 15423 15597 16369 15623
rect 16527 15597 17473 15623
rect 17815 15597 18761 15623
rect 18919 15597 19865 15623
rect 20023 15597 20141 15623
rect 5027 15461 5145 15487
rect 5487 15461 6065 15487
rect 6223 15461 7169 15487
rect 7511 15461 7905 15487
rect 8063 15461 9009 15487
rect 9167 15461 10113 15487
rect 10271 15461 11217 15487
rect 11375 15461 12321 15487
rect 12663 15461 13057 15487
rect 13215 15461 14161 15487
rect 14319 15461 15265 15487
rect 15423 15461 16369 15487
rect 16527 15461 17473 15487
rect 17815 15461 18761 15487
rect 18919 15461 19865 15487
rect 20023 15461 20141 15487
rect 5027 15393 5145 15419
rect 5487 15393 6433 15419
rect 6591 15393 7537 15419
rect 7695 15393 8641 15419
rect 8799 15393 9745 15419
rect 10087 15393 10481 15419
rect 10639 15393 11585 15419
rect 11743 15393 12689 15419
rect 12869 15393 12899 15419
rect 12953 15393 13053 15419
rect 13211 15393 13311 15419
rect 13376 15393 13406 15419
rect 13583 15393 13793 15419
rect 13951 15393 14897 15419
rect 15147 15393 15265 15419
rect 15445 15393 15475 15419
rect 15529 15393 15629 15419
rect 15787 15393 15887 15419
rect 15952 15393 15982 15419
rect 16159 15393 16553 15419
rect 16711 15393 17657 15419
rect 17815 15393 18761 15419
rect 18919 15393 19865 15419
rect 20023 15393 20141 15419
rect 5027 15257 5145 15283
rect 5107 15255 5145 15257
rect 5487 15257 6433 15283
rect 6591 15257 7537 15283
rect 7695 15257 8641 15283
rect 8799 15257 9745 15283
rect 10087 15257 10481 15283
rect 10639 15257 11585 15283
rect 11743 15257 12689 15283
rect 5107 15239 5173 15255
rect 4999 15199 5065 15215
rect 4999 15165 5015 15199
rect 5049 15165 5065 15199
rect 5107 15205 5123 15239
rect 5157 15205 5173 15239
rect 5107 15189 5173 15205
rect 5487 15235 5941 15257
rect 5487 15201 5763 15235
rect 5797 15201 5941 15235
rect 6591 15235 7045 15257
rect 5487 15185 5941 15201
rect 5983 15199 6433 15215
rect 4999 15149 5065 15165
rect 5027 15147 5065 15149
rect 5983 15165 6127 15199
rect 6161 15165 6433 15199
rect 6591 15201 6867 15235
rect 6901 15201 7045 15235
rect 7695 15235 8149 15257
rect 6591 15185 7045 15201
rect 7087 15199 7537 15215
rect 5027 15117 5145 15147
rect 5983 15143 6433 15165
rect 7087 15165 7231 15199
rect 7265 15165 7537 15199
rect 7695 15201 7971 15235
rect 8005 15201 8149 15235
rect 8799 15235 9253 15257
rect 7695 15185 8149 15201
rect 8191 15199 8641 15215
rect 7087 15143 7537 15165
rect 8191 15165 8335 15199
rect 8369 15165 8641 15199
rect 8799 15201 9075 15235
rect 9109 15201 9253 15235
rect 10087 15235 10263 15257
rect 8799 15185 9253 15201
rect 9295 15199 9745 15215
rect 8191 15143 8641 15165
rect 9295 15165 9439 15199
rect 9473 15165 9745 15199
rect 10087 15201 10103 15235
rect 10137 15201 10213 15235
rect 10247 15201 10263 15235
rect 10639 15235 11093 15257
rect 10087 15185 10263 15201
rect 10305 15199 10481 15215
rect 9295 15143 9745 15165
rect 10305 15165 10321 15199
rect 10355 15165 10431 15199
rect 10465 15165 10481 15199
rect 10639 15201 10915 15235
rect 10949 15201 11093 15235
rect 11743 15235 12197 15257
rect 12869 15241 12899 15309
rect 10639 15185 11093 15201
rect 11135 15199 11585 15215
rect 10305 15143 10481 15165
rect 11135 15165 11279 15199
rect 11313 15165 11585 15199
rect 11743 15201 12019 15235
rect 12053 15201 12197 15235
rect 12839 15225 12899 15241
rect 11743 15185 12197 15201
rect 12239 15199 12689 15215
rect 11135 15143 11585 15165
rect 12239 15165 12383 15199
rect 12417 15165 12689 15199
rect 12839 15191 12849 15225
rect 12883 15191 12899 15225
rect 12839 15175 12899 15191
rect 12239 15143 12689 15165
rect 5487 15117 6433 15143
rect 6591 15117 7537 15143
rect 7695 15117 8641 15143
rect 8799 15117 9745 15143
rect 10087 15117 10481 15143
rect 10639 15117 11585 15143
rect 11743 15117 12689 15143
rect 12869 15027 12899 15175
rect 12953 15225 13053 15309
rect 13211 15241 13311 15309
rect 13376 15241 13406 15263
rect 13583 15257 13793 15283
rect 13951 15257 14897 15283
rect 15147 15257 15265 15283
rect 13583 15251 13667 15257
rect 12953 15191 12963 15225
rect 12997 15191 13053 15225
rect 12953 15027 13053 15191
rect 13157 15225 13311 15241
rect 13157 15191 13167 15225
rect 13201 15191 13311 15225
rect 13157 15175 13311 15191
rect 13353 15225 13407 15241
rect 13353 15191 13363 15225
rect 13397 15191 13407 15225
rect 13353 15175 13407 15191
rect 13525 15235 13667 15251
rect 13525 15201 13541 15235
rect 13575 15201 13667 15235
rect 13951 15235 14405 15257
rect 15147 15255 15185 15257
rect 13525 15185 13667 15201
rect 13709 15199 13851 15215
rect 13211 15027 13311 15175
rect 13376 15143 13406 15175
rect 13709 15165 13801 15199
rect 13835 15165 13851 15199
rect 13951 15201 14227 15235
rect 14261 15201 14405 15235
rect 15119 15239 15185 15255
rect 15445 15241 15475 15309
rect 13951 15185 14405 15201
rect 14447 15199 14897 15215
rect 13709 15149 13851 15165
rect 14447 15165 14591 15199
rect 14625 15165 14897 15199
rect 15119 15205 15135 15239
rect 15169 15205 15185 15239
rect 15415 15225 15475 15241
rect 15119 15189 15185 15205
rect 15227 15199 15293 15215
rect 13709 15143 13793 15149
rect 14447 15143 14897 15165
rect 15227 15165 15243 15199
rect 15277 15165 15293 15199
rect 15415 15191 15425 15225
rect 15459 15191 15475 15225
rect 15415 15175 15475 15191
rect 15227 15149 15293 15165
rect 15227 15147 15265 15149
rect 13583 15117 13793 15143
rect 13951 15117 14897 15143
rect 15147 15117 15265 15147
rect 15445 15027 15475 15175
rect 15529 15225 15629 15309
rect 15787 15241 15887 15309
rect 15952 15241 15982 15263
rect 16159 15257 16553 15283
rect 16711 15257 17657 15283
rect 17815 15257 18761 15283
rect 18919 15257 19865 15283
rect 20023 15257 20141 15283
rect 15529 15191 15539 15225
rect 15573 15191 15629 15225
rect 15529 15027 15629 15191
rect 15733 15225 15887 15241
rect 15733 15191 15743 15225
rect 15777 15191 15887 15225
rect 15733 15175 15887 15191
rect 15929 15225 15983 15241
rect 15929 15191 15939 15225
rect 15973 15191 15983 15225
rect 15929 15175 15983 15191
rect 16159 15235 16335 15257
rect 16159 15201 16175 15235
rect 16209 15201 16285 15235
rect 16319 15201 16335 15235
rect 16711 15235 17165 15257
rect 16159 15185 16335 15201
rect 16377 15199 16553 15215
rect 15787 15027 15887 15175
rect 15952 15143 15982 15175
rect 16377 15165 16393 15199
rect 16427 15165 16503 15199
rect 16537 15165 16553 15199
rect 16711 15201 16987 15235
rect 17021 15201 17165 15235
rect 17815 15235 18269 15257
rect 16711 15185 17165 15201
rect 17207 15199 17657 15215
rect 16377 15143 16553 15165
rect 17207 15165 17351 15199
rect 17385 15165 17657 15199
rect 17815 15201 18091 15235
rect 18125 15201 18269 15235
rect 18919 15235 19373 15257
rect 20023 15255 20061 15257
rect 17815 15185 18269 15201
rect 18311 15199 18761 15215
rect 17207 15143 17657 15165
rect 18311 15165 18455 15199
rect 18489 15165 18761 15199
rect 18919 15201 19195 15235
rect 19229 15201 19373 15235
rect 19995 15239 20061 15255
rect 18919 15185 19373 15201
rect 19415 15199 19865 15215
rect 18311 15143 18761 15165
rect 19415 15165 19559 15199
rect 19593 15165 19865 15199
rect 19995 15205 20011 15239
rect 20045 15205 20061 15239
rect 19995 15189 20061 15205
rect 20103 15199 20169 15215
rect 19415 15143 19865 15165
rect 20103 15165 20119 15199
rect 20153 15165 20169 15199
rect 20103 15149 20169 15165
rect 20103 15147 20141 15149
rect 16159 15117 16553 15143
rect 16711 15117 17657 15143
rect 17815 15117 18761 15143
rect 18919 15117 19865 15143
rect 20023 15117 20141 15147
rect 5027 14917 5145 14943
rect 5487 14917 6433 14943
rect 6591 14917 7537 14943
rect 7695 14917 8641 14943
rect 8799 14917 9745 14943
rect 10087 14917 10481 14943
rect 10639 14917 11585 14943
rect 11743 14917 12689 14943
rect 12869 14917 12899 14943
rect 12953 14917 13053 14943
rect 13211 14917 13311 14943
rect 13376 14917 13406 14943
rect 13583 14917 13793 14943
rect 13951 14917 14897 14943
rect 15147 14917 15265 14943
rect 15445 14917 15475 14943
rect 15529 14917 15629 14943
rect 15787 14917 15887 14943
rect 15952 14917 15982 14943
rect 16159 14917 16553 14943
rect 16711 14917 17657 14943
rect 17815 14917 18761 14943
rect 18919 14917 19865 14943
rect 20023 14917 20141 14943
rect 5027 14849 5145 14875
rect 5487 14849 6065 14875
rect 6223 14849 7169 14875
rect 7419 14849 8365 14875
rect 8523 14849 9469 14875
rect 9627 14849 10573 14875
rect 11371 14849 11401 14875
rect 11743 14849 12321 14875
rect 13395 14849 13425 14875
rect 13583 14849 14161 14875
rect 14319 14849 14349 14875
rect 14407 14849 14437 14875
rect 14595 14849 14625 14875
rect 14810 14849 14840 14875
rect 14894 14849 14924 14875
rect 15002 14849 15032 14875
rect 15086 14849 15116 14875
rect 15172 14849 15202 14875
rect 15271 14849 15301 14875
rect 15468 14849 15498 14875
rect 15565 14849 15595 14875
rect 15705 14849 15735 14875
rect 15804 14849 15834 14875
rect 15896 14849 15926 14875
rect 5027 14645 5145 14675
rect 5487 14649 6065 14675
rect 6223 14649 7169 14675
rect 10777 14810 10807 14836
rect 10873 14810 10903 14836
rect 10945 14810 10975 14836
rect 11159 14810 11189 14836
rect 11262 14810 11292 14836
rect 10777 14694 10807 14726
rect 10777 14678 10831 14694
rect 7419 14649 8365 14675
rect 8523 14649 9469 14675
rect 9627 14649 10573 14675
rect 5027 14643 5065 14645
rect 4999 14627 5065 14643
rect 4999 14593 5015 14627
rect 5049 14593 5065 14627
rect 5801 14627 6065 14649
rect 4999 14577 5065 14593
rect 5107 14587 5173 14603
rect 5107 14553 5123 14587
rect 5157 14553 5173 14587
rect 5107 14537 5173 14553
rect 5487 14591 5759 14607
rect 5487 14557 5503 14591
rect 5537 14557 5606 14591
rect 5640 14557 5709 14591
rect 5743 14557 5759 14591
rect 5801 14593 5817 14627
rect 5851 14593 5916 14627
rect 5950 14593 6015 14627
rect 6049 14593 6065 14627
rect 6719 14627 7169 14649
rect 5801 14577 6065 14593
rect 6223 14591 6677 14607
rect 5107 14535 5145 14537
rect 5027 14509 5145 14535
rect 5487 14535 5759 14557
rect 6223 14557 6499 14591
rect 6533 14557 6677 14591
rect 6719 14593 6863 14627
rect 6897 14593 7169 14627
rect 7915 14627 8365 14649
rect 6719 14577 7169 14593
rect 7419 14591 7873 14607
rect 6223 14535 6677 14557
rect 7419 14557 7695 14591
rect 7729 14557 7873 14591
rect 7915 14593 8059 14627
rect 8093 14593 8365 14627
rect 9019 14627 9469 14649
rect 7915 14577 8365 14593
rect 8523 14591 8977 14607
rect 7419 14535 7873 14557
rect 8523 14557 8799 14591
rect 8833 14557 8977 14591
rect 9019 14593 9163 14627
rect 9197 14593 9469 14627
rect 10123 14627 10573 14649
rect 9019 14577 9469 14593
rect 9627 14591 10081 14607
rect 8523 14535 8977 14557
rect 9627 14557 9903 14591
rect 9937 14557 10081 14591
rect 10123 14593 10267 14627
rect 10301 14593 10573 14627
rect 10123 14577 10573 14593
rect 10777 14644 10787 14678
rect 10821 14644 10831 14678
rect 10777 14628 10831 14644
rect 9627 14535 10081 14557
rect 5487 14509 6065 14535
rect 6223 14509 7169 14535
rect 7419 14509 8365 14535
rect 8523 14509 9469 14535
rect 9627 14509 10573 14535
rect 10777 14483 10807 14628
rect 10873 14575 10903 14726
rect 10945 14694 10975 14726
rect 11159 14711 11189 14726
rect 10945 14678 10999 14694
rect 10945 14644 10955 14678
rect 10989 14644 10999 14678
rect 10945 14628 10999 14644
rect 11041 14681 11189 14711
rect 11041 14581 11071 14681
rect 11262 14617 11292 14726
rect 12801 14810 12831 14836
rect 12897 14810 12927 14836
rect 12969 14810 12999 14836
rect 13183 14810 13213 14836
rect 13286 14810 13316 14836
rect 11743 14649 12321 14675
rect 12801 14694 12831 14726
rect 12801 14678 12855 14694
rect 11371 14617 11401 14649
rect 12057 14627 12321 14649
rect 11254 14601 11308 14617
rect 10849 14565 10915 14575
rect 10849 14531 10865 14565
rect 10899 14551 10915 14565
rect 11017 14565 11071 14581
rect 10899 14531 10975 14551
rect 10849 14521 10975 14531
rect 10945 14483 10975 14521
rect 11017 14531 11027 14565
rect 11061 14531 11071 14565
rect 11017 14515 11071 14531
rect 11113 14565 11196 14581
rect 11113 14531 11123 14565
rect 11157 14531 11196 14565
rect 11254 14567 11264 14601
rect 11298 14567 11308 14601
rect 11254 14551 11308 14567
rect 11350 14601 11404 14617
rect 11350 14567 11360 14601
rect 11394 14567 11404 14601
rect 11350 14551 11404 14567
rect 11743 14591 12015 14607
rect 11743 14557 11759 14591
rect 11793 14557 11862 14591
rect 11896 14557 11965 14591
rect 11999 14557 12015 14591
rect 12057 14593 12073 14627
rect 12107 14593 12172 14627
rect 12206 14593 12271 14627
rect 12305 14593 12321 14627
rect 12057 14577 12321 14593
rect 12801 14644 12811 14678
rect 12845 14644 12855 14678
rect 12801 14628 12855 14644
rect 11113 14515 11196 14531
rect 11041 14483 11071 14515
rect 11166 14483 11196 14515
rect 11262 14483 11292 14551
rect 11371 14529 11401 14551
rect 11743 14535 12015 14557
rect 11743 14509 12321 14535
rect 12801 14483 12831 14628
rect 12897 14575 12927 14726
rect 12969 14694 12999 14726
rect 13183 14711 13213 14726
rect 12969 14678 13023 14694
rect 12969 14644 12979 14678
rect 13013 14644 13023 14678
rect 12969 14628 13023 14644
rect 13065 14681 13213 14711
rect 13065 14581 13095 14681
rect 13286 14617 13316 14726
rect 14319 14676 14349 14691
rect 13583 14649 14161 14675
rect 13395 14617 13425 14649
rect 13897 14627 14161 14649
rect 13278 14601 13332 14617
rect 12873 14565 12939 14575
rect 12873 14531 12889 14565
rect 12923 14551 12939 14565
rect 13041 14565 13095 14581
rect 12923 14531 12999 14551
rect 12873 14521 12999 14531
rect 12969 14483 12999 14521
rect 13041 14531 13051 14565
rect 13085 14531 13095 14565
rect 13041 14515 13095 14531
rect 13137 14565 13220 14581
rect 13137 14531 13147 14565
rect 13181 14531 13220 14565
rect 13278 14567 13288 14601
rect 13322 14567 13332 14601
rect 13278 14551 13332 14567
rect 13374 14601 13428 14617
rect 13374 14567 13384 14601
rect 13418 14567 13428 14601
rect 13374 14551 13428 14567
rect 13583 14591 13855 14607
rect 13583 14557 13599 14591
rect 13633 14557 13702 14591
rect 13736 14557 13805 14591
rect 13839 14557 13855 14591
rect 13897 14593 13913 14627
rect 13947 14593 14012 14627
rect 14046 14593 14111 14627
rect 14145 14593 14161 14627
rect 14313 14652 14349 14676
rect 14313 14617 14343 14652
rect 14407 14630 14437 14691
rect 14810 14717 14840 14765
rect 14798 14701 14852 14717
rect 14798 14667 14808 14701
rect 14842 14667 14852 14701
rect 14798 14651 14852 14667
rect 13897 14577 14161 14593
rect 14267 14601 14343 14617
rect 13137 14515 13220 14531
rect 13065 14483 13095 14515
rect 13190 14483 13220 14515
rect 13286 14483 13316 14551
rect 13395 14529 13425 14551
rect 13583 14535 13855 14557
rect 14267 14567 14277 14601
rect 14311 14567 14343 14601
rect 14267 14551 14343 14567
rect 14387 14614 14441 14630
rect 14387 14580 14397 14614
rect 14431 14580 14441 14614
rect 14387 14564 14441 14580
rect 14595 14617 14625 14649
rect 14595 14601 14654 14617
rect 14595 14567 14610 14601
rect 14644 14567 14654 14601
rect 14313 14542 14343 14551
rect 13583 14509 14161 14535
rect 14313 14518 14349 14542
rect 14319 14503 14349 14518
rect 14407 14503 14437 14564
rect 14595 14551 14654 14567
rect 14595 14529 14625 14551
rect 14803 14483 14833 14651
rect 14894 14609 14924 14765
rect 14875 14593 14929 14609
rect 14875 14559 14885 14593
rect 14919 14559 14929 14593
rect 15002 14581 15032 14765
rect 15086 14733 15116 14765
rect 15076 14717 15130 14733
rect 15076 14683 15086 14717
rect 15120 14683 15130 14717
rect 15076 14667 15130 14683
rect 15172 14631 15202 14765
rect 16163 14843 16193 14869
rect 16247 14843 16277 14869
rect 16527 14849 17473 14875
rect 17815 14849 18761 14875
rect 18919 14849 19865 14875
rect 20023 14849 20141 14875
rect 15271 14666 15301 14681
rect 15271 14636 15377 14666
rect 15152 14619 15202 14631
rect 15139 14607 15202 14619
rect 14875 14543 14929 14559
rect 14971 14565 15032 14581
rect 14894 14483 14924 14543
rect 14971 14531 14981 14565
rect 15015 14545 15032 14565
rect 15115 14601 15202 14607
rect 15347 14619 15377 14636
rect 15347 14603 15413 14619
rect 15115 14591 15181 14601
rect 15115 14557 15125 14591
rect 15159 14589 15181 14591
rect 15159 14557 15169 14589
rect 15347 14569 15369 14603
rect 15403 14569 15413 14603
rect 15468 14571 15498 14765
rect 15565 14707 15595 14765
rect 15540 14691 15595 14707
rect 15540 14657 15551 14691
rect 15585 14657 15595 14691
rect 15540 14641 15595 14657
rect 15015 14531 15073 14545
rect 15115 14541 15169 14557
rect 14971 14515 15073 14531
rect 15043 14483 15073 14515
rect 15139 14471 15169 14541
rect 15211 14543 15278 14559
rect 15211 14509 15221 14543
rect 15255 14509 15278 14543
rect 15347 14553 15413 14569
rect 15455 14555 15509 14571
rect 15347 14527 15377 14553
rect 15211 14493 15278 14509
rect 15248 14471 15278 14493
rect 15455 14521 15465 14555
rect 15499 14521 15509 14555
rect 15455 14505 15509 14521
rect 15479 14483 15509 14505
rect 15551 14483 15581 14641
rect 15705 14631 15735 14765
rect 15804 14727 15834 14765
rect 15784 14717 15850 14727
rect 15784 14683 15800 14717
rect 15834 14683 15850 14717
rect 15784 14673 15850 14683
rect 15896 14678 15926 14765
rect 15896 14662 16025 14678
rect 15896 14648 15981 14662
rect 15705 14601 15843 14631
rect 15812 14571 15843 14601
rect 15908 14628 15981 14648
rect 16015 14628 16025 14662
rect 15908 14612 16025 14628
rect 16163 14626 16193 14715
rect 16247 14700 16277 14715
rect 16247 14670 16310 14700
rect 16163 14616 16238 14626
rect 15704 14549 15770 14559
rect 15704 14515 15720 14549
rect 15754 14515 15770 14549
rect 15704 14505 15770 14515
rect 15812 14555 15866 14571
rect 15812 14521 15822 14555
rect 15856 14521 15866 14555
rect 15812 14505 15866 14521
rect 15717 14471 15747 14505
rect 15813 14471 15843 14505
rect 15908 14483 15938 14612
rect 16163 14582 16188 14616
rect 16222 14582 16238 14616
rect 16163 14572 16238 14582
rect 16280 14617 16310 14670
rect 16527 14649 17473 14675
rect 17815 14649 18761 14675
rect 18919 14649 19865 14675
rect 17023 14627 17473 14649
rect 16280 14601 16334 14617
rect 16163 14483 16193 14572
rect 16280 14567 16290 14601
rect 16324 14567 16334 14601
rect 16280 14551 16334 14567
rect 16527 14591 16981 14607
rect 16527 14557 16803 14591
rect 16837 14557 16981 14591
rect 17023 14593 17167 14627
rect 17201 14593 17473 14627
rect 18311 14627 18761 14649
rect 17023 14577 17473 14593
rect 17815 14591 18269 14607
rect 16280 14528 16310 14551
rect 16247 14498 16310 14528
rect 16527 14535 16981 14557
rect 17815 14557 18091 14591
rect 18125 14557 18269 14591
rect 18311 14593 18455 14627
rect 18489 14593 18761 14627
rect 19415 14627 19865 14649
rect 20023 14645 20141 14675
rect 18311 14577 18761 14593
rect 18919 14591 19373 14607
rect 17815 14535 18269 14557
rect 18919 14557 19195 14591
rect 19229 14557 19373 14591
rect 19415 14593 19559 14627
rect 19593 14593 19865 14627
rect 20103 14643 20141 14645
rect 20103 14627 20169 14643
rect 19415 14577 19865 14593
rect 19995 14587 20061 14603
rect 18919 14535 19373 14557
rect 19995 14553 20011 14587
rect 20045 14553 20061 14587
rect 20103 14593 20119 14627
rect 20153 14593 20169 14627
rect 20103 14577 20169 14593
rect 19995 14537 20061 14553
rect 20023 14535 20061 14537
rect 16527 14509 17473 14535
rect 16247 14483 16277 14498
rect 17815 14509 18761 14535
rect 18919 14509 19865 14535
rect 20023 14509 20141 14535
rect 5027 14373 5145 14399
rect 5487 14373 6065 14399
rect 6223 14373 7169 14399
rect 7419 14373 8365 14399
rect 8523 14373 9469 14399
rect 9627 14373 10573 14399
rect 10777 14373 10807 14399
rect 10945 14373 10975 14399
rect 11041 14373 11071 14399
rect 11166 14373 11196 14399
rect 11262 14373 11292 14399
rect 11371 14373 11401 14399
rect 11743 14373 12321 14399
rect 12801 14373 12831 14399
rect 12969 14373 12999 14399
rect 13065 14373 13095 14399
rect 13190 14373 13220 14399
rect 13286 14373 13316 14399
rect 13395 14373 13425 14399
rect 13583 14373 14161 14399
rect 14319 14373 14349 14399
rect 14407 14373 14437 14399
rect 14595 14373 14625 14399
rect 14803 14373 14833 14399
rect 14894 14373 14924 14399
rect 15043 14373 15073 14399
rect 15139 14373 15169 14399
rect 15248 14373 15278 14399
rect 15347 14373 15377 14399
rect 15479 14373 15509 14399
rect 15551 14373 15581 14399
rect 15717 14373 15747 14399
rect 15813 14373 15843 14399
rect 15908 14373 15938 14399
rect 16163 14373 16193 14399
rect 16247 14373 16277 14399
rect 16527 14373 17473 14399
rect 17815 14373 18761 14399
rect 18919 14373 19865 14399
rect 20023 14373 20141 14399
rect 5027 14305 5145 14331
rect 5487 14305 6433 14331
rect 6591 14305 7537 14331
rect 7695 14305 8641 14331
rect 8799 14305 9745 14331
rect 10179 14305 10209 14331
rect 10387 14305 10417 14331
rect 10478 14305 10508 14331
rect 10627 14305 10657 14331
rect 10723 14305 10753 14331
rect 10832 14305 10862 14331
rect 10931 14305 10961 14331
rect 11063 14305 11093 14331
rect 11135 14305 11165 14331
rect 11301 14305 11331 14331
rect 11397 14305 11427 14331
rect 11492 14305 11522 14331
rect 11747 14305 11777 14331
rect 11831 14305 11861 14331
rect 12019 14305 12049 14331
rect 12107 14305 12137 14331
rect 12313 14305 12343 14331
rect 12399 14305 12429 14331
rect 12485 14305 12515 14331
rect 12571 14305 12601 14331
rect 12657 14305 12687 14331
rect 12743 14305 12773 14331
rect 12829 14305 12859 14331
rect 12915 14305 12945 14331
rect 13000 14305 13030 14331
rect 13086 14305 13116 14331
rect 13172 14305 13202 14331
rect 13258 14305 13288 14331
rect 13344 14305 13374 14331
rect 13430 14305 13460 14331
rect 13516 14305 13546 14331
rect 13602 14305 13632 14331
rect 13688 14305 13718 14331
rect 13774 14305 13804 14331
rect 13860 14305 13890 14331
rect 13946 14305 13976 14331
rect 14341 14305 14371 14331
rect 14425 14305 14525 14331
rect 14683 14305 14783 14331
rect 14848 14305 14878 14331
rect 15239 14305 15269 14331
rect 15348 14305 15378 14331
rect 15444 14305 15474 14331
rect 15569 14305 15599 14331
rect 15665 14305 15695 14331
rect 15833 14305 15863 14331
rect 16067 14305 16097 14331
rect 16155 14305 16185 14331
rect 16343 14305 16373 14331
rect 16431 14305 16461 14331
rect 16711 14305 17657 14331
rect 17815 14305 18761 14331
rect 18919 14305 19865 14331
rect 20023 14305 20141 14331
rect 5027 14169 5145 14195
rect 5107 14167 5145 14169
rect 5487 14169 6433 14195
rect 6591 14169 7537 14195
rect 7695 14169 8641 14195
rect 8799 14169 9745 14195
rect 5107 14151 5173 14167
rect 4999 14111 5065 14127
rect 4999 14077 5015 14111
rect 5049 14077 5065 14111
rect 5107 14117 5123 14151
rect 5157 14117 5173 14151
rect 5107 14101 5173 14117
rect 5487 14147 5941 14169
rect 5487 14113 5763 14147
rect 5797 14113 5941 14147
rect 6591 14147 7045 14169
rect 5487 14097 5941 14113
rect 5983 14111 6433 14127
rect 4999 14061 5065 14077
rect 5027 14059 5065 14061
rect 5983 14077 6127 14111
rect 6161 14077 6433 14111
rect 6591 14113 6867 14147
rect 6901 14113 7045 14147
rect 7695 14147 8149 14169
rect 6591 14097 7045 14113
rect 7087 14111 7537 14127
rect 5027 14029 5145 14059
rect 5983 14055 6433 14077
rect 7087 14077 7231 14111
rect 7265 14077 7537 14111
rect 7695 14113 7971 14147
rect 8005 14113 8149 14147
rect 8799 14147 9253 14169
rect 7695 14097 8149 14113
rect 8191 14111 8641 14127
rect 7087 14055 7537 14077
rect 8191 14077 8335 14111
rect 8369 14077 8641 14111
rect 8799 14113 9075 14147
rect 9109 14113 9253 14147
rect 10179 14153 10209 14175
rect 10179 14137 10238 14153
rect 8799 14097 9253 14113
rect 9295 14111 9745 14127
rect 8191 14055 8641 14077
rect 9295 14077 9439 14111
rect 9473 14077 9745 14111
rect 9295 14055 9745 14077
rect 10179 14103 10194 14137
rect 10228 14103 10238 14137
rect 10179 14087 10238 14103
rect 10179 14055 10209 14087
rect 5487 14029 6433 14055
rect 6591 14029 7537 14055
rect 7695 14029 8641 14055
rect 8799 14029 9745 14055
rect 10387 14053 10417 14221
rect 10478 14161 10508 14221
rect 10627 14189 10657 14221
rect 10555 14173 10657 14189
rect 10459 14145 10513 14161
rect 10459 14111 10469 14145
rect 10503 14111 10513 14145
rect 10555 14139 10565 14173
rect 10599 14159 10657 14173
rect 10723 14163 10753 14233
rect 10832 14211 10862 14233
rect 10599 14139 10616 14159
rect 10555 14123 10616 14139
rect 10459 14095 10513 14111
rect 10382 14037 10436 14053
rect 10382 14003 10392 14037
rect 10426 14003 10436 14037
rect 10382 13987 10436 14003
rect 10394 13939 10424 13987
rect 10478 13939 10508 14095
rect 10586 13939 10616 14123
rect 10699 14147 10753 14163
rect 10699 14113 10709 14147
rect 10743 14115 10753 14147
rect 10795 14195 10862 14211
rect 10795 14161 10805 14195
rect 10839 14161 10862 14195
rect 11063 14199 11093 14221
rect 11039 14183 11093 14199
rect 10795 14145 10862 14161
rect 10931 14151 10961 14177
rect 10931 14135 10997 14151
rect 10743 14113 10765 14115
rect 10699 14103 10765 14113
rect 10699 14097 10786 14103
rect 10723 14085 10786 14097
rect 10736 14073 10786 14085
rect 10660 14021 10714 14037
rect 10660 13987 10670 14021
rect 10704 13987 10714 14021
rect 10660 13971 10714 13987
rect 10670 13939 10700 13971
rect 10756 13939 10786 14073
rect 10931 14101 10953 14135
rect 10987 14101 10997 14135
rect 11039 14149 11049 14183
rect 11083 14149 11093 14183
rect 11039 14133 11093 14149
rect 10931 14085 10997 14101
rect 10931 14068 10961 14085
rect 10855 14038 10961 14068
rect 10855 14023 10885 14038
rect 11052 13939 11082 14133
rect 11135 14063 11165 14221
rect 11301 14199 11331 14233
rect 11397 14199 11427 14233
rect 11288 14189 11354 14199
rect 11288 14155 11304 14189
rect 11338 14155 11354 14189
rect 11288 14145 11354 14155
rect 11396 14183 11450 14199
rect 11396 14149 11406 14183
rect 11440 14149 11450 14183
rect 11396 14133 11450 14149
rect 11396 14103 11427 14133
rect 11289 14073 11427 14103
rect 11492 14092 11522 14221
rect 11747 14132 11777 14221
rect 11831 14206 11861 14221
rect 11831 14176 11894 14206
rect 11864 14153 11894 14176
rect 11864 14137 11918 14153
rect 12019 14140 12049 14201
rect 12107 14186 12137 14201
rect 12107 14162 12143 14186
rect 12113 14153 12143 14162
rect 12313 14162 12343 14221
rect 12399 14162 12429 14221
rect 12485 14162 12515 14221
rect 12571 14162 12601 14221
rect 12657 14162 12687 14221
rect 12743 14162 12773 14221
rect 12829 14162 12859 14221
rect 12915 14162 12945 14221
rect 13000 14162 13030 14221
rect 13086 14162 13116 14221
rect 13172 14162 13202 14221
rect 13258 14162 13288 14221
rect 13344 14162 13374 14221
rect 13430 14162 13460 14221
rect 13516 14162 13546 14221
rect 13602 14162 13632 14221
rect 11747 14122 11822 14132
rect 11492 14076 11609 14092
rect 11124 14047 11179 14063
rect 11124 14013 11135 14047
rect 11169 14013 11179 14047
rect 11124 13997 11179 14013
rect 11149 13939 11179 13997
rect 11289 13939 11319 14073
rect 11492 14056 11565 14076
rect 11480 14042 11565 14056
rect 11599 14042 11609 14076
rect 11368 14021 11434 14031
rect 11368 13987 11384 14021
rect 11418 13987 11434 14021
rect 11368 13977 11434 13987
rect 11480 14026 11609 14042
rect 11747 14088 11772 14122
rect 11806 14088 11822 14122
rect 11747 14078 11822 14088
rect 11864 14103 11874 14137
rect 11908 14103 11918 14137
rect 11864 14087 11918 14103
rect 12015 14124 12069 14140
rect 12015 14090 12025 14124
rect 12059 14090 12069 14124
rect 11388 13939 11418 13977
rect 11480 13939 11510 14026
rect 11747 13989 11777 14078
rect 11864 14034 11894 14087
rect 12015 14074 12069 14090
rect 12113 14137 12189 14153
rect 12113 14103 12145 14137
rect 12179 14103 12189 14137
rect 12113 14087 12189 14103
rect 12313 14137 13632 14162
rect 12313 14103 12538 14137
rect 12572 14103 12606 14137
rect 12640 14103 12674 14137
rect 12708 14103 12742 14137
rect 12776 14103 12810 14137
rect 12844 14103 12878 14137
rect 12912 14103 12946 14137
rect 12980 14103 13014 14137
rect 13048 14103 13082 14137
rect 13116 14103 13150 14137
rect 13184 14103 13218 14137
rect 13252 14103 13286 14137
rect 13320 14103 13354 14137
rect 13388 14103 13422 14137
rect 13456 14103 13490 14137
rect 13524 14103 13558 14137
rect 13592 14103 13632 14137
rect 12313 14087 13632 14103
rect 11831 14004 11894 14034
rect 12019 14013 12049 14074
rect 12113 14052 12143 14087
rect 12313 14055 12343 14087
rect 12399 14055 12429 14087
rect 12485 14055 12515 14087
rect 12571 14055 12601 14087
rect 12657 14055 12687 14087
rect 12743 14055 12773 14087
rect 12829 14055 12859 14087
rect 12915 14055 12945 14087
rect 13000 14055 13030 14087
rect 13086 14055 13116 14087
rect 13172 14055 13202 14087
rect 13258 14055 13288 14087
rect 13344 14055 13374 14087
rect 13430 14055 13460 14087
rect 13516 14055 13546 14087
rect 13602 14055 13632 14087
rect 13688 14172 13718 14221
rect 13774 14172 13804 14221
rect 13860 14172 13890 14221
rect 13946 14172 13976 14221
rect 13688 14137 14035 14172
rect 14341 14153 14371 14221
rect 13688 14103 13985 14137
rect 14019 14103 14035 14137
rect 13688 14070 14035 14103
rect 14311 14137 14371 14153
rect 14311 14103 14321 14137
rect 14355 14103 14371 14137
rect 14311 14087 14371 14103
rect 13688 14055 13718 14070
rect 13774 14055 13804 14070
rect 13860 14055 13890 14070
rect 13946 14055 13976 14070
rect 12107 14028 12143 14052
rect 12107 14013 12137 14028
rect 11831 13989 11861 14004
rect 5027 13829 5145 13855
rect 5487 13829 6433 13855
rect 6591 13829 7537 13855
rect 7695 13829 8641 13855
rect 8799 13829 9745 13855
rect 10179 13829 10209 13855
rect 10394 13829 10424 13855
rect 10478 13829 10508 13855
rect 10586 13829 10616 13855
rect 10670 13829 10700 13855
rect 10756 13829 10786 13855
rect 10855 13829 10885 13855
rect 11052 13829 11082 13855
rect 11149 13829 11179 13855
rect 11289 13829 11319 13855
rect 11388 13829 11418 13855
rect 11480 13829 11510 13855
rect 11747 13835 11777 13861
rect 11831 13835 11861 13861
rect 14341 13939 14371 14087
rect 14425 14137 14525 14221
rect 14683 14153 14783 14221
rect 14848 14153 14878 14175
rect 15239 14153 15269 14175
rect 15348 14153 15378 14221
rect 15444 14189 15474 14221
rect 15569 14189 15599 14221
rect 15444 14173 15527 14189
rect 14425 14103 14435 14137
rect 14469 14103 14525 14137
rect 14425 13939 14525 14103
rect 14629 14137 14783 14153
rect 14629 14103 14639 14137
rect 14673 14103 14783 14137
rect 14629 14087 14783 14103
rect 14825 14137 14879 14153
rect 14825 14103 14835 14137
rect 14869 14103 14879 14137
rect 14825 14087 14879 14103
rect 15236 14137 15290 14153
rect 15236 14103 15246 14137
rect 15280 14103 15290 14137
rect 15236 14087 15290 14103
rect 15332 14137 15386 14153
rect 15332 14103 15342 14137
rect 15376 14103 15386 14137
rect 15444 14139 15483 14173
rect 15517 14139 15527 14173
rect 15444 14123 15527 14139
rect 15569 14173 15623 14189
rect 15569 14139 15579 14173
rect 15613 14139 15623 14173
rect 15665 14183 15695 14221
rect 15665 14173 15791 14183
rect 15665 14153 15741 14173
rect 15569 14123 15623 14139
rect 15725 14139 15741 14153
rect 15775 14139 15791 14173
rect 15725 14129 15791 14139
rect 15332 14087 15386 14103
rect 14683 13939 14783 14087
rect 14848 14055 14878 14087
rect 15239 14055 15269 14087
rect 15348 13978 15378 14087
rect 15569 14023 15599 14123
rect 15451 13993 15599 14023
rect 15641 14060 15695 14076
rect 15641 14026 15651 14060
rect 15685 14026 15695 14060
rect 15641 14010 15695 14026
rect 15451 13978 15481 13993
rect 15665 13978 15695 14010
rect 15737 13978 15767 14129
rect 15833 14076 15863 14221
rect 16067 14140 16097 14201
rect 16155 14186 16185 14201
rect 16155 14162 16191 14186
rect 16161 14153 16191 14162
rect 15809 14060 15863 14076
rect 16063 14124 16117 14140
rect 16063 14090 16073 14124
rect 16107 14090 16117 14124
rect 16063 14074 16117 14090
rect 16161 14137 16237 14153
rect 16343 14140 16373 14201
rect 16431 14186 16461 14201
rect 16431 14162 16467 14186
rect 16437 14153 16467 14162
rect 16711 14169 17657 14195
rect 17815 14169 18761 14195
rect 18919 14169 19865 14195
rect 20023 14169 20141 14195
rect 16161 14103 16193 14137
rect 16227 14103 16237 14137
rect 16161 14087 16237 14103
rect 16339 14124 16393 14140
rect 16339 14090 16349 14124
rect 16383 14090 16393 14124
rect 15809 14026 15819 14060
rect 15853 14026 15863 14060
rect 15809 14010 15863 14026
rect 16067 14013 16097 14074
rect 16161 14052 16191 14087
rect 16339 14074 16393 14090
rect 16437 14137 16513 14153
rect 16437 14103 16469 14137
rect 16503 14103 16513 14137
rect 16437 14087 16513 14103
rect 16711 14147 17165 14169
rect 16711 14113 16987 14147
rect 17021 14113 17165 14147
rect 17815 14147 18269 14169
rect 16711 14097 17165 14113
rect 17207 14111 17657 14127
rect 16155 14028 16191 14052
rect 16155 14013 16185 14028
rect 16343 14013 16373 14074
rect 16437 14052 16467 14087
rect 17207 14077 17351 14111
rect 17385 14077 17657 14111
rect 17815 14113 18091 14147
rect 18125 14113 18269 14147
rect 18919 14147 19373 14169
rect 20023 14167 20061 14169
rect 17815 14097 18269 14113
rect 18311 14111 18761 14127
rect 17207 14055 17657 14077
rect 18311 14077 18455 14111
rect 18489 14077 18761 14111
rect 18919 14113 19195 14147
rect 19229 14113 19373 14147
rect 19995 14151 20061 14167
rect 18919 14097 19373 14113
rect 19415 14111 19865 14127
rect 18311 14055 18761 14077
rect 19415 14077 19559 14111
rect 19593 14077 19865 14111
rect 19995 14117 20011 14151
rect 20045 14117 20061 14151
rect 19995 14101 20061 14117
rect 20103 14111 20169 14127
rect 19415 14055 19865 14077
rect 20103 14077 20119 14111
rect 20153 14077 20169 14111
rect 20103 14061 20169 14077
rect 20103 14059 20141 14061
rect 16431 14028 16467 14052
rect 16711 14029 17657 14055
rect 17815 14029 18761 14055
rect 18919 14029 19865 14055
rect 20023 14029 20141 14059
rect 16431 14013 16461 14028
rect 15833 13978 15863 14010
rect 15348 13868 15378 13894
rect 15451 13868 15481 13894
rect 15665 13868 15695 13894
rect 15737 13868 15767 13894
rect 15833 13868 15863 13894
rect 12019 13829 12049 13855
rect 12107 13829 12137 13855
rect 12313 13829 12343 13855
rect 12399 13829 12429 13855
rect 12485 13829 12515 13855
rect 12571 13829 12601 13855
rect 12657 13829 12687 13855
rect 12743 13829 12773 13855
rect 12829 13829 12859 13855
rect 12915 13829 12945 13855
rect 13000 13829 13030 13855
rect 13086 13829 13116 13855
rect 13172 13829 13202 13855
rect 13258 13829 13288 13855
rect 13344 13829 13374 13855
rect 13430 13829 13460 13855
rect 13516 13829 13546 13855
rect 13602 13829 13632 13855
rect 13688 13829 13718 13855
rect 13774 13829 13804 13855
rect 13860 13829 13890 13855
rect 13946 13829 13976 13855
rect 14341 13829 14371 13855
rect 14425 13829 14525 13855
rect 14683 13829 14783 13855
rect 14848 13829 14878 13855
rect 15239 13829 15269 13855
rect 16067 13829 16097 13855
rect 16155 13829 16185 13855
rect 16343 13829 16373 13855
rect 16431 13829 16461 13855
rect 16711 13829 17657 13855
rect 17815 13829 18761 13855
rect 18919 13829 19865 13855
rect 20023 13829 20141 13855
rect 5027 13761 5145 13787
rect 5487 13761 6065 13787
rect 6223 13761 7169 13787
rect 7511 13761 8457 13787
rect 8615 13761 9561 13787
rect 9719 13761 9749 13787
rect 9807 13761 9837 13787
rect 10013 13761 10043 13787
rect 10099 13761 10129 13787
rect 10185 13761 10215 13787
rect 10271 13761 10301 13787
rect 10357 13761 10387 13787
rect 10443 13761 10473 13787
rect 10529 13761 10559 13787
rect 10615 13761 10645 13787
rect 10700 13761 10730 13787
rect 10786 13761 10816 13787
rect 10872 13761 10902 13787
rect 10958 13761 10988 13787
rect 11044 13761 11074 13787
rect 11130 13761 11160 13787
rect 11216 13761 11246 13787
rect 11302 13761 11332 13787
rect 11388 13761 11418 13787
rect 11474 13761 11504 13787
rect 11560 13761 11590 13787
rect 11646 13761 11676 13787
rect 11927 13761 12321 13787
rect 12571 13761 12601 13787
rect 12659 13761 12689 13787
rect 12939 13761 12969 13787
rect 13154 13761 13184 13787
rect 13238 13761 13268 13787
rect 13346 13761 13376 13787
rect 13430 13761 13460 13787
rect 13516 13761 13546 13787
rect 13615 13761 13645 13787
rect 13812 13761 13842 13787
rect 13909 13761 13939 13787
rect 14049 13761 14079 13787
rect 14148 13761 14178 13787
rect 14240 13761 14270 13787
rect 5027 13557 5145 13587
rect 5487 13561 6065 13587
rect 6223 13561 7169 13587
rect 9719 13588 9749 13603
rect 7511 13561 8457 13587
rect 8615 13561 9561 13587
rect 5027 13555 5065 13557
rect 4999 13539 5065 13555
rect 4999 13505 5015 13539
rect 5049 13505 5065 13539
rect 5801 13539 6065 13561
rect 4999 13489 5065 13505
rect 5107 13499 5173 13515
rect 5107 13465 5123 13499
rect 5157 13465 5173 13499
rect 5107 13449 5173 13465
rect 5487 13503 5759 13519
rect 5487 13469 5503 13503
rect 5537 13469 5606 13503
rect 5640 13469 5709 13503
rect 5743 13469 5759 13503
rect 5801 13505 5817 13539
rect 5851 13505 5916 13539
rect 5950 13505 6015 13539
rect 6049 13505 6065 13539
rect 6719 13539 7169 13561
rect 5801 13489 6065 13505
rect 6223 13503 6677 13519
rect 5107 13447 5145 13449
rect 5027 13421 5145 13447
rect 5487 13447 5759 13469
rect 6223 13469 6499 13503
rect 6533 13469 6677 13503
rect 6719 13505 6863 13539
rect 6897 13505 7169 13539
rect 8007 13539 8457 13561
rect 6719 13489 7169 13505
rect 7511 13503 7965 13519
rect 6223 13447 6677 13469
rect 7511 13469 7787 13503
rect 7821 13469 7965 13503
rect 8007 13505 8151 13539
rect 8185 13505 8457 13539
rect 9111 13539 9561 13561
rect 8007 13489 8457 13505
rect 8615 13503 9069 13519
rect 7511 13447 7965 13469
rect 8615 13469 8891 13503
rect 8925 13469 9069 13503
rect 9111 13505 9255 13539
rect 9289 13505 9561 13539
rect 9713 13564 9749 13588
rect 9713 13529 9743 13564
rect 9807 13542 9837 13603
rect 11927 13561 12321 13587
rect 9111 13489 9561 13505
rect 9667 13513 9743 13529
rect 8615 13447 9069 13469
rect 9667 13479 9677 13513
rect 9711 13479 9743 13513
rect 9667 13463 9743 13479
rect 9787 13526 9841 13542
rect 9787 13492 9797 13526
rect 9831 13492 9841 13526
rect 9787 13476 9841 13492
rect 10013 13529 10043 13561
rect 10099 13529 10129 13561
rect 10185 13529 10215 13561
rect 10271 13529 10301 13561
rect 10357 13529 10387 13561
rect 10443 13529 10473 13561
rect 10529 13529 10559 13561
rect 10615 13529 10645 13561
rect 10700 13529 10730 13561
rect 10786 13529 10816 13561
rect 10872 13529 10902 13561
rect 10958 13529 10988 13561
rect 11044 13529 11074 13561
rect 11130 13529 11160 13561
rect 11216 13529 11246 13561
rect 11302 13529 11332 13561
rect 10013 13513 11332 13529
rect 10013 13479 10238 13513
rect 10272 13479 10306 13513
rect 10340 13479 10374 13513
rect 10408 13479 10442 13513
rect 10476 13479 10510 13513
rect 10544 13479 10578 13513
rect 10612 13479 10646 13513
rect 10680 13479 10714 13513
rect 10748 13479 10782 13513
rect 10816 13479 10850 13513
rect 10884 13479 10918 13513
rect 10952 13479 10986 13513
rect 11020 13479 11054 13513
rect 11088 13479 11122 13513
rect 11156 13479 11190 13513
rect 11224 13479 11258 13513
rect 11292 13479 11332 13513
rect 9713 13454 9743 13463
rect 5487 13421 6065 13447
rect 6223 13421 7169 13447
rect 7511 13421 8457 13447
rect 8615 13421 9561 13447
rect 9713 13430 9749 13454
rect 9719 13415 9749 13430
rect 9807 13415 9837 13476
rect 10013 13454 11332 13479
rect 10013 13395 10043 13454
rect 10099 13395 10129 13454
rect 10185 13395 10215 13454
rect 10271 13395 10301 13454
rect 10357 13395 10387 13454
rect 10443 13395 10473 13454
rect 10529 13395 10559 13454
rect 10615 13395 10645 13454
rect 10700 13395 10730 13454
rect 10786 13395 10816 13454
rect 10872 13395 10902 13454
rect 10958 13395 10988 13454
rect 11044 13395 11074 13454
rect 11130 13395 11160 13454
rect 11216 13395 11246 13454
rect 11302 13395 11332 13454
rect 11388 13546 11418 13561
rect 11474 13546 11504 13561
rect 11560 13546 11590 13561
rect 11646 13546 11676 13561
rect 11388 13513 11735 13546
rect 12145 13539 12321 13561
rect 12571 13542 12601 13603
rect 12659 13588 12689 13603
rect 12659 13564 12695 13588
rect 11388 13479 11685 13513
rect 11719 13479 11735 13513
rect 11388 13444 11735 13479
rect 11927 13503 12103 13519
rect 11927 13469 11943 13503
rect 11977 13469 12053 13503
rect 12087 13469 12103 13503
rect 12145 13505 12161 13539
rect 12195 13505 12271 13539
rect 12305 13505 12321 13539
rect 12145 13489 12321 13505
rect 12567 13526 12621 13542
rect 12567 13492 12577 13526
rect 12611 13492 12621 13526
rect 12567 13476 12621 13492
rect 12665 13529 12695 13564
rect 13154 13629 13184 13677
rect 13142 13613 13196 13629
rect 13142 13579 13152 13613
rect 13186 13579 13196 13613
rect 13142 13563 13196 13579
rect 12939 13529 12969 13561
rect 12665 13513 12741 13529
rect 12665 13479 12697 13513
rect 12731 13479 12741 13513
rect 11927 13447 12103 13469
rect 11388 13395 11418 13444
rect 11474 13395 11504 13444
rect 11560 13395 11590 13444
rect 11646 13395 11676 13444
rect 11927 13421 12321 13447
rect 12571 13415 12601 13476
rect 12665 13463 12741 13479
rect 12939 13513 12998 13529
rect 12939 13479 12954 13513
rect 12988 13479 12998 13513
rect 12939 13463 12998 13479
rect 12665 13454 12695 13463
rect 12659 13430 12695 13454
rect 12939 13441 12969 13463
rect 12659 13415 12689 13430
rect 13147 13395 13177 13563
rect 13238 13521 13268 13677
rect 13219 13505 13273 13521
rect 13219 13471 13229 13505
rect 13263 13471 13273 13505
rect 13346 13493 13376 13677
rect 13430 13645 13460 13677
rect 13420 13629 13474 13645
rect 13420 13595 13430 13629
rect 13464 13595 13474 13629
rect 13420 13579 13474 13595
rect 13516 13543 13546 13677
rect 14507 13755 14537 13781
rect 14591 13755 14621 13781
rect 14780 13761 14810 13787
rect 14866 13761 14896 13787
rect 14952 13761 14982 13787
rect 15038 13761 15068 13787
rect 15124 13761 15154 13787
rect 15210 13761 15240 13787
rect 15296 13761 15326 13787
rect 15382 13761 15412 13787
rect 15468 13761 15498 13787
rect 15554 13761 15584 13787
rect 15640 13761 15670 13787
rect 15726 13761 15756 13787
rect 15811 13761 15841 13787
rect 15897 13761 15927 13787
rect 15983 13761 16013 13787
rect 16069 13761 16099 13787
rect 16155 13761 16185 13787
rect 16241 13761 16271 13787
rect 16327 13761 16357 13787
rect 16413 13761 16443 13787
rect 16619 13761 16649 13787
rect 17815 13761 18761 13787
rect 18919 13761 19865 13787
rect 20023 13761 20141 13787
rect 13615 13578 13645 13593
rect 13615 13548 13721 13578
rect 13496 13531 13546 13543
rect 13483 13519 13546 13531
rect 13219 13455 13273 13471
rect 13315 13477 13376 13493
rect 13238 13395 13268 13455
rect 13315 13443 13325 13477
rect 13359 13457 13376 13477
rect 13459 13513 13546 13519
rect 13691 13531 13721 13548
rect 13691 13515 13757 13531
rect 13459 13503 13525 13513
rect 13459 13469 13469 13503
rect 13503 13501 13525 13503
rect 13503 13469 13513 13501
rect 13691 13481 13713 13515
rect 13747 13481 13757 13515
rect 13812 13483 13842 13677
rect 13909 13619 13939 13677
rect 13884 13603 13939 13619
rect 13884 13569 13895 13603
rect 13929 13569 13939 13603
rect 13884 13553 13939 13569
rect 13359 13443 13417 13457
rect 13459 13453 13513 13469
rect 13315 13427 13417 13443
rect 13387 13395 13417 13427
rect 13483 13383 13513 13453
rect 13555 13455 13622 13471
rect 13555 13421 13565 13455
rect 13599 13421 13622 13455
rect 13691 13465 13757 13481
rect 13799 13467 13853 13483
rect 13691 13439 13721 13465
rect 13555 13405 13622 13421
rect 13592 13383 13622 13405
rect 13799 13433 13809 13467
rect 13843 13433 13853 13467
rect 13799 13417 13853 13433
rect 13823 13395 13853 13417
rect 13895 13395 13925 13553
rect 14049 13543 14079 13677
rect 14148 13639 14178 13677
rect 14128 13629 14194 13639
rect 14128 13595 14144 13629
rect 14178 13595 14194 13629
rect 14128 13585 14194 13595
rect 14240 13590 14270 13677
rect 14240 13574 14369 13590
rect 14240 13560 14325 13574
rect 14049 13513 14187 13543
rect 14156 13483 14187 13513
rect 14252 13540 14325 13560
rect 14359 13540 14369 13574
rect 14252 13524 14369 13540
rect 14507 13538 14537 13627
rect 14591 13612 14621 13627
rect 14591 13582 14654 13612
rect 14507 13528 14582 13538
rect 14048 13461 14114 13471
rect 14048 13427 14064 13461
rect 14098 13427 14114 13461
rect 14048 13417 14114 13427
rect 14156 13467 14210 13483
rect 14156 13433 14166 13467
rect 14200 13433 14210 13467
rect 14156 13417 14210 13433
rect 14061 13383 14091 13417
rect 14157 13383 14187 13417
rect 14252 13395 14282 13524
rect 14507 13494 14532 13528
rect 14566 13494 14582 13528
rect 14507 13484 14582 13494
rect 14624 13529 14654 13582
rect 16728 13722 16758 13748
rect 16831 13722 16861 13748
rect 17045 13722 17075 13748
rect 17117 13722 17147 13748
rect 17213 13722 17243 13748
rect 14780 13546 14810 13561
rect 14866 13546 14896 13561
rect 14952 13546 14982 13561
rect 15038 13546 15068 13561
rect 14624 13513 14678 13529
rect 14507 13395 14537 13484
rect 14624 13479 14634 13513
rect 14668 13479 14678 13513
rect 14624 13463 14678 13479
rect 14721 13513 15068 13546
rect 14721 13479 14737 13513
rect 14771 13479 15068 13513
rect 14624 13440 14654 13463
rect 14721 13444 15068 13479
rect 14591 13410 14654 13440
rect 14591 13395 14621 13410
rect 14780 13395 14810 13444
rect 14866 13395 14896 13444
rect 14952 13395 14982 13444
rect 15038 13395 15068 13444
rect 15124 13529 15154 13561
rect 15210 13529 15240 13561
rect 15296 13529 15326 13561
rect 15382 13529 15412 13561
rect 15468 13529 15498 13561
rect 15554 13529 15584 13561
rect 15640 13529 15670 13561
rect 15726 13529 15756 13561
rect 15811 13529 15841 13561
rect 15897 13529 15927 13561
rect 15983 13529 16013 13561
rect 16069 13529 16099 13561
rect 16155 13529 16185 13561
rect 16241 13529 16271 13561
rect 16327 13529 16357 13561
rect 16413 13529 16443 13561
rect 16619 13529 16649 13561
rect 16728 13529 16758 13638
rect 16831 13623 16861 13638
rect 16831 13593 16979 13623
rect 17045 13606 17075 13638
rect 15124 13513 16443 13529
rect 15124 13479 15164 13513
rect 15198 13479 15232 13513
rect 15266 13479 15300 13513
rect 15334 13479 15368 13513
rect 15402 13479 15436 13513
rect 15470 13479 15504 13513
rect 15538 13479 15572 13513
rect 15606 13479 15640 13513
rect 15674 13479 15708 13513
rect 15742 13479 15776 13513
rect 15810 13479 15844 13513
rect 15878 13479 15912 13513
rect 15946 13479 15980 13513
rect 16014 13479 16048 13513
rect 16082 13479 16116 13513
rect 16150 13479 16184 13513
rect 16218 13479 16443 13513
rect 15124 13454 16443 13479
rect 16616 13513 16670 13529
rect 16616 13479 16626 13513
rect 16660 13479 16670 13513
rect 16616 13463 16670 13479
rect 16712 13513 16766 13529
rect 16712 13479 16722 13513
rect 16756 13479 16766 13513
rect 16949 13493 16979 13593
rect 17021 13590 17075 13606
rect 17021 13556 17031 13590
rect 17065 13556 17075 13590
rect 17021 13540 17075 13556
rect 16712 13463 16766 13479
rect 16824 13477 16907 13493
rect 15124 13395 15154 13454
rect 15210 13395 15240 13454
rect 15296 13395 15326 13454
rect 15382 13395 15412 13454
rect 15468 13395 15498 13454
rect 15554 13395 15584 13454
rect 15640 13395 15670 13454
rect 15726 13395 15756 13454
rect 15811 13395 15841 13454
rect 15897 13395 15927 13454
rect 15983 13395 16013 13454
rect 16069 13395 16099 13454
rect 16155 13395 16185 13454
rect 16241 13395 16271 13454
rect 16327 13395 16357 13454
rect 16413 13395 16443 13454
rect 16619 13441 16649 13463
rect 16728 13395 16758 13463
rect 16824 13443 16863 13477
rect 16897 13443 16907 13477
rect 16824 13427 16907 13443
rect 16949 13477 17003 13493
rect 17117 13487 17147 13638
rect 17213 13606 17243 13638
rect 17189 13590 17243 13606
rect 17189 13556 17199 13590
rect 17233 13556 17243 13590
rect 17815 13561 18761 13587
rect 18919 13561 19865 13587
rect 17189 13540 17243 13556
rect 16949 13443 16959 13477
rect 16993 13443 17003 13477
rect 17105 13477 17171 13487
rect 17105 13463 17121 13477
rect 16949 13427 17003 13443
rect 17045 13443 17121 13463
rect 17155 13443 17171 13477
rect 17045 13433 17171 13443
rect 16824 13395 16854 13427
rect 16949 13395 16979 13427
rect 17045 13395 17075 13433
rect 17213 13395 17243 13540
rect 18311 13539 18761 13561
rect 17815 13503 18269 13519
rect 17815 13469 18091 13503
rect 18125 13469 18269 13503
rect 18311 13505 18455 13539
rect 18489 13505 18761 13539
rect 19415 13539 19865 13561
rect 20023 13557 20141 13587
rect 18311 13489 18761 13505
rect 18919 13503 19373 13519
rect 17815 13447 18269 13469
rect 18919 13469 19195 13503
rect 19229 13469 19373 13503
rect 19415 13505 19559 13539
rect 19593 13505 19865 13539
rect 20103 13555 20141 13557
rect 20103 13539 20169 13555
rect 19415 13489 19865 13505
rect 19995 13499 20061 13515
rect 18919 13447 19373 13469
rect 19995 13465 20011 13499
rect 20045 13465 20061 13499
rect 20103 13505 20119 13539
rect 20153 13505 20169 13539
rect 20103 13489 20169 13505
rect 19995 13449 20061 13465
rect 20023 13447 20061 13449
rect 17815 13421 18761 13447
rect 18919 13421 19865 13447
rect 20023 13421 20141 13447
rect 5027 13285 5145 13311
rect 5487 13285 6065 13311
rect 6223 13285 7169 13311
rect 7511 13285 8457 13311
rect 8615 13285 9561 13311
rect 9719 13285 9749 13311
rect 9807 13285 9837 13311
rect 10013 13285 10043 13311
rect 10099 13285 10129 13311
rect 10185 13285 10215 13311
rect 10271 13285 10301 13311
rect 10357 13285 10387 13311
rect 10443 13285 10473 13311
rect 10529 13285 10559 13311
rect 10615 13285 10645 13311
rect 10700 13285 10730 13311
rect 10786 13285 10816 13311
rect 10872 13285 10902 13311
rect 10958 13285 10988 13311
rect 11044 13285 11074 13311
rect 11130 13285 11160 13311
rect 11216 13285 11246 13311
rect 11302 13285 11332 13311
rect 11388 13285 11418 13311
rect 11474 13285 11504 13311
rect 11560 13285 11590 13311
rect 11646 13285 11676 13311
rect 11927 13285 12321 13311
rect 12571 13285 12601 13311
rect 12659 13285 12689 13311
rect 12939 13285 12969 13311
rect 13147 13285 13177 13311
rect 13238 13285 13268 13311
rect 13387 13285 13417 13311
rect 13483 13285 13513 13311
rect 13592 13285 13622 13311
rect 13691 13285 13721 13311
rect 13823 13285 13853 13311
rect 13895 13285 13925 13311
rect 14061 13285 14091 13311
rect 14157 13285 14187 13311
rect 14252 13285 14282 13311
rect 14507 13285 14537 13311
rect 14591 13285 14621 13311
rect 14780 13285 14810 13311
rect 14866 13285 14896 13311
rect 14952 13285 14982 13311
rect 15038 13285 15068 13311
rect 15124 13285 15154 13311
rect 15210 13285 15240 13311
rect 15296 13285 15326 13311
rect 15382 13285 15412 13311
rect 15468 13285 15498 13311
rect 15554 13285 15584 13311
rect 15640 13285 15670 13311
rect 15726 13285 15756 13311
rect 15811 13285 15841 13311
rect 15897 13285 15927 13311
rect 15983 13285 16013 13311
rect 16069 13285 16099 13311
rect 16155 13285 16185 13311
rect 16241 13285 16271 13311
rect 16327 13285 16357 13311
rect 16413 13285 16443 13311
rect 16619 13285 16649 13311
rect 16728 13285 16758 13311
rect 16824 13285 16854 13311
rect 16949 13285 16979 13311
rect 17045 13285 17075 13311
rect 17213 13285 17243 13311
rect 17815 13285 18761 13311
rect 18919 13285 19865 13311
rect 20023 13285 20141 13311
rect 5027 13217 5145 13243
rect 5303 13217 5697 13243
rect 5855 13217 6801 13243
rect 6959 13217 7905 13243
rect 8063 13217 9009 13243
rect 9189 13217 9219 13243
rect 9273 13217 9373 13243
rect 9531 13217 9631 13243
rect 9696 13217 9726 13243
rect 10087 13217 10297 13243
rect 10455 13217 10485 13243
rect 10663 13217 10693 13243
rect 10754 13217 10784 13243
rect 10903 13217 10933 13243
rect 10999 13217 11029 13243
rect 11108 13217 11138 13243
rect 11207 13217 11237 13243
rect 11339 13217 11369 13243
rect 11411 13217 11441 13243
rect 11577 13217 11607 13243
rect 11673 13217 11703 13243
rect 11768 13217 11798 13243
rect 12023 13217 12053 13243
rect 12107 13217 12137 13243
rect 12295 13217 12325 13243
rect 12379 13217 12409 13243
rect 12634 13217 12664 13243
rect 12729 13217 12759 13243
rect 12825 13217 12855 13243
rect 12991 13217 13021 13243
rect 13063 13217 13093 13243
rect 13195 13217 13225 13243
rect 13294 13217 13324 13243
rect 13403 13217 13433 13243
rect 13499 13217 13529 13243
rect 13648 13217 13678 13243
rect 13739 13217 13769 13243
rect 13947 13217 13977 13243
rect 14135 13217 14165 13243
rect 14244 13217 14274 13243
rect 14340 13217 14370 13243
rect 14465 13217 14495 13243
rect 14561 13217 14591 13243
rect 14729 13217 14759 13243
rect 15147 13217 15177 13243
rect 15355 13217 15385 13243
rect 15446 13217 15476 13243
rect 15595 13217 15625 13243
rect 15691 13217 15721 13243
rect 15800 13217 15830 13243
rect 15899 13217 15929 13243
rect 16031 13217 16061 13243
rect 16103 13217 16133 13243
rect 16269 13217 16299 13243
rect 16365 13217 16395 13243
rect 16460 13217 16490 13243
rect 16715 13217 16745 13243
rect 16799 13217 16829 13243
rect 17006 13217 17036 13243
rect 17101 13217 17201 13243
rect 17359 13217 17459 13243
rect 17513 13217 17543 13243
rect 17815 13217 18761 13243
rect 18919 13217 19865 13243
rect 20023 13217 20141 13243
rect 5027 13081 5145 13107
rect 5107 13079 5145 13081
rect 5303 13081 5697 13107
rect 5855 13081 6801 13107
rect 6959 13081 7905 13107
rect 8063 13081 9009 13107
rect 5107 13063 5173 13079
rect 4999 13023 5065 13039
rect 4999 12989 5015 13023
rect 5049 12989 5065 13023
rect 5107 13029 5123 13063
rect 5157 13029 5173 13063
rect 5107 13013 5173 13029
rect 5303 13059 5479 13081
rect 5303 13025 5319 13059
rect 5353 13025 5429 13059
rect 5463 13025 5479 13059
rect 5855 13059 6309 13081
rect 5303 13009 5479 13025
rect 5521 13023 5697 13039
rect 4999 12973 5065 12989
rect 5027 12971 5065 12973
rect 5521 12989 5537 13023
rect 5571 12989 5647 13023
rect 5681 12989 5697 13023
rect 5855 13025 6131 13059
rect 6165 13025 6309 13059
rect 6959 13059 7413 13081
rect 5855 13009 6309 13025
rect 6351 13023 6801 13039
rect 5027 12941 5145 12971
rect 5521 12967 5697 12989
rect 6351 12989 6495 13023
rect 6529 12989 6801 13023
rect 6959 13025 7235 13059
rect 7269 13025 7413 13059
rect 8063 13059 8517 13081
rect 9189 13065 9219 13133
rect 6959 13009 7413 13025
rect 7455 13023 7905 13039
rect 6351 12967 6801 12989
rect 7455 12989 7599 13023
rect 7633 12989 7905 13023
rect 8063 13025 8339 13059
rect 8373 13025 8517 13059
rect 9159 13049 9219 13065
rect 8063 13009 8517 13025
rect 8559 13023 9009 13039
rect 7455 12967 7905 12989
rect 8559 12989 8703 13023
rect 8737 12989 9009 13023
rect 9159 13015 9169 13049
rect 9203 13015 9219 13049
rect 9159 12999 9219 13015
rect 8559 12967 9009 12989
rect 5303 12941 5697 12967
rect 5855 12941 6801 12967
rect 6959 12941 7905 12967
rect 8063 12941 9009 12967
rect 9189 12851 9219 12999
rect 9273 13049 9373 13133
rect 9531 13065 9631 13133
rect 9696 13065 9726 13087
rect 10087 13081 10297 13107
rect 10087 13075 10171 13081
rect 9273 13015 9283 13049
rect 9317 13015 9373 13049
rect 9273 12851 9373 13015
rect 9477 13049 9631 13065
rect 9477 13015 9487 13049
rect 9521 13015 9631 13049
rect 9477 12999 9631 13015
rect 9673 13049 9727 13065
rect 9673 13015 9683 13049
rect 9717 13015 9727 13049
rect 9673 12999 9727 13015
rect 10029 13059 10171 13075
rect 10029 13025 10045 13059
rect 10079 13025 10171 13059
rect 10455 13065 10485 13087
rect 10455 13049 10514 13065
rect 10029 13009 10171 13025
rect 10213 13023 10355 13039
rect 9531 12851 9631 12999
rect 9696 12967 9726 12999
rect 10213 12989 10305 13023
rect 10339 12989 10355 13023
rect 10213 12973 10355 12989
rect 10455 13015 10470 13049
rect 10504 13015 10514 13049
rect 10455 12999 10514 13015
rect 10213 12967 10297 12973
rect 10455 12967 10485 12999
rect 10087 12941 10297 12967
rect 10663 12965 10693 13133
rect 10754 13073 10784 13133
rect 10903 13101 10933 13133
rect 10831 13085 10933 13101
rect 10735 13057 10789 13073
rect 10735 13023 10745 13057
rect 10779 13023 10789 13057
rect 10831 13051 10841 13085
rect 10875 13071 10933 13085
rect 10999 13075 11029 13145
rect 11108 13123 11138 13145
rect 10875 13051 10892 13071
rect 10831 13035 10892 13051
rect 10735 13007 10789 13023
rect 10658 12949 10712 12965
rect 10658 12915 10668 12949
rect 10702 12915 10712 12949
rect 10658 12899 10712 12915
rect 10670 12851 10700 12899
rect 10754 12851 10784 13007
rect 10862 12851 10892 13035
rect 10975 13059 11029 13075
rect 10975 13025 10985 13059
rect 11019 13027 11029 13059
rect 11071 13107 11138 13123
rect 11071 13073 11081 13107
rect 11115 13073 11138 13107
rect 11339 13111 11369 13133
rect 11315 13095 11369 13111
rect 11071 13057 11138 13073
rect 11207 13063 11237 13089
rect 11207 13047 11273 13063
rect 11019 13025 11041 13027
rect 10975 13015 11041 13025
rect 10975 13009 11062 13015
rect 10999 12997 11062 13009
rect 11012 12985 11062 12997
rect 10936 12933 10990 12949
rect 10936 12899 10946 12933
rect 10980 12899 10990 12933
rect 10936 12883 10990 12899
rect 10946 12851 10976 12883
rect 11032 12851 11062 12985
rect 11207 13013 11229 13047
rect 11263 13013 11273 13047
rect 11315 13061 11325 13095
rect 11359 13061 11369 13095
rect 11315 13045 11369 13061
rect 11207 12997 11273 13013
rect 11207 12980 11237 12997
rect 11131 12950 11237 12980
rect 11131 12935 11161 12950
rect 11328 12851 11358 13045
rect 11411 12975 11441 13133
rect 11577 13111 11607 13145
rect 11673 13111 11703 13145
rect 11564 13101 11630 13111
rect 11564 13067 11580 13101
rect 11614 13067 11630 13101
rect 11564 13057 11630 13067
rect 11672 13095 11726 13111
rect 11672 13061 11682 13095
rect 11716 13061 11726 13095
rect 11672 13045 11726 13061
rect 11672 13015 11703 13045
rect 11565 12985 11703 13015
rect 11768 13004 11798 13133
rect 12023 13044 12053 13133
rect 12107 13118 12137 13133
rect 12295 13118 12325 13133
rect 12107 13088 12170 13118
rect 12140 13065 12170 13088
rect 12262 13088 12325 13118
rect 12262 13065 12292 13088
rect 12140 13049 12194 13065
rect 12023 13034 12098 13044
rect 11768 12988 11885 13004
rect 11400 12959 11455 12975
rect 11400 12925 11411 12959
rect 11445 12925 11455 12959
rect 11400 12909 11455 12925
rect 11425 12851 11455 12909
rect 11565 12851 11595 12985
rect 11768 12968 11841 12988
rect 11756 12954 11841 12968
rect 11875 12954 11885 12988
rect 11644 12933 11710 12943
rect 11644 12899 11660 12933
rect 11694 12899 11710 12933
rect 11644 12889 11710 12899
rect 11756 12938 11885 12954
rect 12023 13000 12048 13034
rect 12082 13000 12098 13034
rect 12023 12990 12098 13000
rect 12140 13015 12150 13049
rect 12184 13015 12194 13049
rect 12140 12999 12194 13015
rect 12238 13049 12292 13065
rect 12238 13015 12248 13049
rect 12282 13015 12292 13049
rect 12379 13044 12409 13133
rect 12238 12999 12292 13015
rect 11664 12851 11694 12889
rect 11756 12851 11786 12938
rect 12023 12901 12053 12990
rect 12140 12946 12170 12999
rect 12107 12916 12170 12946
rect 12262 12946 12292 12999
rect 12334 13034 12409 13044
rect 12334 13000 12350 13034
rect 12384 13000 12409 13034
rect 12634 13004 12664 13133
rect 12729 13111 12759 13145
rect 12825 13111 12855 13145
rect 12706 13095 12760 13111
rect 12706 13061 12716 13095
rect 12750 13061 12760 13095
rect 12706 13045 12760 13061
rect 12802 13101 12868 13111
rect 12802 13067 12818 13101
rect 12852 13067 12868 13101
rect 12802 13057 12868 13067
rect 12334 12990 12409 13000
rect 12262 12916 12325 12946
rect 12107 12901 12137 12916
rect 12295 12901 12325 12916
rect 12379 12901 12409 12990
rect 12547 12988 12664 13004
rect 12547 12954 12557 12988
rect 12591 12968 12664 12988
rect 12729 13015 12760 13045
rect 12729 12985 12867 13015
rect 12591 12954 12676 12968
rect 12547 12938 12676 12954
rect 12646 12851 12676 12938
rect 12722 12933 12788 12943
rect 12722 12899 12738 12933
rect 12772 12899 12788 12933
rect 12722 12889 12788 12899
rect 12738 12851 12768 12889
rect 12837 12851 12867 12985
rect 12991 12975 13021 13133
rect 13063 13111 13093 13133
rect 13063 13095 13117 13111
rect 13063 13061 13073 13095
rect 13107 13061 13117 13095
rect 13294 13123 13324 13145
rect 13294 13107 13361 13123
rect 13195 13063 13225 13089
rect 13063 13045 13117 13061
rect 13159 13047 13225 13063
rect 13294 13073 13317 13107
rect 13351 13073 13361 13107
rect 13294 13057 13361 13073
rect 13403 13075 13433 13145
rect 13499 13101 13529 13133
rect 13499 13085 13601 13101
rect 13403 13059 13457 13075
rect 13499 13071 13557 13085
rect 12977 12959 13032 12975
rect 12977 12925 12987 12959
rect 13021 12925 13032 12959
rect 12977 12909 13032 12925
rect 12977 12851 13007 12909
rect 13074 12851 13104 13045
rect 13159 13013 13169 13047
rect 13203 13013 13225 13047
rect 13403 13027 13413 13059
rect 13391 13025 13413 13027
rect 13447 13025 13457 13059
rect 13391 13015 13457 13025
rect 13159 12997 13225 13013
rect 13195 12980 13225 12997
rect 13370 13009 13457 13015
rect 13540 13051 13557 13071
rect 13591 13051 13601 13085
rect 13648 13073 13678 13133
rect 13540 13035 13601 13051
rect 13643 13057 13697 13073
rect 13370 12997 13433 13009
rect 13370 12985 13420 12997
rect 13195 12950 13301 12980
rect 13271 12935 13301 12950
rect 5027 12741 5145 12767
rect 5303 12741 5697 12767
rect 5855 12741 6801 12767
rect 6959 12741 7905 12767
rect 8063 12741 9009 12767
rect 9189 12741 9219 12767
rect 9273 12741 9373 12767
rect 9531 12741 9631 12767
rect 9696 12741 9726 12767
rect 10087 12741 10297 12767
rect 10455 12741 10485 12767
rect 10670 12741 10700 12767
rect 10754 12741 10784 12767
rect 10862 12741 10892 12767
rect 10946 12741 10976 12767
rect 11032 12741 11062 12767
rect 11131 12741 11161 12767
rect 11328 12741 11358 12767
rect 11425 12741 11455 12767
rect 11565 12741 11595 12767
rect 11664 12741 11694 12767
rect 11756 12741 11786 12767
rect 12023 12747 12053 12773
rect 12107 12747 12137 12773
rect 12295 12747 12325 12773
rect 12379 12747 12409 12773
rect 13370 12851 13400 12985
rect 13442 12933 13496 12949
rect 13442 12899 13452 12933
rect 13486 12899 13496 12933
rect 13442 12883 13496 12899
rect 13456 12851 13486 12883
rect 13540 12851 13570 13035
rect 13643 13023 13653 13057
rect 13687 13023 13697 13057
rect 13643 13007 13697 13023
rect 13648 12851 13678 13007
rect 13739 12965 13769 13133
rect 13947 13065 13977 13087
rect 14135 13065 14165 13087
rect 14244 13065 14274 13133
rect 14340 13101 14370 13133
rect 14465 13101 14495 13133
rect 14340 13085 14423 13101
rect 13918 13049 13977 13065
rect 13918 13015 13928 13049
rect 13962 13015 13977 13049
rect 13918 12999 13977 13015
rect 14132 13049 14186 13065
rect 14132 13015 14142 13049
rect 14176 13015 14186 13049
rect 14132 12999 14186 13015
rect 14228 13049 14282 13065
rect 14228 13015 14238 13049
rect 14272 13015 14282 13049
rect 14340 13051 14379 13085
rect 14413 13051 14423 13085
rect 14340 13035 14423 13051
rect 14465 13085 14519 13101
rect 14465 13051 14475 13085
rect 14509 13051 14519 13085
rect 14561 13095 14591 13133
rect 14561 13085 14687 13095
rect 14561 13065 14637 13085
rect 14465 13035 14519 13051
rect 14621 13051 14637 13065
rect 14671 13051 14687 13085
rect 14621 13041 14687 13051
rect 14228 12999 14282 13015
rect 13947 12967 13977 12999
rect 14135 12967 14165 12999
rect 13720 12949 13774 12965
rect 13720 12915 13730 12949
rect 13764 12915 13774 12949
rect 13720 12899 13774 12915
rect 13732 12851 13762 12899
rect 14244 12890 14274 12999
rect 14465 12935 14495 13035
rect 14347 12905 14495 12935
rect 14537 12972 14591 12988
rect 14537 12938 14547 12972
rect 14581 12938 14591 12972
rect 14537 12922 14591 12938
rect 14347 12890 14377 12905
rect 14561 12890 14591 12922
rect 14633 12890 14663 13041
rect 14729 12988 14759 13133
rect 14705 12972 14759 12988
rect 14705 12938 14715 12972
rect 14749 12938 14759 12972
rect 15147 13065 15177 13087
rect 15147 13049 15206 13065
rect 15147 13015 15162 13049
rect 15196 13015 15206 13049
rect 15147 12999 15206 13015
rect 15147 12967 15177 12999
rect 14705 12922 14759 12938
rect 14729 12890 14759 12922
rect 14244 12780 14274 12806
rect 14347 12780 14377 12806
rect 14561 12780 14591 12806
rect 14633 12780 14663 12806
rect 14729 12780 14759 12806
rect 15355 12965 15385 13133
rect 15446 13073 15476 13133
rect 15595 13101 15625 13133
rect 15523 13085 15625 13101
rect 15427 13057 15481 13073
rect 15427 13023 15437 13057
rect 15471 13023 15481 13057
rect 15523 13051 15533 13085
rect 15567 13071 15625 13085
rect 15691 13075 15721 13145
rect 15800 13123 15830 13145
rect 15567 13051 15584 13071
rect 15523 13035 15584 13051
rect 15427 13007 15481 13023
rect 15350 12949 15404 12965
rect 15350 12915 15360 12949
rect 15394 12915 15404 12949
rect 15350 12899 15404 12915
rect 15362 12851 15392 12899
rect 15446 12851 15476 13007
rect 15554 12851 15584 13035
rect 15667 13059 15721 13075
rect 15667 13025 15677 13059
rect 15711 13027 15721 13059
rect 15763 13107 15830 13123
rect 15763 13073 15773 13107
rect 15807 13073 15830 13107
rect 16031 13111 16061 13133
rect 16007 13095 16061 13111
rect 15763 13057 15830 13073
rect 15899 13063 15929 13089
rect 15899 13047 15965 13063
rect 15711 13025 15733 13027
rect 15667 13015 15733 13025
rect 15667 13009 15754 13015
rect 15691 12997 15754 13009
rect 15704 12985 15754 12997
rect 15628 12933 15682 12949
rect 15628 12899 15638 12933
rect 15672 12899 15682 12933
rect 15628 12883 15682 12899
rect 15638 12851 15668 12883
rect 15724 12851 15754 12985
rect 15899 13013 15921 13047
rect 15955 13013 15965 13047
rect 16007 13061 16017 13095
rect 16051 13061 16061 13095
rect 16007 13045 16061 13061
rect 15899 12997 15965 13013
rect 15899 12980 15929 12997
rect 15823 12950 15929 12980
rect 15823 12935 15853 12950
rect 16020 12851 16050 13045
rect 16103 12975 16133 13133
rect 16269 13111 16299 13145
rect 16365 13111 16395 13145
rect 16256 13101 16322 13111
rect 16256 13067 16272 13101
rect 16306 13067 16322 13101
rect 16256 13057 16322 13067
rect 16364 13095 16418 13111
rect 16364 13061 16374 13095
rect 16408 13061 16418 13095
rect 16364 13045 16418 13061
rect 16364 13015 16395 13045
rect 16257 12985 16395 13015
rect 16460 13004 16490 13133
rect 16715 13044 16745 13133
rect 16799 13118 16829 13133
rect 16799 13088 16862 13118
rect 16832 13065 16862 13088
rect 17006 13065 17036 13087
rect 17101 13065 17201 13133
rect 16832 13049 16886 13065
rect 16715 13034 16790 13044
rect 16460 12988 16577 13004
rect 16092 12959 16147 12975
rect 16092 12925 16103 12959
rect 16137 12925 16147 12959
rect 16092 12909 16147 12925
rect 16117 12851 16147 12909
rect 16257 12851 16287 12985
rect 16460 12968 16533 12988
rect 16448 12954 16533 12968
rect 16567 12954 16577 12988
rect 16336 12933 16402 12943
rect 16336 12899 16352 12933
rect 16386 12899 16402 12933
rect 16336 12889 16402 12899
rect 16448 12938 16577 12954
rect 16715 13000 16740 13034
rect 16774 13000 16790 13034
rect 16715 12990 16790 13000
rect 16832 13015 16842 13049
rect 16876 13015 16886 13049
rect 16832 12999 16886 13015
rect 17005 13049 17059 13065
rect 17005 13015 17015 13049
rect 17049 13015 17059 13049
rect 17005 12999 17059 13015
rect 17101 13049 17255 13065
rect 17101 13015 17211 13049
rect 17245 13015 17255 13049
rect 17101 12999 17255 13015
rect 17359 13049 17459 13133
rect 17359 13015 17415 13049
rect 17449 13015 17459 13049
rect 16356 12851 16386 12889
rect 16448 12851 16478 12938
rect 16715 12901 16745 12990
rect 16832 12946 16862 12999
rect 17006 12967 17036 12999
rect 16799 12916 16862 12946
rect 16799 12901 16829 12916
rect 12646 12741 12676 12767
rect 12738 12741 12768 12767
rect 12837 12741 12867 12767
rect 12977 12741 13007 12767
rect 13074 12741 13104 12767
rect 13271 12741 13301 12767
rect 13370 12741 13400 12767
rect 13456 12741 13486 12767
rect 13540 12741 13570 12767
rect 13648 12741 13678 12767
rect 13732 12741 13762 12767
rect 13947 12741 13977 12767
rect 14135 12741 14165 12767
rect 15147 12741 15177 12767
rect 15362 12741 15392 12767
rect 15446 12741 15476 12767
rect 15554 12741 15584 12767
rect 15638 12741 15668 12767
rect 15724 12741 15754 12767
rect 15823 12741 15853 12767
rect 16020 12741 16050 12767
rect 16117 12741 16147 12767
rect 16257 12741 16287 12767
rect 16356 12741 16386 12767
rect 16448 12741 16478 12767
rect 16715 12747 16745 12773
rect 16799 12747 16829 12773
rect 17101 12851 17201 12999
rect 17359 12851 17459 13015
rect 17513 13065 17543 13133
rect 17815 13081 18761 13107
rect 18919 13081 19865 13107
rect 20023 13081 20141 13107
rect 17513 13049 17573 13065
rect 17513 13015 17529 13049
rect 17563 13015 17573 13049
rect 17513 12999 17573 13015
rect 17815 13059 18269 13081
rect 17815 13025 18091 13059
rect 18125 13025 18269 13059
rect 18919 13059 19373 13081
rect 20023 13079 20061 13081
rect 17815 13009 18269 13025
rect 18311 13023 18761 13039
rect 17513 12851 17543 12999
rect 18311 12989 18455 13023
rect 18489 12989 18761 13023
rect 18919 13025 19195 13059
rect 19229 13025 19373 13059
rect 19995 13063 20061 13079
rect 18919 13009 19373 13025
rect 19415 13023 19865 13039
rect 18311 12967 18761 12989
rect 19415 12989 19559 13023
rect 19593 12989 19865 13023
rect 19995 13029 20011 13063
rect 20045 13029 20061 13063
rect 19995 13013 20061 13029
rect 20103 13023 20169 13039
rect 19415 12967 19865 12989
rect 20103 12989 20119 13023
rect 20153 12989 20169 13023
rect 20103 12973 20169 12989
rect 20103 12971 20141 12973
rect 17815 12941 18761 12967
rect 18919 12941 19865 12967
rect 20023 12941 20141 12971
rect 17006 12741 17036 12767
rect 17101 12741 17201 12767
rect 17359 12741 17459 12767
rect 17513 12741 17543 12767
rect 17815 12741 18761 12767
rect 18919 12741 19865 12767
rect 20023 12741 20141 12767
rect 5027 12673 5145 12699
rect 5245 12660 5341 12699
rect 5245 12626 5295 12660
rect 5329 12626 5341 12660
rect 5245 12592 5341 12626
rect 5245 12558 5295 12592
rect 5329 12558 5341 12592
rect 5027 12469 5145 12499
rect 5027 12467 5065 12469
rect 4999 12451 5065 12467
rect 4999 12417 5015 12451
rect 5049 12417 5065 12451
rect 4999 12401 5065 12417
rect 5107 12411 5173 12427
rect 5107 12377 5123 12411
rect 5157 12377 5173 12411
rect 5107 12361 5173 12377
rect 5245 12417 5341 12558
rect 5107 12359 5145 12361
rect 5027 12333 5145 12359
rect 5245 12325 5341 12408
rect 5245 12291 5295 12325
rect 5329 12291 5341 12325
rect 5245 12257 5341 12291
rect 5245 12223 5295 12257
rect 5329 12223 5341 12257
rect 5027 12197 5145 12223
rect 5245 12197 5341 12223
rect 5383 12660 5479 12699
rect 5671 12673 6617 12699
rect 6784 12673 6814 12699
rect 6870 12673 6900 12699
rect 6956 12673 6986 12699
rect 7042 12673 7072 12699
rect 7138 12673 7168 12699
rect 7419 12673 7629 12699
rect 7787 12673 8733 12699
rect 8900 12673 8930 12699
rect 8986 12673 9016 12699
rect 9072 12673 9102 12699
rect 9158 12673 9188 12699
rect 9254 12673 9284 12699
rect 9535 12673 9745 12699
rect 10004 12673 10034 12699
rect 10090 12673 10120 12699
rect 10176 12673 10206 12699
rect 10262 12673 10292 12699
rect 10358 12673 10388 12699
rect 10547 12673 10577 12699
rect 12107 12673 12137 12699
rect 12764 12673 12794 12699
rect 12850 12673 12880 12699
rect 12936 12673 12966 12699
rect 13022 12673 13052 12699
rect 13118 12673 13148 12699
rect 13308 12673 13338 12699
rect 13404 12673 13434 12699
rect 13490 12673 13520 12699
rect 13576 12673 13606 12699
rect 13662 12673 13692 12699
rect 13859 12673 13889 12699
rect 13947 12673 13977 12699
rect 14157 12673 14187 12699
rect 14241 12673 14341 12699
rect 14499 12673 14599 12699
rect 14664 12673 14694 12699
rect 5383 12626 5395 12660
rect 5429 12626 5479 12660
rect 5383 12592 5479 12626
rect 5383 12558 5395 12592
rect 5429 12558 5479 12592
rect 5383 12417 5479 12558
rect 5671 12473 6617 12499
rect 7419 12473 7629 12499
rect 7787 12473 8733 12499
rect 9535 12473 9745 12499
rect 10656 12634 10686 12660
rect 10759 12634 10789 12660
rect 10973 12634 11003 12660
rect 11045 12634 11075 12660
rect 11141 12634 11171 12660
rect 11513 12634 11543 12660
rect 11609 12634 11639 12660
rect 11681 12634 11711 12660
rect 11895 12634 11925 12660
rect 11998 12634 12028 12660
rect 6167 12451 6617 12473
rect 5383 12329 5479 12408
rect 5671 12415 6125 12431
rect 5671 12381 5947 12415
rect 5981 12381 6125 12415
rect 6167 12417 6311 12451
rect 6345 12417 6617 12451
rect 6167 12401 6617 12417
rect 6784 12435 6814 12473
rect 6870 12435 6900 12473
rect 6956 12435 6986 12473
rect 7042 12435 7072 12473
rect 7138 12441 7168 12473
rect 7545 12467 7629 12473
rect 7545 12451 7687 12467
rect 6784 12425 7072 12435
rect 6784 12413 6847 12425
rect 5671 12359 6125 12381
rect 6783 12391 6847 12413
rect 6881 12391 6915 12425
rect 6949 12391 6983 12425
rect 7017 12391 7072 12425
rect 6783 12386 7072 12391
rect 7119 12425 7179 12441
rect 7119 12391 7129 12425
rect 7163 12391 7179 12425
rect 6783 12380 7071 12386
rect 5671 12333 6617 12359
rect 5383 12295 5395 12329
rect 5429 12295 5479 12329
rect 5383 12261 5479 12295
rect 5383 12227 5395 12261
rect 5429 12227 5479 12261
rect 5383 12197 5479 12227
rect 6783 12307 6813 12380
rect 6869 12307 6899 12380
rect 6955 12307 6985 12380
rect 7041 12307 7071 12380
rect 7119 12375 7179 12391
rect 7361 12415 7503 12431
rect 7361 12381 7377 12415
rect 7411 12381 7503 12415
rect 7545 12417 7637 12451
rect 7671 12417 7687 12451
rect 8283 12451 8733 12473
rect 7545 12401 7687 12417
rect 7787 12415 8241 12431
rect 7138 12307 7168 12375
rect 7361 12365 7503 12381
rect 7419 12359 7503 12365
rect 7787 12381 8063 12415
rect 8097 12381 8241 12415
rect 8283 12417 8427 12451
rect 8461 12417 8733 12451
rect 8283 12401 8733 12417
rect 8900 12435 8930 12473
rect 8986 12435 9016 12473
rect 9072 12435 9102 12473
rect 9158 12435 9188 12473
rect 9254 12441 9284 12473
rect 9661 12467 9745 12473
rect 9661 12451 9803 12467
rect 8900 12425 9188 12435
rect 8900 12413 8963 12425
rect 7787 12359 8241 12381
rect 8899 12391 8963 12413
rect 8997 12391 9031 12425
rect 9065 12391 9099 12425
rect 9133 12391 9188 12425
rect 8899 12386 9188 12391
rect 9235 12425 9295 12441
rect 9235 12391 9245 12425
rect 9279 12391 9295 12425
rect 8899 12380 9187 12386
rect 7419 12333 7629 12359
rect 7787 12333 8733 12359
rect 8899 12307 8929 12380
rect 8985 12307 9015 12380
rect 9071 12307 9101 12380
rect 9157 12307 9187 12380
rect 9235 12375 9295 12391
rect 9477 12415 9619 12431
rect 9477 12381 9493 12415
rect 9527 12381 9619 12415
rect 9661 12417 9753 12451
rect 9787 12417 9803 12451
rect 9661 12401 9803 12417
rect 10004 12435 10034 12473
rect 10090 12435 10120 12473
rect 10176 12435 10206 12473
rect 10262 12435 10292 12473
rect 10358 12441 10388 12473
rect 10547 12441 10577 12473
rect 10656 12441 10686 12550
rect 10759 12535 10789 12550
rect 10759 12505 10907 12535
rect 10973 12518 11003 12550
rect 10004 12425 10292 12435
rect 10004 12413 10067 12425
rect 9254 12307 9284 12375
rect 9477 12365 9619 12381
rect 9535 12359 9619 12365
rect 10003 12391 10067 12413
rect 10101 12391 10135 12425
rect 10169 12391 10203 12425
rect 10237 12391 10292 12425
rect 10003 12386 10292 12391
rect 10339 12425 10399 12441
rect 10339 12391 10349 12425
rect 10383 12391 10399 12425
rect 10003 12380 10291 12386
rect 9535 12333 9745 12359
rect 10003 12307 10033 12380
rect 10089 12307 10119 12380
rect 10175 12307 10205 12380
rect 10261 12307 10291 12380
rect 10339 12375 10399 12391
rect 10544 12425 10598 12441
rect 10544 12391 10554 12425
rect 10588 12391 10598 12425
rect 10544 12375 10598 12391
rect 10640 12425 10694 12441
rect 10640 12391 10650 12425
rect 10684 12391 10694 12425
rect 10877 12405 10907 12505
rect 10949 12502 11003 12518
rect 10949 12468 10959 12502
rect 10993 12468 11003 12502
rect 10949 12452 11003 12468
rect 10640 12375 10694 12391
rect 10752 12389 10835 12405
rect 10358 12307 10388 12375
rect 10547 12353 10577 12375
rect 10656 12307 10686 12375
rect 10752 12355 10791 12389
rect 10825 12355 10835 12389
rect 10752 12339 10835 12355
rect 10877 12389 10931 12405
rect 11045 12399 11075 12550
rect 11141 12518 11171 12550
rect 11117 12502 11171 12518
rect 11117 12468 11127 12502
rect 11161 12468 11171 12502
rect 11117 12452 11171 12468
rect 10877 12355 10887 12389
rect 10921 12355 10931 12389
rect 11033 12389 11099 12399
rect 11033 12375 11049 12389
rect 10877 12339 10931 12355
rect 10973 12355 11049 12375
rect 11083 12355 11099 12389
rect 10973 12345 11099 12355
rect 10752 12307 10782 12339
rect 10877 12307 10907 12339
rect 10973 12307 11003 12345
rect 11141 12307 11171 12452
rect 11513 12518 11543 12550
rect 11513 12502 11567 12518
rect 11513 12468 11523 12502
rect 11557 12468 11567 12502
rect 11513 12452 11567 12468
rect 11513 12307 11543 12452
rect 11609 12399 11639 12550
rect 11681 12518 11711 12550
rect 11895 12535 11925 12550
rect 11681 12502 11735 12518
rect 11681 12468 11691 12502
rect 11725 12468 11735 12502
rect 11681 12452 11735 12468
rect 11777 12505 11925 12535
rect 11777 12405 11807 12505
rect 11998 12441 12028 12550
rect 13859 12500 13889 12515
rect 13853 12476 13889 12500
rect 12107 12441 12137 12473
rect 11990 12425 12044 12441
rect 11585 12389 11651 12399
rect 11585 12355 11601 12389
rect 11635 12375 11651 12389
rect 11753 12389 11807 12405
rect 11635 12355 11711 12375
rect 11585 12345 11711 12355
rect 11681 12307 11711 12345
rect 11753 12355 11763 12389
rect 11797 12355 11807 12389
rect 11753 12339 11807 12355
rect 11849 12389 11932 12405
rect 11849 12355 11859 12389
rect 11893 12355 11932 12389
rect 11990 12391 12000 12425
rect 12034 12391 12044 12425
rect 11990 12375 12044 12391
rect 12086 12425 12140 12441
rect 12086 12391 12096 12425
rect 12130 12391 12140 12425
rect 12764 12435 12794 12473
rect 12850 12435 12880 12473
rect 12936 12435 12966 12473
rect 13022 12435 13052 12473
rect 13118 12441 13148 12473
rect 13308 12441 13338 12473
rect 12764 12425 13052 12435
rect 12764 12413 12827 12425
rect 12086 12375 12140 12391
rect 12763 12391 12827 12413
rect 12861 12391 12895 12425
rect 12929 12391 12963 12425
rect 12997 12391 13052 12425
rect 12763 12386 13052 12391
rect 13099 12425 13159 12441
rect 13099 12391 13109 12425
rect 13143 12391 13159 12425
rect 12763 12380 13051 12386
rect 11849 12339 11932 12355
rect 11777 12307 11807 12339
rect 11902 12307 11932 12339
rect 11998 12307 12028 12375
rect 12107 12353 12137 12375
rect 12763 12307 12793 12380
rect 12849 12307 12879 12380
rect 12935 12307 12965 12380
rect 13021 12307 13051 12380
rect 13099 12375 13159 12391
rect 13297 12425 13357 12441
rect 13297 12391 13313 12425
rect 13347 12391 13357 12425
rect 13297 12375 13357 12391
rect 13404 12435 13434 12473
rect 13490 12435 13520 12473
rect 13576 12435 13606 12473
rect 13662 12435 13692 12473
rect 13853 12441 13883 12476
rect 13947 12454 13977 12515
rect 13404 12425 13692 12435
rect 13404 12391 13459 12425
rect 13493 12391 13527 12425
rect 13561 12391 13595 12425
rect 13629 12413 13692 12425
rect 13807 12425 13883 12441
rect 13629 12391 13693 12413
rect 13404 12386 13693 12391
rect 13405 12380 13693 12386
rect 13118 12307 13148 12375
rect 13308 12307 13338 12375
rect 13405 12307 13435 12380
rect 13491 12307 13521 12380
rect 13577 12307 13607 12380
rect 13663 12307 13693 12380
rect 13807 12391 13817 12425
rect 13851 12391 13883 12425
rect 13807 12375 13883 12391
rect 13927 12438 13981 12454
rect 14157 12441 14187 12589
rect 13927 12404 13937 12438
rect 13971 12404 13981 12438
rect 13927 12388 13981 12404
rect 14127 12425 14187 12441
rect 14127 12391 14137 12425
rect 14171 12391 14187 12425
rect 13853 12366 13883 12375
rect 13853 12342 13889 12366
rect 13859 12327 13889 12342
rect 13947 12327 13977 12388
rect 14127 12375 14187 12391
rect 14157 12307 14187 12375
rect 14241 12425 14341 12589
rect 14499 12441 14599 12589
rect 15147 12667 15177 12693
rect 15231 12667 15261 12693
rect 15498 12673 15528 12699
rect 15590 12673 15620 12699
rect 15689 12673 15719 12699
rect 15829 12673 15859 12699
rect 15926 12673 15956 12699
rect 16123 12673 16153 12699
rect 16222 12673 16252 12699
rect 16308 12673 16338 12699
rect 16392 12673 16422 12699
rect 16500 12673 16530 12699
rect 16584 12673 16614 12699
rect 16799 12673 16829 12699
rect 17080 12673 17110 12699
rect 17176 12673 17206 12699
rect 17262 12673 17292 12699
rect 17348 12673 17378 12699
rect 17434 12673 17464 12699
rect 17815 12673 18209 12699
rect 18367 12673 19313 12699
rect 19472 12673 19502 12699
rect 19568 12673 19598 12699
rect 19654 12673 19684 12699
rect 19740 12673 19770 12699
rect 19826 12673 19856 12699
rect 20023 12673 20141 12699
rect 15147 12524 15177 12539
rect 15114 12494 15177 12524
rect 14664 12441 14694 12473
rect 15114 12441 15144 12494
rect 15231 12450 15261 12539
rect 15498 12502 15528 12589
rect 15590 12551 15620 12589
rect 14241 12391 14251 12425
rect 14285 12391 14341 12425
rect 14241 12307 14341 12391
rect 14445 12425 14599 12441
rect 14445 12391 14455 12425
rect 14489 12391 14599 12425
rect 14445 12375 14599 12391
rect 14641 12425 14695 12441
rect 14641 12391 14651 12425
rect 14685 12391 14695 12425
rect 14641 12375 14695 12391
rect 15090 12425 15144 12441
rect 15090 12391 15100 12425
rect 15134 12391 15144 12425
rect 15186 12440 15261 12450
rect 15186 12406 15202 12440
rect 15236 12406 15261 12440
rect 15399 12486 15528 12502
rect 15574 12541 15640 12551
rect 15574 12507 15590 12541
rect 15624 12507 15640 12541
rect 15574 12497 15640 12507
rect 15399 12452 15409 12486
rect 15443 12472 15528 12486
rect 15443 12452 15516 12472
rect 15689 12455 15719 12589
rect 15829 12531 15859 12589
rect 15829 12515 15884 12531
rect 15829 12481 15839 12515
rect 15873 12481 15884 12515
rect 15829 12465 15884 12481
rect 15399 12436 15516 12452
rect 15186 12396 15261 12406
rect 15090 12375 15144 12391
rect 14499 12307 14599 12375
rect 14664 12353 14694 12375
rect 15114 12352 15144 12375
rect 15114 12322 15177 12352
rect 15147 12307 15177 12322
rect 15231 12307 15261 12396
rect 15486 12307 15516 12436
rect 15581 12425 15719 12455
rect 15581 12395 15612 12425
rect 15558 12379 15612 12395
rect 15558 12345 15568 12379
rect 15602 12345 15612 12379
rect 15558 12329 15612 12345
rect 15654 12373 15720 12383
rect 15654 12339 15670 12373
rect 15704 12339 15720 12373
rect 15654 12329 15720 12339
rect 15581 12295 15611 12329
rect 15677 12295 15707 12329
rect 15843 12307 15873 12465
rect 15926 12395 15956 12589
rect 16123 12490 16153 12505
rect 16047 12460 16153 12490
rect 16047 12443 16077 12460
rect 16011 12427 16077 12443
rect 15915 12379 15969 12395
rect 15915 12345 15925 12379
rect 15959 12345 15969 12379
rect 16011 12393 16021 12427
rect 16055 12393 16077 12427
rect 16222 12455 16252 12589
rect 16308 12557 16338 12589
rect 16294 12541 16348 12557
rect 16294 12507 16304 12541
rect 16338 12507 16348 12541
rect 16294 12491 16348 12507
rect 16222 12443 16272 12455
rect 16222 12431 16285 12443
rect 16222 12425 16309 12431
rect 16243 12415 16309 12425
rect 16243 12413 16265 12415
rect 16011 12377 16077 12393
rect 16047 12351 16077 12377
rect 16146 12367 16213 12383
rect 15915 12329 15969 12345
rect 15915 12307 15945 12329
rect 16146 12333 16169 12367
rect 16203 12333 16213 12367
rect 16146 12317 16213 12333
rect 16255 12381 16265 12413
rect 16299 12381 16309 12415
rect 16255 12365 16309 12381
rect 16392 12405 16422 12589
rect 16500 12433 16530 12589
rect 16584 12541 16614 12589
rect 16572 12525 16626 12541
rect 16572 12491 16582 12525
rect 16616 12491 16626 12525
rect 16572 12475 16626 12491
rect 16495 12417 16549 12433
rect 16392 12389 16453 12405
rect 16392 12369 16409 12389
rect 16146 12295 16176 12317
rect 16255 12295 16285 12365
rect 16351 12355 16409 12369
rect 16443 12355 16453 12389
rect 16495 12383 16505 12417
rect 16539 12383 16549 12417
rect 16495 12367 16549 12383
rect 16351 12339 16453 12355
rect 16351 12307 16381 12339
rect 16500 12307 16530 12367
rect 16591 12307 16621 12475
rect 17815 12473 18209 12499
rect 18367 12473 19313 12499
rect 16799 12441 16829 12473
rect 17080 12441 17110 12473
rect 16770 12425 16829 12441
rect 16770 12391 16780 12425
rect 16814 12391 16829 12425
rect 16770 12375 16829 12391
rect 17069 12425 17129 12441
rect 17069 12391 17085 12425
rect 17119 12391 17129 12425
rect 17069 12375 17129 12391
rect 17176 12435 17206 12473
rect 17262 12435 17292 12473
rect 17348 12435 17378 12473
rect 17434 12435 17464 12473
rect 17176 12425 17464 12435
rect 18033 12451 18209 12473
rect 17176 12391 17231 12425
rect 17265 12391 17299 12425
rect 17333 12391 17367 12425
rect 17401 12413 17464 12425
rect 17815 12415 17991 12431
rect 17401 12391 17465 12413
rect 17176 12386 17465 12391
rect 17177 12380 17465 12386
rect 16799 12353 16829 12375
rect 17080 12307 17110 12375
rect 17177 12307 17207 12380
rect 17263 12307 17293 12380
rect 17349 12307 17379 12380
rect 17435 12307 17465 12380
rect 17815 12381 17831 12415
rect 17865 12381 17941 12415
rect 17975 12381 17991 12415
rect 18033 12417 18049 12451
rect 18083 12417 18159 12451
rect 18193 12417 18209 12451
rect 18863 12451 19313 12473
rect 18033 12401 18209 12417
rect 18367 12415 18821 12431
rect 17815 12359 17991 12381
rect 18367 12381 18643 12415
rect 18677 12381 18821 12415
rect 18863 12417 19007 12451
rect 19041 12417 19313 12451
rect 19472 12441 19502 12473
rect 18863 12401 19313 12417
rect 19461 12425 19521 12441
rect 18367 12359 18821 12381
rect 19461 12391 19477 12425
rect 19511 12391 19521 12425
rect 19461 12375 19521 12391
rect 19568 12435 19598 12473
rect 19654 12435 19684 12473
rect 19740 12435 19770 12473
rect 19826 12435 19856 12473
rect 20023 12469 20141 12499
rect 19568 12425 19856 12435
rect 20103 12467 20141 12469
rect 20103 12451 20169 12467
rect 19568 12391 19623 12425
rect 19657 12391 19691 12425
rect 19725 12391 19759 12425
rect 19793 12413 19856 12425
rect 19793 12391 19857 12413
rect 19568 12386 19857 12391
rect 19569 12380 19857 12386
rect 17815 12333 18209 12359
rect 18367 12333 19313 12359
rect 19472 12307 19502 12375
rect 19569 12307 19599 12380
rect 19655 12307 19685 12380
rect 19741 12307 19771 12380
rect 19827 12307 19857 12380
rect 19995 12411 20061 12427
rect 19995 12377 20011 12411
rect 20045 12377 20061 12411
rect 20103 12417 20119 12451
rect 20153 12417 20169 12451
rect 20103 12401 20169 12417
rect 19995 12361 20061 12377
rect 20023 12359 20061 12361
rect 20023 12333 20141 12359
rect 5671 12197 6617 12223
rect 6783 12197 6813 12223
rect 6869 12197 6899 12223
rect 6955 12197 6985 12223
rect 7041 12197 7071 12223
rect 7138 12197 7168 12223
rect 7419 12197 7629 12223
rect 7787 12197 8733 12223
rect 8899 12197 8929 12223
rect 8985 12197 9015 12223
rect 9071 12197 9101 12223
rect 9157 12197 9187 12223
rect 9254 12197 9284 12223
rect 9535 12197 9745 12223
rect 10003 12197 10033 12223
rect 10089 12197 10119 12223
rect 10175 12197 10205 12223
rect 10261 12197 10291 12223
rect 10358 12197 10388 12223
rect 10547 12197 10577 12223
rect 10656 12197 10686 12223
rect 10752 12197 10782 12223
rect 10877 12197 10907 12223
rect 10973 12197 11003 12223
rect 11141 12197 11171 12223
rect 11513 12197 11543 12223
rect 11681 12197 11711 12223
rect 11777 12197 11807 12223
rect 11902 12197 11932 12223
rect 11998 12197 12028 12223
rect 12107 12197 12137 12223
rect 12763 12197 12793 12223
rect 12849 12197 12879 12223
rect 12935 12197 12965 12223
rect 13021 12197 13051 12223
rect 13118 12197 13148 12223
rect 13308 12197 13338 12223
rect 13405 12197 13435 12223
rect 13491 12197 13521 12223
rect 13577 12197 13607 12223
rect 13663 12197 13693 12223
rect 13859 12197 13889 12223
rect 13947 12197 13977 12223
rect 14157 12197 14187 12223
rect 14241 12197 14341 12223
rect 14499 12197 14599 12223
rect 14664 12197 14694 12223
rect 15147 12197 15177 12223
rect 15231 12197 15261 12223
rect 15486 12197 15516 12223
rect 15581 12197 15611 12223
rect 15677 12197 15707 12223
rect 15843 12197 15873 12223
rect 15915 12197 15945 12223
rect 16047 12197 16077 12223
rect 16146 12197 16176 12223
rect 16255 12197 16285 12223
rect 16351 12197 16381 12223
rect 16500 12197 16530 12223
rect 16591 12197 16621 12223
rect 16799 12197 16829 12223
rect 17080 12197 17110 12223
rect 17177 12197 17207 12223
rect 17263 12197 17293 12223
rect 17349 12197 17379 12223
rect 17435 12197 17465 12223
rect 17815 12197 18209 12223
rect 18367 12197 19313 12223
rect 19472 12197 19502 12223
rect 19569 12197 19599 12223
rect 19655 12197 19685 12223
rect 19741 12197 19771 12223
rect 19827 12197 19857 12223
rect 20023 12197 20141 12223
rect 29814 6831 30014 6847
rect 29814 6797 29830 6831
rect 29998 6797 30014 6831
rect 29814 6750 30014 6797
rect 30194 6831 30394 6847
rect 30194 6797 30210 6831
rect 30378 6797 30394 6831
rect 30194 6750 30394 6797
rect 30452 6831 30652 6847
rect 30452 6797 30468 6831
rect 30636 6797 30652 6831
rect 30452 6750 30652 6797
rect 30834 6831 31034 6847
rect 30834 6797 30850 6831
rect 31018 6797 31034 6831
rect 30834 6750 31034 6797
rect 31092 6831 31292 6847
rect 31092 6797 31108 6831
rect 31276 6797 31292 6831
rect 31092 6750 31292 6797
rect 31350 6831 31550 6847
rect 31350 6797 31366 6831
rect 31534 6797 31550 6831
rect 31350 6750 31550 6797
rect 31734 6831 31934 6847
rect 31734 6797 31750 6831
rect 31918 6797 31934 6831
rect 31734 6750 31934 6797
rect 31992 6831 32192 6847
rect 31992 6797 32008 6831
rect 32176 6797 32192 6831
rect 31992 6750 32192 6797
rect 32250 6831 32450 6847
rect 32250 6797 32266 6831
rect 32434 6797 32450 6831
rect 32250 6750 32450 6797
rect 32508 6831 32708 6847
rect 32508 6797 32524 6831
rect 32692 6797 32708 6831
rect 32508 6750 32708 6797
rect 32766 6831 32966 6847
rect 32766 6797 32782 6831
rect 32950 6797 32966 6831
rect 32766 6750 32966 6797
rect 33024 6831 33224 6847
rect 33024 6797 33040 6831
rect 33208 6797 33224 6831
rect 33024 6750 33224 6797
rect 33282 6831 33482 6847
rect 33282 6797 33298 6831
rect 33466 6797 33482 6831
rect 33282 6750 33482 6797
rect 33540 6831 33740 6847
rect 33540 6797 33556 6831
rect 33724 6797 33740 6831
rect 33540 6750 33740 6797
rect 33798 6831 33998 6847
rect 33798 6797 33814 6831
rect 33982 6797 33998 6831
rect 33798 6750 33998 6797
rect 34056 6831 34256 6847
rect 34056 6797 34072 6831
rect 34240 6797 34256 6831
rect 34056 6750 34256 6797
rect 34434 6831 34634 6847
rect 34434 6797 34450 6831
rect 34618 6797 34634 6831
rect 34434 6750 34634 6797
rect 29814 6103 30014 6150
rect 29814 6069 29830 6103
rect 29998 6069 30014 6103
rect 29814 6053 30014 6069
rect 30194 6103 30394 6150
rect 30194 6069 30210 6103
rect 30378 6069 30394 6103
rect 30194 6053 30394 6069
rect 30452 6103 30652 6150
rect 30452 6069 30468 6103
rect 30636 6069 30652 6103
rect 30452 6053 30652 6069
rect 30834 6103 31034 6150
rect 30834 6069 30850 6103
rect 31018 6069 31034 6103
rect 30834 6053 31034 6069
rect 31092 6103 31292 6150
rect 31092 6069 31108 6103
rect 31276 6069 31292 6103
rect 31092 6053 31292 6069
rect 31350 6103 31550 6150
rect 31350 6069 31366 6103
rect 31534 6069 31550 6103
rect 31350 6053 31550 6069
rect 31734 6103 31934 6150
rect 31734 6069 31750 6103
rect 31918 6069 31934 6103
rect 31734 6053 31934 6069
rect 31992 6103 32192 6150
rect 31992 6069 32008 6103
rect 32176 6069 32192 6103
rect 31992 6053 32192 6069
rect 32250 6103 32450 6150
rect 32250 6069 32266 6103
rect 32434 6069 32450 6103
rect 32250 6053 32450 6069
rect 32508 6103 32708 6150
rect 32508 6069 32524 6103
rect 32692 6069 32708 6103
rect 32508 6053 32708 6069
rect 32766 6103 32966 6150
rect 32766 6069 32782 6103
rect 32950 6069 32966 6103
rect 32766 6053 32966 6069
rect 33024 6103 33224 6150
rect 33024 6069 33040 6103
rect 33208 6069 33224 6103
rect 33024 6053 33224 6069
rect 33282 6103 33482 6150
rect 33282 6069 33298 6103
rect 33466 6069 33482 6103
rect 33282 6053 33482 6069
rect 33540 6103 33740 6150
rect 33540 6069 33556 6103
rect 33724 6069 33740 6103
rect 33540 6053 33740 6069
rect 33798 6103 33998 6150
rect 33798 6069 33814 6103
rect 33982 6069 33998 6103
rect 33798 6053 33998 6069
rect 34056 6103 34256 6150
rect 34056 6069 34072 6103
rect 34240 6069 34256 6103
rect 34056 6053 34256 6069
rect 34434 6103 34634 6150
rect 34434 6069 34450 6103
rect 34618 6069 34634 6103
rect 34434 6053 34634 6069
rect 30056 5811 30122 5827
rect 30056 5777 30072 5811
rect 30106 5777 30122 5811
rect 30056 5761 30122 5777
rect 30376 5811 30442 5827
rect 30376 5777 30392 5811
rect 30426 5777 30442 5811
rect 30376 5761 30442 5777
rect 30776 5811 30842 5827
rect 30776 5777 30792 5811
rect 30826 5777 30842 5811
rect 30776 5761 30842 5777
rect 31076 5811 31142 5827
rect 31076 5777 31092 5811
rect 31126 5777 31142 5811
rect 31076 5761 31142 5777
rect 30074 5730 30104 5761
rect 30298 5730 30328 5756
rect 30394 5730 30424 5761
rect 30490 5730 30520 5756
rect 30698 5730 30728 5756
rect 30794 5730 30824 5761
rect 30890 5730 30920 5756
rect 31094 5730 31124 5761
rect 30074 5099 30104 5130
rect 30298 5110 30328 5130
rect 30394 5110 30424 5130
rect 30490 5110 30520 5130
rect 30698 5110 30728 5130
rect 30794 5110 30824 5130
rect 30890 5110 30920 5130
rect 30290 5099 30520 5110
rect 30056 5083 30122 5099
rect 30056 5049 30072 5083
rect 30106 5049 30122 5083
rect 30056 5033 30122 5049
rect 30280 5083 30538 5099
rect 30280 5049 30296 5083
rect 30330 5049 30488 5083
rect 30522 5049 30538 5083
rect 30280 5040 30538 5049
rect 30280 5033 30346 5040
rect 30472 5033 30538 5040
rect 30680 5083 30940 5110
rect 31094 5099 31124 5130
rect 30680 5049 30696 5083
rect 30730 5050 30888 5083
rect 30730 5049 30746 5050
rect 30680 5033 30746 5049
rect 30872 5049 30888 5050
rect 30922 5050 30940 5083
rect 31076 5083 31142 5099
rect 30922 5049 30938 5050
rect 30872 5033 30938 5049
rect 31076 5049 31092 5083
rect 31126 5049 31142 5083
rect 31076 5033 31142 5049
rect 1466 4311 1532 4327
rect 1466 4277 1482 4311
rect 1516 4277 1532 4311
rect 1979 4310 2045 4320
rect 2171 4310 2237 4320
rect 2363 4310 2429 4320
rect 2555 4310 2621 4320
rect 2747 4310 2813 4320
rect 2939 4310 3005 4320
rect 1466 4261 1532 4277
rect 1900 4304 3005 4310
rect 1900 4270 1995 4304
rect 2029 4270 2187 4304
rect 2221 4270 2379 4304
rect 2413 4270 2571 4304
rect 2605 4270 2763 4304
rect 2797 4270 2955 4304
rect 2989 4270 3005 4304
rect 1484 4230 1514 4261
rect 1900 4260 3005 4270
rect 3166 4311 3232 4327
rect 3166 4277 3182 4311
rect 3216 4277 3232 4311
rect 3166 4261 3232 4277
rect 1900 4240 1934 4260
rect 1979 4254 2045 4260
rect 1901 4223 1931 4240
rect 1997 4223 2027 4254
rect 2093 4223 2123 4260
rect 2171 4254 2237 4260
rect 2189 4223 2219 4254
rect 2285 4223 2315 4260
rect 2363 4254 2429 4260
rect 2381 4223 2411 4254
rect 2477 4223 2507 4260
rect 2555 4254 2621 4260
rect 2573 4223 2603 4254
rect 2669 4223 2699 4260
rect 2747 4254 2813 4260
rect 2765 4223 2795 4254
rect 2861 4223 2891 4260
rect 2939 4254 3005 4260
rect 2957 4223 2987 4254
rect 3184 4230 3214 4261
rect 1666 3911 1732 3927
rect 1666 3877 1682 3911
rect 1716 3877 1732 3911
rect 1666 3861 1732 3877
rect 1684 3830 1714 3861
rect 1484 3199 1514 3230
rect 1684 3199 1714 3230
rect 1466 3183 1532 3199
rect 1466 3149 1482 3183
rect 1516 3149 1532 3183
rect 1466 3133 1532 3149
rect 1666 3183 1732 3199
rect 1901 3192 1931 3223
rect 1997 3197 2027 3223
rect 2093 3192 2123 3223
rect 2189 3197 2219 3223
rect 2285 3192 2315 3223
rect 2381 3197 2411 3223
rect 2477 3192 2507 3223
rect 2573 3197 2603 3223
rect 2669 3192 2699 3223
rect 2765 3197 2795 3223
rect 2861 3192 2891 3223
rect 2957 3197 2987 3223
rect 3184 3199 3214 3230
rect 1666 3149 1682 3183
rect 1716 3149 1732 3183
rect 1666 3133 1732 3149
rect 1883 3176 1949 3192
rect 1883 3142 1899 3176
rect 1933 3142 1949 3176
rect 1883 3126 1949 3142
rect 2075 3176 2141 3192
rect 2075 3142 2091 3176
rect 2125 3142 2141 3176
rect 2075 3126 2141 3142
rect 2267 3176 2333 3192
rect 2267 3142 2283 3176
rect 2317 3142 2333 3176
rect 2267 3126 2333 3142
rect 2459 3176 2525 3192
rect 2459 3142 2475 3176
rect 2509 3142 2525 3176
rect 2459 3126 2525 3142
rect 2651 3176 2717 3192
rect 2651 3142 2667 3176
rect 2701 3142 2717 3176
rect 2651 3126 2717 3142
rect 2843 3176 2909 3192
rect 2843 3142 2859 3176
rect 2893 3142 2909 3176
rect 2843 3126 2909 3142
rect 3166 3183 3232 3199
rect 3166 3149 3182 3183
rect 3216 3149 3232 3183
rect 3166 3133 3232 3149
rect 4766 4311 4832 4327
rect 4766 4277 4782 4311
rect 4816 4277 4832 4311
rect 5279 4310 5345 4320
rect 5471 4310 5537 4320
rect 5663 4310 5729 4320
rect 5855 4310 5921 4320
rect 6047 4310 6113 4320
rect 6239 4310 6305 4320
rect 4766 4261 4832 4277
rect 5200 4304 6305 4310
rect 5200 4270 5295 4304
rect 5329 4270 5487 4304
rect 5521 4270 5679 4304
rect 5713 4270 5871 4304
rect 5905 4270 6063 4304
rect 6097 4270 6255 4304
rect 6289 4270 6305 4304
rect 4784 4230 4814 4261
rect 5200 4260 6305 4270
rect 6466 4311 6532 4327
rect 6466 4277 6482 4311
rect 6516 4277 6532 4311
rect 6466 4261 6532 4277
rect 5200 4240 5234 4260
rect 5279 4254 5345 4260
rect 5201 4223 5231 4240
rect 5297 4223 5327 4254
rect 5393 4223 5423 4260
rect 5471 4254 5537 4260
rect 5489 4223 5519 4254
rect 5585 4223 5615 4260
rect 5663 4254 5729 4260
rect 5681 4223 5711 4254
rect 5777 4223 5807 4260
rect 5855 4254 5921 4260
rect 5873 4223 5903 4254
rect 5969 4223 5999 4260
rect 6047 4254 6113 4260
rect 6065 4223 6095 4254
rect 6161 4223 6191 4260
rect 6239 4254 6305 4260
rect 6257 4223 6287 4254
rect 6484 4230 6514 4261
rect 4966 3911 5032 3927
rect 4966 3877 4982 3911
rect 5016 3877 5032 3911
rect 4966 3861 5032 3877
rect 4984 3830 5014 3861
rect 4784 3199 4814 3230
rect 4984 3199 5014 3230
rect 4766 3183 4832 3199
rect 4766 3149 4782 3183
rect 4816 3149 4832 3183
rect 4766 3133 4832 3149
rect 4966 3183 5032 3199
rect 5201 3192 5231 3223
rect 5297 3197 5327 3223
rect 5393 3192 5423 3223
rect 5489 3197 5519 3223
rect 5585 3192 5615 3223
rect 5681 3197 5711 3223
rect 5777 3192 5807 3223
rect 5873 3197 5903 3223
rect 5969 3192 5999 3223
rect 6065 3197 6095 3223
rect 6161 3192 6191 3223
rect 6257 3197 6287 3223
rect 6484 3199 6514 3230
rect 4966 3149 4982 3183
rect 5016 3149 5032 3183
rect 4966 3133 5032 3149
rect 5183 3176 5249 3192
rect 5183 3142 5199 3176
rect 5233 3142 5249 3176
rect 5183 3126 5249 3142
rect 5375 3176 5441 3192
rect 5375 3142 5391 3176
rect 5425 3142 5441 3176
rect 5375 3126 5441 3142
rect 5567 3176 5633 3192
rect 5567 3142 5583 3176
rect 5617 3142 5633 3176
rect 5567 3126 5633 3142
rect 5759 3176 5825 3192
rect 5759 3142 5775 3176
rect 5809 3142 5825 3176
rect 5759 3126 5825 3142
rect 5951 3176 6017 3192
rect 5951 3142 5967 3176
rect 6001 3142 6017 3176
rect 5951 3126 6017 3142
rect 6143 3176 6209 3192
rect 6143 3142 6159 3176
rect 6193 3142 6209 3176
rect 6143 3126 6209 3142
rect 6466 3183 6532 3199
rect 6466 3149 6482 3183
rect 6516 3149 6532 3183
rect 6466 3133 6532 3149
rect 8066 4311 8132 4327
rect 8066 4277 8082 4311
rect 8116 4277 8132 4311
rect 8579 4310 8645 4320
rect 8771 4310 8837 4320
rect 8963 4310 9029 4320
rect 9155 4310 9221 4320
rect 9347 4310 9413 4320
rect 9539 4310 9605 4320
rect 8066 4261 8132 4277
rect 8500 4304 9605 4310
rect 8500 4270 8595 4304
rect 8629 4270 8787 4304
rect 8821 4270 8979 4304
rect 9013 4270 9171 4304
rect 9205 4270 9363 4304
rect 9397 4270 9555 4304
rect 9589 4270 9605 4304
rect 8084 4230 8114 4261
rect 8500 4260 9605 4270
rect 9766 4311 9832 4327
rect 9766 4277 9782 4311
rect 9816 4277 9832 4311
rect 9766 4261 9832 4277
rect 8500 4240 8534 4260
rect 8579 4254 8645 4260
rect 8501 4223 8531 4240
rect 8597 4223 8627 4254
rect 8693 4223 8723 4260
rect 8771 4254 8837 4260
rect 8789 4223 8819 4254
rect 8885 4223 8915 4260
rect 8963 4254 9029 4260
rect 8981 4223 9011 4254
rect 9077 4223 9107 4260
rect 9155 4254 9221 4260
rect 9173 4223 9203 4254
rect 9269 4223 9299 4260
rect 9347 4254 9413 4260
rect 9365 4223 9395 4254
rect 9461 4223 9491 4260
rect 9539 4254 9605 4260
rect 9557 4223 9587 4254
rect 9784 4230 9814 4261
rect 8266 3911 8332 3927
rect 8266 3877 8282 3911
rect 8316 3877 8332 3911
rect 8266 3861 8332 3877
rect 8284 3830 8314 3861
rect 8084 3199 8114 3230
rect 8284 3199 8314 3230
rect 8066 3183 8132 3199
rect 8066 3149 8082 3183
rect 8116 3149 8132 3183
rect 8066 3133 8132 3149
rect 8266 3183 8332 3199
rect 8501 3192 8531 3223
rect 8597 3197 8627 3223
rect 8693 3192 8723 3223
rect 8789 3197 8819 3223
rect 8885 3192 8915 3223
rect 8981 3197 9011 3223
rect 9077 3192 9107 3223
rect 9173 3197 9203 3223
rect 9269 3192 9299 3223
rect 9365 3197 9395 3223
rect 9461 3192 9491 3223
rect 9557 3197 9587 3223
rect 9784 3199 9814 3230
rect 8266 3149 8282 3183
rect 8316 3149 8332 3183
rect 8266 3133 8332 3149
rect 8483 3176 8549 3192
rect 8483 3142 8499 3176
rect 8533 3142 8549 3176
rect 8483 3126 8549 3142
rect 8675 3176 8741 3192
rect 8675 3142 8691 3176
rect 8725 3142 8741 3176
rect 8675 3126 8741 3142
rect 8867 3176 8933 3192
rect 8867 3142 8883 3176
rect 8917 3142 8933 3176
rect 8867 3126 8933 3142
rect 9059 3176 9125 3192
rect 9059 3142 9075 3176
rect 9109 3142 9125 3176
rect 9059 3126 9125 3142
rect 9251 3176 9317 3192
rect 9251 3142 9267 3176
rect 9301 3142 9317 3176
rect 9251 3126 9317 3142
rect 9443 3176 9509 3192
rect 9443 3142 9459 3176
rect 9493 3142 9509 3176
rect 9443 3126 9509 3142
rect 9766 3183 9832 3199
rect 9766 3149 9782 3183
rect 9816 3149 9832 3183
rect 9766 3133 9832 3149
rect 11366 4311 11432 4327
rect 11366 4277 11382 4311
rect 11416 4277 11432 4311
rect 11879 4310 11945 4320
rect 12071 4310 12137 4320
rect 12263 4310 12329 4320
rect 12455 4310 12521 4320
rect 12647 4310 12713 4320
rect 12839 4310 12905 4320
rect 11366 4261 11432 4277
rect 11800 4304 12905 4310
rect 11800 4270 11895 4304
rect 11929 4270 12087 4304
rect 12121 4270 12279 4304
rect 12313 4270 12471 4304
rect 12505 4270 12663 4304
rect 12697 4270 12855 4304
rect 12889 4270 12905 4304
rect 11384 4230 11414 4261
rect 11800 4260 12905 4270
rect 13066 4311 13132 4327
rect 13066 4277 13082 4311
rect 13116 4277 13132 4311
rect 13066 4261 13132 4277
rect 11800 4240 11834 4260
rect 11879 4254 11945 4260
rect 11801 4223 11831 4240
rect 11897 4223 11927 4254
rect 11993 4223 12023 4260
rect 12071 4254 12137 4260
rect 12089 4223 12119 4254
rect 12185 4223 12215 4260
rect 12263 4254 12329 4260
rect 12281 4223 12311 4254
rect 12377 4223 12407 4260
rect 12455 4254 12521 4260
rect 12473 4223 12503 4254
rect 12569 4223 12599 4260
rect 12647 4254 12713 4260
rect 12665 4223 12695 4254
rect 12761 4223 12791 4260
rect 12839 4254 12905 4260
rect 12857 4223 12887 4254
rect 13084 4230 13114 4261
rect 11566 3911 11632 3927
rect 11566 3877 11582 3911
rect 11616 3877 11632 3911
rect 11566 3861 11632 3877
rect 11584 3830 11614 3861
rect 11384 3199 11414 3230
rect 11584 3199 11614 3230
rect 11366 3183 11432 3199
rect 11366 3149 11382 3183
rect 11416 3149 11432 3183
rect 11366 3133 11432 3149
rect 11566 3183 11632 3199
rect 11801 3192 11831 3223
rect 11897 3197 11927 3223
rect 11993 3192 12023 3223
rect 12089 3197 12119 3223
rect 12185 3192 12215 3223
rect 12281 3197 12311 3223
rect 12377 3192 12407 3223
rect 12473 3197 12503 3223
rect 12569 3192 12599 3223
rect 12665 3197 12695 3223
rect 12761 3192 12791 3223
rect 12857 3197 12887 3223
rect 13084 3199 13114 3230
rect 11566 3149 11582 3183
rect 11616 3149 11632 3183
rect 11566 3133 11632 3149
rect 11783 3176 11849 3192
rect 11783 3142 11799 3176
rect 11833 3142 11849 3176
rect 11783 3126 11849 3142
rect 11975 3176 12041 3192
rect 11975 3142 11991 3176
rect 12025 3142 12041 3176
rect 11975 3126 12041 3142
rect 12167 3176 12233 3192
rect 12167 3142 12183 3176
rect 12217 3142 12233 3176
rect 12167 3126 12233 3142
rect 12359 3176 12425 3192
rect 12359 3142 12375 3176
rect 12409 3142 12425 3176
rect 12359 3126 12425 3142
rect 12551 3176 12617 3192
rect 12551 3142 12567 3176
rect 12601 3142 12617 3176
rect 12551 3126 12617 3142
rect 12743 3176 12809 3192
rect 12743 3142 12759 3176
rect 12793 3142 12809 3176
rect 12743 3126 12809 3142
rect 13066 3183 13132 3199
rect 13066 3149 13082 3183
rect 13116 3149 13132 3183
rect 13066 3133 13132 3149
rect 14966 4311 15032 4327
rect 14966 4277 14982 4311
rect 15016 4277 15032 4311
rect 15479 4310 15545 4320
rect 15671 4310 15737 4320
rect 15863 4310 15929 4320
rect 16055 4310 16121 4320
rect 16247 4310 16313 4320
rect 16439 4310 16505 4320
rect 14966 4261 15032 4277
rect 15400 4304 16505 4310
rect 15400 4270 15495 4304
rect 15529 4270 15687 4304
rect 15721 4270 15879 4304
rect 15913 4270 16071 4304
rect 16105 4270 16263 4304
rect 16297 4270 16455 4304
rect 16489 4270 16505 4304
rect 14984 4230 15014 4261
rect 15400 4260 16505 4270
rect 16666 4311 16732 4327
rect 16666 4277 16682 4311
rect 16716 4277 16732 4311
rect 16666 4261 16732 4277
rect 15400 4240 15434 4260
rect 15479 4254 15545 4260
rect 15401 4223 15431 4240
rect 15497 4223 15527 4254
rect 15593 4223 15623 4260
rect 15671 4254 15737 4260
rect 15689 4223 15719 4254
rect 15785 4223 15815 4260
rect 15863 4254 15929 4260
rect 15881 4223 15911 4254
rect 15977 4223 16007 4260
rect 16055 4254 16121 4260
rect 16073 4223 16103 4254
rect 16169 4223 16199 4260
rect 16247 4254 16313 4260
rect 16265 4223 16295 4254
rect 16361 4223 16391 4260
rect 16439 4254 16505 4260
rect 16457 4223 16487 4254
rect 16684 4230 16714 4261
rect 15166 3911 15232 3927
rect 15166 3877 15182 3911
rect 15216 3877 15232 3911
rect 15166 3861 15232 3877
rect 15184 3830 15214 3861
rect 14984 3199 15014 3230
rect 15184 3199 15214 3230
rect 14966 3183 15032 3199
rect 14966 3149 14982 3183
rect 15016 3149 15032 3183
rect 14966 3133 15032 3149
rect 15166 3183 15232 3199
rect 15401 3192 15431 3223
rect 15497 3197 15527 3223
rect 15593 3192 15623 3223
rect 15689 3197 15719 3223
rect 15785 3192 15815 3223
rect 15881 3197 15911 3223
rect 15977 3192 16007 3223
rect 16073 3197 16103 3223
rect 16169 3192 16199 3223
rect 16265 3197 16295 3223
rect 16361 3192 16391 3223
rect 16457 3197 16487 3223
rect 16684 3199 16714 3230
rect 15166 3149 15182 3183
rect 15216 3149 15232 3183
rect 15166 3133 15232 3149
rect 15383 3176 15449 3192
rect 15383 3142 15399 3176
rect 15433 3142 15449 3176
rect 15383 3126 15449 3142
rect 15575 3176 15641 3192
rect 15575 3142 15591 3176
rect 15625 3142 15641 3176
rect 15575 3126 15641 3142
rect 15767 3176 15833 3192
rect 15767 3142 15783 3176
rect 15817 3142 15833 3176
rect 15767 3126 15833 3142
rect 15959 3176 16025 3192
rect 15959 3142 15975 3176
rect 16009 3142 16025 3176
rect 15959 3126 16025 3142
rect 16151 3176 16217 3192
rect 16151 3142 16167 3176
rect 16201 3142 16217 3176
rect 16151 3126 16217 3142
rect 16343 3176 16409 3192
rect 16343 3142 16359 3176
rect 16393 3142 16409 3176
rect 16343 3126 16409 3142
rect 16666 3183 16732 3199
rect 16666 3149 16682 3183
rect 16716 3149 16732 3183
rect 16666 3133 16732 3149
rect 18466 4311 18532 4327
rect 18466 4277 18482 4311
rect 18516 4277 18532 4311
rect 18979 4310 19045 4320
rect 19171 4310 19237 4320
rect 19363 4310 19429 4320
rect 19555 4310 19621 4320
rect 19747 4310 19813 4320
rect 19939 4310 20005 4320
rect 18466 4261 18532 4277
rect 18900 4304 20005 4310
rect 18900 4270 18995 4304
rect 19029 4270 19187 4304
rect 19221 4270 19379 4304
rect 19413 4270 19571 4304
rect 19605 4270 19763 4304
rect 19797 4270 19955 4304
rect 19989 4270 20005 4304
rect 18484 4230 18514 4261
rect 18900 4260 20005 4270
rect 20166 4311 20232 4327
rect 20166 4277 20182 4311
rect 20216 4277 20232 4311
rect 20166 4261 20232 4277
rect 18900 4240 18934 4260
rect 18979 4254 19045 4260
rect 18901 4223 18931 4240
rect 18997 4223 19027 4254
rect 19093 4223 19123 4260
rect 19171 4254 19237 4260
rect 19189 4223 19219 4254
rect 19285 4223 19315 4260
rect 19363 4254 19429 4260
rect 19381 4223 19411 4254
rect 19477 4223 19507 4260
rect 19555 4254 19621 4260
rect 19573 4223 19603 4254
rect 19669 4223 19699 4260
rect 19747 4254 19813 4260
rect 19765 4223 19795 4254
rect 19861 4223 19891 4260
rect 19939 4254 20005 4260
rect 19957 4223 19987 4254
rect 20184 4230 20214 4261
rect 18666 3911 18732 3927
rect 18666 3877 18682 3911
rect 18716 3877 18732 3911
rect 18666 3861 18732 3877
rect 18684 3830 18714 3861
rect 18484 3199 18514 3230
rect 18684 3199 18714 3230
rect 18466 3183 18532 3199
rect 18466 3149 18482 3183
rect 18516 3149 18532 3183
rect 18466 3133 18532 3149
rect 18666 3183 18732 3199
rect 18901 3192 18931 3223
rect 18997 3197 19027 3223
rect 19093 3192 19123 3223
rect 19189 3197 19219 3223
rect 19285 3192 19315 3223
rect 19381 3197 19411 3223
rect 19477 3192 19507 3223
rect 19573 3197 19603 3223
rect 19669 3192 19699 3223
rect 19765 3197 19795 3223
rect 19861 3192 19891 3223
rect 19957 3197 19987 3223
rect 20184 3199 20214 3230
rect 18666 3149 18682 3183
rect 18716 3149 18732 3183
rect 18666 3133 18732 3149
rect 18883 3176 18949 3192
rect 18883 3142 18899 3176
rect 18933 3142 18949 3176
rect 18883 3126 18949 3142
rect 19075 3176 19141 3192
rect 19075 3142 19091 3176
rect 19125 3142 19141 3176
rect 19075 3126 19141 3142
rect 19267 3176 19333 3192
rect 19267 3142 19283 3176
rect 19317 3142 19333 3176
rect 19267 3126 19333 3142
rect 19459 3176 19525 3192
rect 19459 3142 19475 3176
rect 19509 3142 19525 3176
rect 19459 3126 19525 3142
rect 19651 3176 19717 3192
rect 19651 3142 19667 3176
rect 19701 3142 19717 3176
rect 19651 3126 19717 3142
rect 19843 3176 19909 3192
rect 19843 3142 19859 3176
rect 19893 3142 19909 3176
rect 19843 3126 19909 3142
rect 20166 3183 20232 3199
rect 20166 3149 20182 3183
rect 20216 3149 20232 3183
rect 20166 3133 20232 3149
rect 22166 4311 22232 4327
rect 22166 4277 22182 4311
rect 22216 4277 22232 4311
rect 22679 4310 22745 4320
rect 22871 4310 22937 4320
rect 23063 4310 23129 4320
rect 23255 4310 23321 4320
rect 23447 4310 23513 4320
rect 23639 4310 23705 4320
rect 22166 4261 22232 4277
rect 22600 4304 23705 4310
rect 22600 4270 22695 4304
rect 22729 4270 22887 4304
rect 22921 4270 23079 4304
rect 23113 4270 23271 4304
rect 23305 4270 23463 4304
rect 23497 4270 23655 4304
rect 23689 4270 23705 4304
rect 22184 4230 22214 4261
rect 22600 4260 23705 4270
rect 23866 4311 23932 4327
rect 23866 4277 23882 4311
rect 23916 4277 23932 4311
rect 23866 4261 23932 4277
rect 22600 4240 22634 4260
rect 22679 4254 22745 4260
rect 22601 4223 22631 4240
rect 22697 4223 22727 4254
rect 22793 4223 22823 4260
rect 22871 4254 22937 4260
rect 22889 4223 22919 4254
rect 22985 4223 23015 4260
rect 23063 4254 23129 4260
rect 23081 4223 23111 4254
rect 23177 4223 23207 4260
rect 23255 4254 23321 4260
rect 23273 4223 23303 4254
rect 23369 4223 23399 4260
rect 23447 4254 23513 4260
rect 23465 4223 23495 4254
rect 23561 4223 23591 4260
rect 23639 4254 23705 4260
rect 23657 4223 23687 4254
rect 23884 4230 23914 4261
rect 22366 3911 22432 3927
rect 22366 3877 22382 3911
rect 22416 3877 22432 3911
rect 22366 3861 22432 3877
rect 22384 3830 22414 3861
rect 22184 3199 22214 3230
rect 22384 3199 22414 3230
rect 22166 3183 22232 3199
rect 22166 3149 22182 3183
rect 22216 3149 22232 3183
rect 22166 3133 22232 3149
rect 22366 3183 22432 3199
rect 22601 3192 22631 3223
rect 22697 3197 22727 3223
rect 22793 3192 22823 3223
rect 22889 3197 22919 3223
rect 22985 3192 23015 3223
rect 23081 3197 23111 3223
rect 23177 3192 23207 3223
rect 23273 3197 23303 3223
rect 23369 3192 23399 3223
rect 23465 3197 23495 3223
rect 23561 3192 23591 3223
rect 23657 3197 23687 3223
rect 23884 3199 23914 3230
rect 22366 3149 22382 3183
rect 22416 3149 22432 3183
rect 22366 3133 22432 3149
rect 22583 3176 22649 3192
rect 22583 3142 22599 3176
rect 22633 3142 22649 3176
rect 22583 3126 22649 3142
rect 22775 3176 22841 3192
rect 22775 3142 22791 3176
rect 22825 3142 22841 3176
rect 22775 3126 22841 3142
rect 22967 3176 23033 3192
rect 22967 3142 22983 3176
rect 23017 3142 23033 3176
rect 22967 3126 23033 3142
rect 23159 3176 23225 3192
rect 23159 3142 23175 3176
rect 23209 3142 23225 3176
rect 23159 3126 23225 3142
rect 23351 3176 23417 3192
rect 23351 3142 23367 3176
rect 23401 3142 23417 3176
rect 23351 3126 23417 3142
rect 23543 3176 23609 3192
rect 23543 3142 23559 3176
rect 23593 3142 23609 3176
rect 23543 3126 23609 3142
rect 23866 3183 23932 3199
rect 23866 3149 23882 3183
rect 23916 3149 23932 3183
rect 23866 3133 23932 3149
rect 25966 4311 26032 4327
rect 25966 4277 25982 4311
rect 26016 4277 26032 4311
rect 26479 4310 26545 4320
rect 26671 4310 26737 4320
rect 26863 4310 26929 4320
rect 27055 4310 27121 4320
rect 27247 4310 27313 4320
rect 27439 4310 27505 4320
rect 25966 4261 26032 4277
rect 26400 4304 27505 4310
rect 26400 4270 26495 4304
rect 26529 4270 26687 4304
rect 26721 4270 26879 4304
rect 26913 4270 27071 4304
rect 27105 4270 27263 4304
rect 27297 4270 27455 4304
rect 27489 4270 27505 4304
rect 25984 4230 26014 4261
rect 26400 4260 27505 4270
rect 27666 4311 27732 4327
rect 27666 4277 27682 4311
rect 27716 4277 27732 4311
rect 27666 4261 27732 4277
rect 26400 4240 26434 4260
rect 26479 4254 26545 4260
rect 26401 4223 26431 4240
rect 26497 4223 26527 4254
rect 26593 4223 26623 4260
rect 26671 4254 26737 4260
rect 26689 4223 26719 4254
rect 26785 4223 26815 4260
rect 26863 4254 26929 4260
rect 26881 4223 26911 4254
rect 26977 4223 27007 4260
rect 27055 4254 27121 4260
rect 27073 4223 27103 4254
rect 27169 4223 27199 4260
rect 27247 4254 27313 4260
rect 27265 4223 27295 4254
rect 27361 4223 27391 4260
rect 27439 4254 27505 4260
rect 27457 4223 27487 4254
rect 27684 4230 27714 4261
rect 26166 3911 26232 3927
rect 26166 3877 26182 3911
rect 26216 3877 26232 3911
rect 26166 3861 26232 3877
rect 26184 3830 26214 3861
rect 25984 3199 26014 3230
rect 26184 3199 26214 3230
rect 25966 3183 26032 3199
rect 25966 3149 25982 3183
rect 26016 3149 26032 3183
rect 25966 3133 26032 3149
rect 26166 3183 26232 3199
rect 26401 3192 26431 3223
rect 26497 3197 26527 3223
rect 26593 3192 26623 3223
rect 26689 3197 26719 3223
rect 26785 3192 26815 3223
rect 26881 3197 26911 3223
rect 26977 3192 27007 3223
rect 27073 3197 27103 3223
rect 27169 3192 27199 3223
rect 27265 3197 27295 3223
rect 27361 3192 27391 3223
rect 27457 3197 27487 3223
rect 27684 3199 27714 3230
rect 26166 3149 26182 3183
rect 26216 3149 26232 3183
rect 26166 3133 26232 3149
rect 26383 3176 26449 3192
rect 26383 3142 26399 3176
rect 26433 3142 26449 3176
rect 26383 3126 26449 3142
rect 26575 3176 26641 3192
rect 26575 3142 26591 3176
rect 26625 3142 26641 3176
rect 26575 3126 26641 3142
rect 26767 3176 26833 3192
rect 26767 3142 26783 3176
rect 26817 3142 26833 3176
rect 26767 3126 26833 3142
rect 26959 3176 27025 3192
rect 26959 3142 26975 3176
rect 27009 3142 27025 3176
rect 26959 3126 27025 3142
rect 27151 3176 27217 3192
rect 27151 3142 27167 3176
rect 27201 3142 27217 3176
rect 27151 3126 27217 3142
rect 27343 3176 27409 3192
rect 27343 3142 27359 3176
rect 27393 3142 27409 3176
rect 27343 3126 27409 3142
rect 27666 3183 27732 3199
rect 27666 3149 27682 3183
rect 27716 3149 27732 3183
rect 27666 3133 27732 3149
rect 29918 4630 30118 4646
rect 29918 4596 29934 4630
rect 30102 4596 30118 4630
rect 29918 4558 30118 4596
rect 30298 4630 30498 4646
rect 30298 4596 30314 4630
rect 30482 4596 30498 4630
rect 30298 4558 30498 4596
rect 30698 4630 30898 4646
rect 30698 4596 30714 4630
rect 30882 4596 30898 4630
rect 30698 4558 30898 4596
rect 31078 4630 31278 4646
rect 31078 4596 31094 4630
rect 31262 4596 31278 4630
rect 31078 4558 31278 4596
rect 31336 4630 31536 4646
rect 31336 4596 31352 4630
rect 31520 4596 31536 4630
rect 31336 4558 31536 4596
rect 31594 4630 31794 4646
rect 31594 4596 31610 4630
rect 31778 4596 31794 4630
rect 31594 4558 31794 4596
rect 31852 4630 32052 4646
rect 31852 4596 31868 4630
rect 32036 4596 32052 4630
rect 31852 4558 32052 4596
rect 32110 4630 32310 4646
rect 32110 4596 32126 4630
rect 32294 4596 32310 4630
rect 32110 4558 32310 4596
rect 32368 4630 32568 4646
rect 32368 4596 32384 4630
rect 32552 4596 32568 4630
rect 32368 4558 32568 4596
rect 32626 4630 32826 4646
rect 32626 4596 32642 4630
rect 32810 4596 32826 4630
rect 32626 4558 32826 4596
rect 32884 4630 33084 4646
rect 32884 4596 32900 4630
rect 33068 4596 33084 4630
rect 32884 4558 33084 4596
rect 33142 4630 33342 4646
rect 33142 4596 33158 4630
rect 33326 4596 33342 4630
rect 33142 4558 33342 4596
rect 33518 4630 33718 4646
rect 33518 4596 33534 4630
rect 33702 4596 33718 4630
rect 33518 4558 33718 4596
rect 29918 4320 30118 4358
rect 29918 4286 29934 4320
rect 30102 4286 30118 4320
rect 29918 4270 30118 4286
rect 30298 4320 30498 4358
rect 30298 4286 30314 4320
rect 30482 4286 30498 4320
rect 30298 4270 30498 4286
rect 30698 4320 30898 4358
rect 30698 4286 30714 4320
rect 30882 4286 30898 4320
rect 30698 4270 30898 4286
rect 31078 4320 31278 4358
rect 31078 4286 31094 4320
rect 31262 4286 31278 4320
rect 31078 4270 31278 4286
rect 31336 4320 31536 4358
rect 31336 4286 31352 4320
rect 31520 4286 31536 4320
rect 31336 4270 31536 4286
rect 31594 4320 31794 4358
rect 31594 4286 31610 4320
rect 31778 4286 31794 4320
rect 31594 4270 31794 4286
rect 31852 4320 32052 4358
rect 31852 4286 31868 4320
rect 32036 4286 32052 4320
rect 31852 4270 32052 4286
rect 32110 4320 32310 4358
rect 32110 4286 32126 4320
rect 32294 4286 32310 4320
rect 32110 4270 32310 4286
rect 32368 4320 32568 4358
rect 32368 4286 32384 4320
rect 32552 4286 32568 4320
rect 32368 4270 32568 4286
rect 32626 4320 32826 4358
rect 32626 4286 32642 4320
rect 32810 4286 32826 4320
rect 32626 4270 32826 4286
rect 32884 4320 33084 4358
rect 32884 4286 32900 4320
rect 33068 4286 33084 4320
rect 32884 4270 33084 4286
rect 33142 4320 33342 4358
rect 33142 4286 33158 4320
rect 33326 4286 33342 4320
rect 33142 4270 33342 4286
rect 33518 4320 33718 4358
rect 33518 4286 33534 4320
rect 33702 4286 33718 4320
rect 33518 4270 33718 4286
rect 1470 2780 1536 2796
rect 1470 2746 1486 2780
rect 1520 2746 1536 2780
rect 1470 2730 1536 2746
rect 1670 2780 1736 2796
rect 1670 2746 1686 2780
rect 1720 2746 1736 2780
rect 1670 2730 1736 2746
rect 1983 2773 2049 2789
rect 1983 2739 1999 2773
rect 2033 2739 2049 2773
rect 1488 2708 1518 2730
rect 1688 2708 1718 2730
rect 1905 2701 1935 2727
rect 1983 2723 2049 2739
rect 2175 2773 2241 2789
rect 2175 2739 2191 2773
rect 2225 2739 2241 2773
rect 2001 2701 2031 2723
rect 2097 2701 2127 2727
rect 2175 2723 2241 2739
rect 2367 2773 2433 2789
rect 2367 2739 2383 2773
rect 2417 2739 2433 2773
rect 2193 2701 2223 2723
rect 2289 2701 2319 2727
rect 2367 2723 2433 2739
rect 2559 2773 2625 2789
rect 2559 2739 2575 2773
rect 2609 2739 2625 2773
rect 2385 2701 2415 2723
rect 2481 2701 2511 2727
rect 2559 2723 2625 2739
rect 2751 2773 2817 2789
rect 2751 2739 2767 2773
rect 2801 2739 2817 2773
rect 2577 2701 2607 2723
rect 2673 2701 2703 2727
rect 2751 2723 2817 2739
rect 2943 2773 3009 2789
rect 2943 2739 2959 2773
rect 2993 2739 3009 2773
rect 2769 2701 2799 2723
rect 2865 2701 2895 2727
rect 2943 2723 3009 2739
rect 3150 2780 3216 2796
rect 3150 2746 3166 2780
rect 3200 2746 3216 2780
rect 3150 2730 3216 2746
rect 2961 2701 2991 2723
rect 3168 2708 3198 2730
rect 1688 2486 1718 2508
rect 1670 2470 1736 2486
rect 1670 2436 1686 2470
rect 1720 2436 1736 2470
rect 1670 2420 1736 2436
rect 1488 1686 1518 1708
rect 1470 1670 1536 1686
rect 1905 1680 1935 1701
rect 2001 1680 2031 1701
rect 2097 1680 2127 1701
rect 2193 1680 2223 1701
rect 2289 1680 2319 1701
rect 2385 1680 2415 1701
rect 2481 1680 2511 1701
rect 2577 1680 2607 1701
rect 2673 1680 2703 1701
rect 2769 1680 2799 1701
rect 2865 1680 2895 1701
rect 1900 1679 2896 1680
rect 1470 1636 1486 1670
rect 1520 1636 1536 1670
rect 1470 1620 1536 1636
rect 1887 1670 2913 1679
rect 2961 1670 2991 1701
rect 3168 1686 3198 1708
rect 1887 1663 2991 1670
rect 1887 1629 1903 1663
rect 1937 1629 2095 1663
rect 2129 1629 2287 1663
rect 2321 1629 2479 1663
rect 2513 1629 2671 1663
rect 2705 1629 2863 1663
rect 2897 1629 2991 1663
rect 1887 1620 2991 1629
rect 3150 1670 3216 1686
rect 3150 1636 3166 1670
rect 3200 1636 3216 1670
rect 3150 1620 3216 1636
rect 1887 1613 2990 1620
rect 1900 1610 2990 1613
rect 4770 2780 4836 2796
rect 4770 2746 4786 2780
rect 4820 2746 4836 2780
rect 4770 2730 4836 2746
rect 4970 2780 5036 2796
rect 4970 2746 4986 2780
rect 5020 2746 5036 2780
rect 4970 2730 5036 2746
rect 5283 2773 5349 2789
rect 5283 2739 5299 2773
rect 5333 2739 5349 2773
rect 4788 2708 4818 2730
rect 4988 2708 5018 2730
rect 5205 2701 5235 2727
rect 5283 2723 5349 2739
rect 5475 2773 5541 2789
rect 5475 2739 5491 2773
rect 5525 2739 5541 2773
rect 5301 2701 5331 2723
rect 5397 2701 5427 2727
rect 5475 2723 5541 2739
rect 5667 2773 5733 2789
rect 5667 2739 5683 2773
rect 5717 2739 5733 2773
rect 5493 2701 5523 2723
rect 5589 2701 5619 2727
rect 5667 2723 5733 2739
rect 5859 2773 5925 2789
rect 5859 2739 5875 2773
rect 5909 2739 5925 2773
rect 5685 2701 5715 2723
rect 5781 2701 5811 2727
rect 5859 2723 5925 2739
rect 6051 2773 6117 2789
rect 6051 2739 6067 2773
rect 6101 2739 6117 2773
rect 5877 2701 5907 2723
rect 5973 2701 6003 2727
rect 6051 2723 6117 2739
rect 6243 2773 6309 2789
rect 6243 2739 6259 2773
rect 6293 2739 6309 2773
rect 6069 2701 6099 2723
rect 6165 2701 6195 2727
rect 6243 2723 6309 2739
rect 6450 2780 6516 2796
rect 6450 2746 6466 2780
rect 6500 2746 6516 2780
rect 6450 2730 6516 2746
rect 6261 2701 6291 2723
rect 6468 2708 6498 2730
rect 4988 2486 5018 2508
rect 4970 2470 5036 2486
rect 4970 2436 4986 2470
rect 5020 2436 5036 2470
rect 4970 2420 5036 2436
rect 4788 1686 4818 1708
rect 4770 1670 4836 1686
rect 5205 1680 5235 1701
rect 5301 1680 5331 1701
rect 5397 1680 5427 1701
rect 5493 1680 5523 1701
rect 5589 1680 5619 1701
rect 5685 1680 5715 1701
rect 5781 1680 5811 1701
rect 5877 1680 5907 1701
rect 5973 1680 6003 1701
rect 6069 1680 6099 1701
rect 6165 1680 6195 1701
rect 5200 1679 6196 1680
rect 4770 1636 4786 1670
rect 4820 1636 4836 1670
rect 4770 1620 4836 1636
rect 5187 1670 6213 1679
rect 6261 1670 6291 1701
rect 6468 1686 6498 1708
rect 5187 1663 6291 1670
rect 5187 1629 5203 1663
rect 5237 1629 5395 1663
rect 5429 1629 5587 1663
rect 5621 1629 5779 1663
rect 5813 1629 5971 1663
rect 6005 1629 6163 1663
rect 6197 1629 6291 1663
rect 5187 1620 6291 1629
rect 6450 1670 6516 1686
rect 6450 1636 6466 1670
rect 6500 1636 6516 1670
rect 6450 1620 6516 1636
rect 5187 1613 6290 1620
rect 5200 1610 6290 1613
rect 8070 2780 8136 2796
rect 8070 2746 8086 2780
rect 8120 2746 8136 2780
rect 8070 2730 8136 2746
rect 8270 2780 8336 2796
rect 8270 2746 8286 2780
rect 8320 2746 8336 2780
rect 8270 2730 8336 2746
rect 8583 2773 8649 2789
rect 8583 2739 8599 2773
rect 8633 2739 8649 2773
rect 8088 2708 8118 2730
rect 8288 2708 8318 2730
rect 8505 2701 8535 2727
rect 8583 2723 8649 2739
rect 8775 2773 8841 2789
rect 8775 2739 8791 2773
rect 8825 2739 8841 2773
rect 8601 2701 8631 2723
rect 8697 2701 8727 2727
rect 8775 2723 8841 2739
rect 8967 2773 9033 2789
rect 8967 2739 8983 2773
rect 9017 2739 9033 2773
rect 8793 2701 8823 2723
rect 8889 2701 8919 2727
rect 8967 2723 9033 2739
rect 9159 2773 9225 2789
rect 9159 2739 9175 2773
rect 9209 2739 9225 2773
rect 8985 2701 9015 2723
rect 9081 2701 9111 2727
rect 9159 2723 9225 2739
rect 9351 2773 9417 2789
rect 9351 2739 9367 2773
rect 9401 2739 9417 2773
rect 9177 2701 9207 2723
rect 9273 2701 9303 2727
rect 9351 2723 9417 2739
rect 9543 2773 9609 2789
rect 9543 2739 9559 2773
rect 9593 2739 9609 2773
rect 9369 2701 9399 2723
rect 9465 2701 9495 2727
rect 9543 2723 9609 2739
rect 9750 2780 9816 2796
rect 9750 2746 9766 2780
rect 9800 2746 9816 2780
rect 9750 2730 9816 2746
rect 9561 2701 9591 2723
rect 9768 2708 9798 2730
rect 8288 2486 8318 2508
rect 8270 2470 8336 2486
rect 8270 2436 8286 2470
rect 8320 2436 8336 2470
rect 8270 2420 8336 2436
rect 8088 1686 8118 1708
rect 8070 1670 8136 1686
rect 8505 1680 8535 1701
rect 8601 1680 8631 1701
rect 8697 1680 8727 1701
rect 8793 1680 8823 1701
rect 8889 1680 8919 1701
rect 8985 1680 9015 1701
rect 9081 1680 9111 1701
rect 9177 1680 9207 1701
rect 9273 1680 9303 1701
rect 9369 1680 9399 1701
rect 9465 1680 9495 1701
rect 8500 1679 9496 1680
rect 8070 1636 8086 1670
rect 8120 1636 8136 1670
rect 8070 1620 8136 1636
rect 8487 1670 9513 1679
rect 9561 1670 9591 1701
rect 9768 1686 9798 1708
rect 8487 1663 9591 1670
rect 8487 1629 8503 1663
rect 8537 1629 8695 1663
rect 8729 1629 8887 1663
rect 8921 1629 9079 1663
rect 9113 1629 9271 1663
rect 9305 1629 9463 1663
rect 9497 1629 9591 1663
rect 8487 1620 9591 1629
rect 9750 1670 9816 1686
rect 9750 1636 9766 1670
rect 9800 1636 9816 1670
rect 9750 1620 9816 1636
rect 8487 1613 9590 1620
rect 8500 1610 9590 1613
rect 11370 2780 11436 2796
rect 11370 2746 11386 2780
rect 11420 2746 11436 2780
rect 11370 2730 11436 2746
rect 11570 2780 11636 2796
rect 11570 2746 11586 2780
rect 11620 2746 11636 2780
rect 11570 2730 11636 2746
rect 11883 2773 11949 2789
rect 11883 2739 11899 2773
rect 11933 2739 11949 2773
rect 11388 2708 11418 2730
rect 11588 2708 11618 2730
rect 11805 2701 11835 2727
rect 11883 2723 11949 2739
rect 12075 2773 12141 2789
rect 12075 2739 12091 2773
rect 12125 2739 12141 2773
rect 11901 2701 11931 2723
rect 11997 2701 12027 2727
rect 12075 2723 12141 2739
rect 12267 2773 12333 2789
rect 12267 2739 12283 2773
rect 12317 2739 12333 2773
rect 12093 2701 12123 2723
rect 12189 2701 12219 2727
rect 12267 2723 12333 2739
rect 12459 2773 12525 2789
rect 12459 2739 12475 2773
rect 12509 2739 12525 2773
rect 12285 2701 12315 2723
rect 12381 2701 12411 2727
rect 12459 2723 12525 2739
rect 12651 2773 12717 2789
rect 12651 2739 12667 2773
rect 12701 2739 12717 2773
rect 12477 2701 12507 2723
rect 12573 2701 12603 2727
rect 12651 2723 12717 2739
rect 12843 2773 12909 2789
rect 12843 2739 12859 2773
rect 12893 2739 12909 2773
rect 12669 2701 12699 2723
rect 12765 2701 12795 2727
rect 12843 2723 12909 2739
rect 13050 2780 13116 2796
rect 13050 2746 13066 2780
rect 13100 2746 13116 2780
rect 13050 2730 13116 2746
rect 12861 2701 12891 2723
rect 13068 2708 13098 2730
rect 11588 2486 11618 2508
rect 11570 2470 11636 2486
rect 11570 2436 11586 2470
rect 11620 2436 11636 2470
rect 11570 2420 11636 2436
rect 11388 1686 11418 1708
rect 11370 1670 11436 1686
rect 11805 1680 11835 1701
rect 11901 1680 11931 1701
rect 11997 1680 12027 1701
rect 12093 1680 12123 1701
rect 12189 1680 12219 1701
rect 12285 1680 12315 1701
rect 12381 1680 12411 1701
rect 12477 1680 12507 1701
rect 12573 1680 12603 1701
rect 12669 1680 12699 1701
rect 12765 1680 12795 1701
rect 11800 1679 12796 1680
rect 11370 1636 11386 1670
rect 11420 1636 11436 1670
rect 11370 1620 11436 1636
rect 11787 1670 12813 1679
rect 12861 1670 12891 1701
rect 13068 1686 13098 1708
rect 11787 1663 12891 1670
rect 11787 1629 11803 1663
rect 11837 1629 11995 1663
rect 12029 1629 12187 1663
rect 12221 1629 12379 1663
rect 12413 1629 12571 1663
rect 12605 1629 12763 1663
rect 12797 1629 12891 1663
rect 11787 1620 12891 1629
rect 13050 1670 13116 1686
rect 13050 1636 13066 1670
rect 13100 1636 13116 1670
rect 13050 1620 13116 1636
rect 11787 1613 12890 1620
rect 11800 1610 12890 1613
rect 14970 2780 15036 2796
rect 14970 2746 14986 2780
rect 15020 2746 15036 2780
rect 14970 2730 15036 2746
rect 15170 2780 15236 2796
rect 15170 2746 15186 2780
rect 15220 2746 15236 2780
rect 15170 2730 15236 2746
rect 15483 2773 15549 2789
rect 15483 2739 15499 2773
rect 15533 2739 15549 2773
rect 14988 2708 15018 2730
rect 15188 2708 15218 2730
rect 15405 2701 15435 2727
rect 15483 2723 15549 2739
rect 15675 2773 15741 2789
rect 15675 2739 15691 2773
rect 15725 2739 15741 2773
rect 15501 2701 15531 2723
rect 15597 2701 15627 2727
rect 15675 2723 15741 2739
rect 15867 2773 15933 2789
rect 15867 2739 15883 2773
rect 15917 2739 15933 2773
rect 15693 2701 15723 2723
rect 15789 2701 15819 2727
rect 15867 2723 15933 2739
rect 16059 2773 16125 2789
rect 16059 2739 16075 2773
rect 16109 2739 16125 2773
rect 15885 2701 15915 2723
rect 15981 2701 16011 2727
rect 16059 2723 16125 2739
rect 16251 2773 16317 2789
rect 16251 2739 16267 2773
rect 16301 2739 16317 2773
rect 16077 2701 16107 2723
rect 16173 2701 16203 2727
rect 16251 2723 16317 2739
rect 16443 2773 16509 2789
rect 16443 2739 16459 2773
rect 16493 2739 16509 2773
rect 16269 2701 16299 2723
rect 16365 2701 16395 2727
rect 16443 2723 16509 2739
rect 16650 2780 16716 2796
rect 16650 2746 16666 2780
rect 16700 2746 16716 2780
rect 16650 2730 16716 2746
rect 16461 2701 16491 2723
rect 16668 2708 16698 2730
rect 15188 2486 15218 2508
rect 15170 2470 15236 2486
rect 15170 2436 15186 2470
rect 15220 2436 15236 2470
rect 15170 2420 15236 2436
rect 14988 1686 15018 1708
rect 14970 1670 15036 1686
rect 15405 1680 15435 1701
rect 15501 1680 15531 1701
rect 15597 1680 15627 1701
rect 15693 1680 15723 1701
rect 15789 1680 15819 1701
rect 15885 1680 15915 1701
rect 15981 1680 16011 1701
rect 16077 1680 16107 1701
rect 16173 1680 16203 1701
rect 16269 1680 16299 1701
rect 16365 1680 16395 1701
rect 15400 1679 16396 1680
rect 14970 1636 14986 1670
rect 15020 1636 15036 1670
rect 14970 1620 15036 1636
rect 15387 1670 16413 1679
rect 16461 1670 16491 1701
rect 16668 1686 16698 1708
rect 15387 1663 16491 1670
rect 15387 1629 15403 1663
rect 15437 1629 15595 1663
rect 15629 1629 15787 1663
rect 15821 1629 15979 1663
rect 16013 1629 16171 1663
rect 16205 1629 16363 1663
rect 16397 1629 16491 1663
rect 15387 1620 16491 1629
rect 16650 1670 16716 1686
rect 16650 1636 16666 1670
rect 16700 1636 16716 1670
rect 16650 1620 16716 1636
rect 15387 1613 16490 1620
rect 15400 1610 16490 1613
rect 18470 2780 18536 2796
rect 18470 2746 18486 2780
rect 18520 2746 18536 2780
rect 18470 2730 18536 2746
rect 18670 2780 18736 2796
rect 18670 2746 18686 2780
rect 18720 2746 18736 2780
rect 18670 2730 18736 2746
rect 18983 2773 19049 2789
rect 18983 2739 18999 2773
rect 19033 2739 19049 2773
rect 18488 2708 18518 2730
rect 18688 2708 18718 2730
rect 18905 2701 18935 2727
rect 18983 2723 19049 2739
rect 19175 2773 19241 2789
rect 19175 2739 19191 2773
rect 19225 2739 19241 2773
rect 19001 2701 19031 2723
rect 19097 2701 19127 2727
rect 19175 2723 19241 2739
rect 19367 2773 19433 2789
rect 19367 2739 19383 2773
rect 19417 2739 19433 2773
rect 19193 2701 19223 2723
rect 19289 2701 19319 2727
rect 19367 2723 19433 2739
rect 19559 2773 19625 2789
rect 19559 2739 19575 2773
rect 19609 2739 19625 2773
rect 19385 2701 19415 2723
rect 19481 2701 19511 2727
rect 19559 2723 19625 2739
rect 19751 2773 19817 2789
rect 19751 2739 19767 2773
rect 19801 2739 19817 2773
rect 19577 2701 19607 2723
rect 19673 2701 19703 2727
rect 19751 2723 19817 2739
rect 19943 2773 20009 2789
rect 19943 2739 19959 2773
rect 19993 2739 20009 2773
rect 19769 2701 19799 2723
rect 19865 2701 19895 2727
rect 19943 2723 20009 2739
rect 20150 2780 20216 2796
rect 20150 2746 20166 2780
rect 20200 2746 20216 2780
rect 20150 2730 20216 2746
rect 19961 2701 19991 2723
rect 20168 2708 20198 2730
rect 18688 2486 18718 2508
rect 18670 2470 18736 2486
rect 18670 2436 18686 2470
rect 18720 2436 18736 2470
rect 18670 2420 18736 2436
rect 18488 1686 18518 1708
rect 18470 1670 18536 1686
rect 18905 1680 18935 1701
rect 19001 1680 19031 1701
rect 19097 1680 19127 1701
rect 19193 1680 19223 1701
rect 19289 1680 19319 1701
rect 19385 1680 19415 1701
rect 19481 1680 19511 1701
rect 19577 1680 19607 1701
rect 19673 1680 19703 1701
rect 19769 1680 19799 1701
rect 19865 1680 19895 1701
rect 18900 1679 19896 1680
rect 18470 1636 18486 1670
rect 18520 1636 18536 1670
rect 18470 1620 18536 1636
rect 18887 1670 19913 1679
rect 19961 1670 19991 1701
rect 20168 1686 20198 1708
rect 18887 1663 19991 1670
rect 18887 1629 18903 1663
rect 18937 1629 19095 1663
rect 19129 1629 19287 1663
rect 19321 1629 19479 1663
rect 19513 1629 19671 1663
rect 19705 1629 19863 1663
rect 19897 1629 19991 1663
rect 18887 1620 19991 1629
rect 20150 1670 20216 1686
rect 20150 1636 20166 1670
rect 20200 1636 20216 1670
rect 20150 1620 20216 1636
rect 18887 1613 19990 1620
rect 18900 1610 19990 1613
rect 22170 2780 22236 2796
rect 22170 2746 22186 2780
rect 22220 2746 22236 2780
rect 22170 2730 22236 2746
rect 22370 2780 22436 2796
rect 22370 2746 22386 2780
rect 22420 2746 22436 2780
rect 22370 2730 22436 2746
rect 22683 2773 22749 2789
rect 22683 2739 22699 2773
rect 22733 2739 22749 2773
rect 22188 2708 22218 2730
rect 22388 2708 22418 2730
rect 22605 2701 22635 2727
rect 22683 2723 22749 2739
rect 22875 2773 22941 2789
rect 22875 2739 22891 2773
rect 22925 2739 22941 2773
rect 22701 2701 22731 2723
rect 22797 2701 22827 2727
rect 22875 2723 22941 2739
rect 23067 2773 23133 2789
rect 23067 2739 23083 2773
rect 23117 2739 23133 2773
rect 22893 2701 22923 2723
rect 22989 2701 23019 2727
rect 23067 2723 23133 2739
rect 23259 2773 23325 2789
rect 23259 2739 23275 2773
rect 23309 2739 23325 2773
rect 23085 2701 23115 2723
rect 23181 2701 23211 2727
rect 23259 2723 23325 2739
rect 23451 2773 23517 2789
rect 23451 2739 23467 2773
rect 23501 2739 23517 2773
rect 23277 2701 23307 2723
rect 23373 2701 23403 2727
rect 23451 2723 23517 2739
rect 23643 2773 23709 2789
rect 23643 2739 23659 2773
rect 23693 2739 23709 2773
rect 23469 2701 23499 2723
rect 23565 2701 23595 2727
rect 23643 2723 23709 2739
rect 23850 2780 23916 2796
rect 23850 2746 23866 2780
rect 23900 2746 23916 2780
rect 23850 2730 23916 2746
rect 23661 2701 23691 2723
rect 23868 2708 23898 2730
rect 22388 2486 22418 2508
rect 22370 2470 22436 2486
rect 22370 2436 22386 2470
rect 22420 2436 22436 2470
rect 22370 2420 22436 2436
rect 22188 1686 22218 1708
rect 22170 1670 22236 1686
rect 22605 1680 22635 1701
rect 22701 1680 22731 1701
rect 22797 1680 22827 1701
rect 22893 1680 22923 1701
rect 22989 1680 23019 1701
rect 23085 1680 23115 1701
rect 23181 1680 23211 1701
rect 23277 1680 23307 1701
rect 23373 1680 23403 1701
rect 23469 1680 23499 1701
rect 23565 1680 23595 1701
rect 22600 1679 23596 1680
rect 22170 1636 22186 1670
rect 22220 1636 22236 1670
rect 22170 1620 22236 1636
rect 22587 1670 23613 1679
rect 23661 1670 23691 1701
rect 23868 1686 23898 1708
rect 22587 1663 23691 1670
rect 22587 1629 22603 1663
rect 22637 1629 22795 1663
rect 22829 1629 22987 1663
rect 23021 1629 23179 1663
rect 23213 1629 23371 1663
rect 23405 1629 23563 1663
rect 23597 1629 23691 1663
rect 22587 1620 23691 1629
rect 23850 1670 23916 1686
rect 23850 1636 23866 1670
rect 23900 1636 23916 1670
rect 23850 1620 23916 1636
rect 22587 1613 23690 1620
rect 22600 1610 23690 1613
rect 25970 2780 26036 2796
rect 25970 2746 25986 2780
rect 26020 2746 26036 2780
rect 25970 2730 26036 2746
rect 26170 2780 26236 2796
rect 26170 2746 26186 2780
rect 26220 2746 26236 2780
rect 26170 2730 26236 2746
rect 26483 2773 26549 2789
rect 26483 2739 26499 2773
rect 26533 2739 26549 2773
rect 25988 2708 26018 2730
rect 26188 2708 26218 2730
rect 26405 2701 26435 2727
rect 26483 2723 26549 2739
rect 26675 2773 26741 2789
rect 26675 2739 26691 2773
rect 26725 2739 26741 2773
rect 26501 2701 26531 2723
rect 26597 2701 26627 2727
rect 26675 2723 26741 2739
rect 26867 2773 26933 2789
rect 26867 2739 26883 2773
rect 26917 2739 26933 2773
rect 26693 2701 26723 2723
rect 26789 2701 26819 2727
rect 26867 2723 26933 2739
rect 27059 2773 27125 2789
rect 27059 2739 27075 2773
rect 27109 2739 27125 2773
rect 26885 2701 26915 2723
rect 26981 2701 27011 2727
rect 27059 2723 27125 2739
rect 27251 2773 27317 2789
rect 27251 2739 27267 2773
rect 27301 2739 27317 2773
rect 27077 2701 27107 2723
rect 27173 2701 27203 2727
rect 27251 2723 27317 2739
rect 27443 2773 27509 2789
rect 27443 2739 27459 2773
rect 27493 2739 27509 2773
rect 27269 2701 27299 2723
rect 27365 2701 27395 2727
rect 27443 2723 27509 2739
rect 27650 2780 27716 2796
rect 27650 2746 27666 2780
rect 27700 2746 27716 2780
rect 27650 2730 27716 2746
rect 27461 2701 27491 2723
rect 27668 2708 27698 2730
rect 26188 2486 26218 2508
rect 26170 2470 26236 2486
rect 26170 2436 26186 2470
rect 26220 2436 26236 2470
rect 26170 2420 26236 2436
rect 25988 1686 26018 1708
rect 25970 1670 26036 1686
rect 26405 1680 26435 1701
rect 26501 1680 26531 1701
rect 26597 1680 26627 1701
rect 26693 1680 26723 1701
rect 26789 1680 26819 1701
rect 26885 1680 26915 1701
rect 26981 1680 27011 1701
rect 27077 1680 27107 1701
rect 27173 1680 27203 1701
rect 27269 1680 27299 1701
rect 27365 1680 27395 1701
rect 26400 1679 27396 1680
rect 25970 1636 25986 1670
rect 26020 1636 26036 1670
rect 25970 1620 26036 1636
rect 26387 1670 27413 1679
rect 27461 1670 27491 1701
rect 27668 1686 27698 1708
rect 26387 1663 27491 1670
rect 26387 1629 26403 1663
rect 26437 1629 26595 1663
rect 26629 1629 26787 1663
rect 26821 1629 26979 1663
rect 27013 1629 27171 1663
rect 27205 1629 27363 1663
rect 27397 1629 27491 1663
rect 26387 1620 27491 1629
rect 27650 1670 27716 1686
rect 27650 1636 27666 1670
rect 27700 1636 27716 1670
rect 27650 1620 27716 1636
rect 26387 1613 27490 1620
rect 26400 1610 27490 1613
<< polycont >>
rect 5015 27133 5049 27167
rect 5123 27173 5157 27207
rect 5291 27173 5325 27207
rect 5399 27133 5433 27167
rect 5651 27159 5685 27193
rect 5719 27159 5753 27193
rect 5787 27159 5821 27193
rect 5933 27159 5967 27193
rect 6499 27169 6533 27203
rect 6863 27133 6897 27167
rect 7407 27173 7441 27207
rect 7515 27133 7549 27167
rect 7971 27169 8005 27203
rect 8335 27133 8369 27167
rect 9075 27169 9109 27203
rect 9439 27133 9473 27167
rect 10137 27159 10171 27193
rect 10255 27146 10289 27180
rect 10655 27169 10689 27203
rect 10758 27169 10792 27203
rect 10861 27169 10895 27203
rect 10969 27133 11003 27167
rect 11068 27133 11102 27167
rect 11167 27133 11201 27167
rect 11651 27169 11685 27203
rect 12015 27133 12049 27167
rect 12559 27173 12593 27207
rect 12667 27133 12701 27167
rect 13123 27169 13157 27203
rect 13487 27133 13521 27167
rect 14227 27169 14261 27203
rect 14591 27133 14625 27167
rect 15135 27173 15169 27207
rect 15243 27133 15277 27167
rect 15699 27169 15733 27203
rect 16063 27133 16097 27167
rect 16803 27169 16837 27203
rect 17167 27133 17201 27167
rect 17831 27169 17865 27203
rect 17934 27169 17968 27203
rect 18037 27169 18071 27203
rect 18145 27133 18179 27167
rect 18244 27133 18278 27167
rect 18343 27133 18377 27167
rect 18623 27159 18657 27193
rect 18691 27159 18725 27193
rect 18759 27159 18793 27193
rect 18905 27159 18939 27193
rect 19303 27169 19337 27203
rect 19406 27169 19440 27203
rect 19509 27169 19543 27203
rect 19617 27133 19651 27167
rect 19716 27133 19750 27167
rect 19815 27133 19849 27167
rect 20011 27173 20045 27207
rect 20119 27133 20153 27167
rect 5015 26561 5049 26595
rect 5123 26521 5157 26555
rect 5503 26525 5537 26559
rect 5606 26525 5640 26559
rect 5709 26525 5743 26559
rect 5817 26561 5851 26595
rect 5916 26561 5950 26595
rect 6015 26561 6049 26595
rect 6499 26525 6533 26559
rect 6863 26561 6897 26595
rect 7527 26525 7561 26559
rect 7637 26525 7671 26559
rect 7745 26561 7779 26595
rect 7855 26561 7889 26595
rect 8339 26525 8373 26559
rect 8703 26561 8737 26595
rect 9443 26525 9477 26559
rect 9807 26561 9841 26595
rect 10547 26525 10581 26559
rect 10911 26561 10945 26595
rect 11651 26525 11685 26559
rect 12015 26561 12049 26595
rect 12679 26525 12713 26559
rect 12789 26525 12823 26559
rect 12897 26561 12931 26595
rect 13007 26561 13041 26595
rect 13491 26525 13525 26559
rect 13855 26561 13889 26595
rect 14595 26525 14629 26559
rect 14959 26561 14993 26595
rect 15699 26525 15733 26559
rect 16063 26561 16097 26595
rect 16803 26525 16837 26559
rect 17167 26561 17201 26595
rect 18091 26525 18125 26559
rect 18455 26561 18489 26595
rect 19195 26525 19229 26559
rect 19559 26561 19593 26595
rect 20011 26521 20045 26555
rect 20119 26561 20153 26595
rect 5015 26045 5049 26079
rect 5123 26085 5157 26119
rect 5763 26081 5797 26115
rect 6127 26045 6161 26079
rect 6867 26081 6901 26115
rect 7231 26045 7265 26079
rect 7971 26081 8005 26115
rect 8335 26045 8369 26079
rect 9075 26081 9109 26115
rect 9439 26045 9473 26079
rect 10103 26081 10137 26115
rect 10213 26081 10247 26115
rect 10321 26045 10355 26079
rect 10431 26045 10465 26079
rect 10915 26081 10949 26115
rect 11279 26045 11313 26079
rect 12019 26081 12053 26115
rect 12383 26045 12417 26079
rect 13123 26081 13157 26115
rect 13487 26045 13521 26079
rect 14227 26081 14261 26115
rect 14591 26045 14625 26079
rect 15197 26081 15231 26115
rect 15457 26045 15491 26079
rect 15883 26081 15917 26115
rect 16247 26045 16281 26079
rect 16987 26081 17021 26115
rect 17351 26045 17385 26079
rect 18091 26081 18125 26115
rect 18455 26045 18489 26079
rect 19195 26081 19229 26115
rect 19559 26045 19593 26079
rect 20011 26085 20045 26119
rect 20119 26045 20153 26079
rect 5015 25473 5049 25507
rect 5123 25433 5157 25467
rect 5503 25437 5537 25471
rect 5606 25437 5640 25471
rect 5709 25437 5743 25471
rect 5817 25473 5851 25507
rect 5916 25473 5950 25507
rect 6015 25473 6049 25507
rect 6499 25437 6533 25471
rect 6863 25473 6897 25507
rect 7527 25437 7561 25471
rect 7637 25437 7671 25471
rect 7745 25473 7779 25507
rect 7855 25473 7889 25507
rect 8339 25437 8373 25471
rect 8703 25473 8737 25507
rect 9443 25437 9477 25471
rect 9807 25473 9841 25507
rect 10547 25437 10581 25471
rect 10911 25473 10945 25507
rect 11651 25437 11685 25471
rect 12015 25473 12049 25507
rect 12679 25437 12713 25471
rect 12789 25437 12823 25471
rect 12897 25473 12931 25507
rect 13007 25473 13041 25507
rect 13491 25437 13525 25471
rect 13855 25473 13889 25507
rect 14595 25437 14629 25471
rect 14959 25473 14993 25507
rect 15699 25437 15733 25471
rect 16063 25473 16097 25507
rect 16803 25437 16837 25471
rect 17167 25473 17201 25507
rect 18091 25437 18125 25471
rect 18455 25473 18489 25507
rect 19195 25437 19229 25471
rect 19559 25473 19593 25507
rect 20011 25433 20045 25467
rect 20119 25473 20153 25507
rect 5015 24957 5049 24991
rect 5123 24997 5157 25031
rect 5763 24993 5797 25027
rect 6127 24957 6161 24991
rect 6867 24993 6901 25027
rect 7231 24957 7265 24991
rect 7971 24993 8005 25027
rect 8335 24957 8369 24991
rect 9075 24993 9109 25027
rect 9439 24957 9473 24991
rect 10103 24993 10137 25027
rect 10213 24993 10247 25027
rect 10321 24957 10355 24991
rect 10431 24957 10465 24991
rect 10915 24993 10949 25027
rect 11279 24957 11313 24991
rect 12019 24993 12053 25027
rect 12383 24957 12417 24991
rect 13123 24993 13157 25027
rect 13487 24957 13521 24991
rect 14227 24993 14261 25027
rect 14591 24957 14625 24991
rect 15197 24993 15231 25027
rect 15457 24957 15491 24991
rect 15883 24993 15917 25027
rect 16247 24957 16281 24991
rect 16987 24993 17021 25027
rect 17351 24957 17385 24991
rect 18091 24993 18125 25027
rect 18455 24957 18489 24991
rect 19195 24993 19229 25027
rect 19559 24957 19593 24991
rect 20011 24997 20045 25031
rect 20119 24957 20153 24991
rect 5015 24385 5049 24419
rect 5123 24345 5157 24379
rect 5503 24349 5537 24383
rect 5606 24349 5640 24383
rect 5709 24349 5743 24383
rect 5817 24385 5851 24419
rect 5916 24385 5950 24419
rect 6015 24385 6049 24419
rect 6499 24349 6533 24383
rect 6863 24385 6897 24419
rect 7527 24349 7561 24383
rect 7637 24349 7671 24383
rect 7745 24385 7779 24419
rect 7855 24385 7889 24419
rect 8339 24349 8373 24383
rect 8703 24385 8737 24419
rect 9443 24349 9477 24383
rect 9807 24385 9841 24419
rect 10547 24349 10581 24383
rect 10911 24385 10945 24419
rect 11651 24349 11685 24383
rect 12015 24385 12049 24419
rect 12679 24349 12713 24383
rect 12789 24349 12823 24383
rect 12897 24385 12931 24419
rect 13007 24385 13041 24419
rect 13491 24349 13525 24383
rect 13855 24385 13889 24419
rect 14595 24349 14629 24383
rect 14959 24385 14993 24419
rect 15699 24349 15733 24383
rect 16063 24385 16097 24419
rect 16803 24349 16837 24383
rect 17167 24385 17201 24419
rect 18091 24349 18125 24383
rect 18455 24385 18489 24419
rect 19195 24349 19229 24383
rect 19559 24385 19593 24419
rect 20011 24345 20045 24379
rect 20119 24385 20153 24419
rect 5015 23869 5049 23903
rect 5123 23909 5157 23943
rect 5763 23905 5797 23939
rect 6127 23869 6161 23903
rect 6867 23905 6901 23939
rect 7231 23869 7265 23903
rect 7971 23905 8005 23939
rect 8335 23869 8369 23903
rect 9075 23905 9109 23939
rect 9439 23869 9473 23903
rect 10103 23905 10137 23939
rect 10213 23905 10247 23939
rect 10321 23869 10355 23903
rect 10431 23869 10465 23903
rect 10915 23905 10949 23939
rect 11279 23869 11313 23903
rect 12019 23905 12053 23939
rect 12383 23869 12417 23903
rect 13123 23905 13157 23939
rect 13487 23869 13521 23903
rect 14227 23905 14261 23939
rect 14591 23869 14625 23903
rect 15197 23905 15231 23939
rect 15457 23869 15491 23903
rect 15883 23905 15917 23939
rect 16247 23869 16281 23903
rect 16987 23905 17021 23939
rect 17351 23869 17385 23903
rect 18091 23905 18125 23939
rect 18455 23869 18489 23903
rect 19195 23905 19229 23939
rect 19559 23869 19593 23903
rect 20011 23909 20045 23943
rect 20119 23869 20153 23903
rect 5015 23297 5049 23331
rect 5123 23257 5157 23291
rect 5503 23261 5537 23295
rect 5606 23261 5640 23295
rect 5709 23261 5743 23295
rect 5817 23297 5851 23331
rect 5916 23297 5950 23331
rect 6015 23297 6049 23331
rect 6499 23261 6533 23295
rect 6863 23297 6897 23331
rect 7527 23261 7561 23295
rect 7637 23261 7671 23295
rect 7745 23297 7779 23331
rect 7855 23297 7889 23331
rect 8339 23261 8373 23295
rect 8703 23297 8737 23331
rect 9443 23261 9477 23295
rect 9807 23297 9841 23331
rect 10547 23261 10581 23295
rect 10911 23297 10945 23331
rect 11651 23261 11685 23295
rect 12015 23297 12049 23331
rect 12679 23261 12713 23295
rect 12789 23261 12823 23295
rect 12897 23297 12931 23331
rect 13007 23297 13041 23331
rect 13491 23261 13525 23295
rect 13855 23297 13889 23331
rect 14595 23261 14629 23295
rect 14959 23297 14993 23331
rect 15699 23261 15733 23295
rect 16063 23297 16097 23331
rect 16803 23261 16837 23295
rect 17167 23297 17201 23331
rect 18091 23261 18125 23295
rect 18455 23297 18489 23331
rect 19195 23261 19229 23295
rect 19559 23297 19593 23331
rect 20011 23257 20045 23291
rect 20119 23297 20153 23331
rect 5015 22781 5049 22815
rect 5123 22821 5157 22855
rect 5763 22817 5797 22851
rect 6127 22781 6161 22815
rect 6867 22817 6901 22851
rect 7231 22781 7265 22815
rect 7971 22817 8005 22851
rect 8335 22781 8369 22815
rect 9075 22817 9109 22851
rect 9439 22781 9473 22815
rect 10103 22817 10137 22851
rect 10213 22817 10247 22851
rect 10321 22781 10355 22815
rect 10431 22781 10465 22815
rect 10915 22817 10949 22851
rect 11279 22781 11313 22815
rect 12019 22817 12053 22851
rect 12383 22781 12417 22815
rect 13123 22817 13157 22851
rect 13487 22781 13521 22815
rect 14227 22817 14261 22851
rect 14591 22781 14625 22815
rect 15197 22817 15231 22851
rect 15457 22781 15491 22815
rect 15883 22817 15917 22851
rect 16247 22781 16281 22815
rect 16987 22817 17021 22851
rect 17351 22781 17385 22815
rect 18091 22817 18125 22851
rect 18455 22781 18489 22815
rect 19195 22817 19229 22851
rect 19559 22781 19593 22815
rect 20011 22821 20045 22855
rect 20119 22781 20153 22815
rect 5015 22209 5049 22243
rect 5123 22169 5157 22203
rect 5503 22173 5537 22207
rect 5606 22173 5640 22207
rect 5709 22173 5743 22207
rect 5817 22209 5851 22243
rect 5916 22209 5950 22243
rect 6015 22209 6049 22243
rect 6499 22173 6533 22207
rect 6863 22209 6897 22243
rect 7527 22173 7561 22207
rect 7637 22173 7671 22207
rect 7745 22209 7779 22243
rect 7855 22209 7889 22243
rect 8339 22173 8373 22207
rect 8703 22209 8737 22243
rect 9443 22173 9477 22207
rect 9807 22209 9841 22243
rect 10547 22173 10581 22207
rect 10911 22209 10945 22243
rect 11651 22173 11685 22207
rect 12015 22209 12049 22243
rect 12679 22173 12713 22207
rect 12789 22173 12823 22207
rect 12897 22209 12931 22243
rect 13007 22209 13041 22243
rect 13491 22173 13525 22207
rect 13855 22209 13889 22243
rect 14595 22173 14629 22207
rect 14959 22209 14993 22243
rect 15699 22173 15733 22207
rect 16063 22209 16097 22243
rect 16803 22173 16837 22207
rect 17167 22209 17201 22243
rect 18091 22173 18125 22207
rect 18455 22209 18489 22243
rect 19195 22173 19229 22207
rect 19559 22209 19593 22243
rect 20011 22169 20045 22203
rect 20119 22209 20153 22243
rect 5015 21693 5049 21727
rect 5123 21733 5157 21767
rect 5763 21729 5797 21763
rect 6127 21693 6161 21727
rect 6867 21729 6901 21763
rect 7231 21693 7265 21727
rect 7971 21729 8005 21763
rect 8335 21693 8369 21727
rect 9075 21729 9109 21763
rect 9439 21693 9473 21727
rect 10103 21729 10137 21763
rect 10213 21729 10247 21763
rect 10321 21693 10355 21727
rect 10431 21693 10465 21727
rect 10915 21729 10949 21763
rect 11279 21693 11313 21727
rect 12019 21729 12053 21763
rect 12383 21693 12417 21727
rect 13123 21729 13157 21763
rect 13487 21693 13521 21727
rect 14227 21729 14261 21763
rect 14591 21693 14625 21727
rect 15197 21729 15231 21763
rect 15457 21693 15491 21727
rect 15883 21729 15917 21763
rect 16247 21693 16281 21727
rect 16987 21729 17021 21763
rect 17351 21693 17385 21727
rect 18091 21729 18125 21763
rect 18455 21693 18489 21727
rect 19195 21729 19229 21763
rect 19559 21693 19593 21727
rect 20011 21733 20045 21767
rect 20119 21693 20153 21727
rect 5015 21121 5049 21155
rect 5123 21081 5157 21115
rect 5503 21085 5537 21119
rect 5606 21085 5640 21119
rect 5709 21085 5743 21119
rect 5817 21121 5851 21155
rect 5916 21121 5950 21155
rect 6015 21121 6049 21155
rect 6499 21085 6533 21119
rect 6863 21121 6897 21155
rect 7527 21085 7561 21119
rect 7637 21085 7671 21119
rect 7745 21121 7779 21155
rect 7855 21121 7889 21155
rect 8339 21085 8373 21119
rect 8703 21121 8737 21155
rect 9443 21085 9477 21119
rect 9807 21121 9841 21155
rect 10547 21085 10581 21119
rect 10911 21121 10945 21155
rect 11651 21085 11685 21119
rect 12015 21121 12049 21155
rect 12679 21085 12713 21119
rect 12789 21085 12823 21119
rect 12897 21121 12931 21155
rect 13007 21121 13041 21155
rect 13491 21085 13525 21119
rect 13855 21121 13889 21155
rect 14595 21085 14629 21119
rect 14959 21121 14993 21155
rect 15699 21085 15733 21119
rect 16063 21121 16097 21155
rect 16803 21085 16837 21119
rect 17167 21121 17201 21155
rect 18091 21085 18125 21119
rect 18455 21121 18489 21155
rect 19195 21085 19229 21119
rect 19559 21121 19593 21155
rect 20011 21081 20045 21115
rect 20119 21121 20153 21155
rect 5015 20605 5049 20639
rect 5123 20645 5157 20679
rect 5763 20641 5797 20675
rect 6127 20605 6161 20639
rect 6867 20641 6901 20675
rect 7231 20605 7265 20639
rect 7971 20641 8005 20675
rect 8335 20605 8369 20639
rect 9075 20641 9109 20675
rect 9439 20605 9473 20639
rect 10103 20641 10137 20675
rect 10213 20641 10247 20675
rect 10321 20605 10355 20639
rect 10431 20605 10465 20639
rect 10915 20641 10949 20675
rect 11279 20605 11313 20639
rect 12019 20641 12053 20675
rect 12383 20605 12417 20639
rect 13123 20641 13157 20675
rect 13487 20605 13521 20639
rect 14227 20641 14261 20675
rect 14591 20605 14625 20639
rect 15197 20641 15231 20675
rect 15457 20605 15491 20639
rect 15883 20641 15917 20675
rect 16247 20605 16281 20639
rect 16987 20641 17021 20675
rect 17351 20605 17385 20639
rect 18091 20641 18125 20675
rect 18455 20605 18489 20639
rect 19195 20641 19229 20675
rect 19559 20605 19593 20639
rect 20011 20645 20045 20679
rect 20119 20605 20153 20639
rect 5015 20033 5049 20067
rect 5123 19993 5157 20027
rect 5503 19997 5537 20031
rect 5606 19997 5640 20031
rect 5709 19997 5743 20031
rect 5817 20033 5851 20067
rect 5916 20033 5950 20067
rect 6015 20033 6049 20067
rect 6499 19997 6533 20031
rect 6863 20033 6897 20067
rect 7527 19997 7561 20031
rect 7637 19997 7671 20031
rect 7745 20033 7779 20067
rect 7855 20033 7889 20067
rect 8339 19997 8373 20031
rect 8703 20033 8737 20067
rect 9443 19997 9477 20031
rect 9807 20033 9841 20067
rect 10547 19997 10581 20031
rect 10911 20033 10945 20067
rect 11651 19997 11685 20031
rect 12015 20033 12049 20067
rect 12679 19997 12713 20031
rect 12789 19997 12823 20031
rect 12897 20033 12931 20067
rect 13007 20033 13041 20067
rect 13491 19997 13525 20031
rect 13855 20033 13889 20067
rect 14595 19997 14629 20031
rect 14959 20033 14993 20067
rect 15699 19997 15733 20031
rect 16063 20033 16097 20067
rect 16803 19997 16837 20031
rect 17167 20033 17201 20067
rect 18091 19997 18125 20031
rect 18455 20033 18489 20067
rect 19195 19997 19229 20031
rect 19559 20033 19593 20067
rect 20011 19993 20045 20027
rect 20119 20033 20153 20067
rect 5015 19517 5049 19551
rect 5123 19557 5157 19591
rect 5763 19553 5797 19587
rect 6127 19517 6161 19551
rect 6867 19553 6901 19587
rect 7231 19517 7265 19551
rect 7971 19553 8005 19587
rect 8335 19517 8369 19551
rect 9075 19553 9109 19587
rect 9439 19517 9473 19551
rect 10103 19553 10137 19587
rect 10213 19553 10247 19587
rect 10321 19517 10355 19551
rect 10431 19517 10465 19551
rect 10915 19553 10949 19587
rect 11279 19517 11313 19551
rect 12019 19553 12053 19587
rect 12383 19517 12417 19551
rect 13123 19553 13157 19587
rect 13487 19517 13521 19551
rect 14227 19553 14261 19587
rect 14591 19517 14625 19551
rect 15197 19553 15231 19587
rect 15457 19517 15491 19551
rect 15883 19553 15917 19587
rect 16247 19517 16281 19551
rect 16987 19553 17021 19587
rect 17351 19517 17385 19551
rect 18091 19553 18125 19587
rect 18455 19517 18489 19551
rect 19195 19553 19229 19587
rect 19559 19517 19593 19551
rect 20011 19557 20045 19591
rect 20119 19517 20153 19551
rect 5015 18945 5049 18979
rect 5123 18905 5157 18939
rect 5503 18909 5537 18943
rect 5606 18909 5640 18943
rect 5709 18909 5743 18943
rect 5817 18945 5851 18979
rect 5916 18945 5950 18979
rect 6015 18945 6049 18979
rect 6499 18909 6533 18943
rect 6863 18945 6897 18979
rect 7527 18909 7561 18943
rect 7637 18909 7671 18943
rect 7745 18945 7779 18979
rect 7855 18945 7889 18979
rect 8339 18909 8373 18943
rect 8703 18945 8737 18979
rect 9443 18909 9477 18943
rect 9807 18945 9841 18979
rect 10547 18909 10581 18943
rect 10911 18945 10945 18979
rect 11651 18909 11685 18943
rect 12015 18945 12049 18979
rect 12679 18909 12713 18943
rect 12789 18909 12823 18943
rect 12897 18945 12931 18979
rect 13007 18945 13041 18979
rect 13491 18909 13525 18943
rect 13855 18945 13889 18979
rect 14595 18909 14629 18943
rect 14959 18945 14993 18979
rect 15699 18909 15733 18943
rect 16063 18945 16097 18979
rect 16803 18909 16837 18943
rect 17167 18945 17201 18979
rect 18091 18909 18125 18943
rect 18455 18945 18489 18979
rect 19195 18909 19229 18943
rect 19559 18945 19593 18979
rect 20011 18905 20045 18939
rect 20119 18945 20153 18979
rect 5015 18429 5049 18463
rect 5123 18469 5157 18503
rect 5763 18465 5797 18499
rect 6127 18429 6161 18463
rect 6867 18465 6901 18499
rect 7231 18429 7265 18463
rect 7971 18465 8005 18499
rect 8335 18429 8369 18463
rect 9075 18465 9109 18499
rect 9439 18429 9473 18463
rect 10103 18465 10137 18499
rect 10213 18465 10247 18499
rect 10321 18429 10355 18463
rect 10431 18429 10465 18463
rect 10915 18465 10949 18499
rect 11279 18429 11313 18463
rect 12019 18465 12053 18499
rect 12383 18429 12417 18463
rect 13123 18465 13157 18499
rect 13487 18429 13521 18463
rect 14227 18465 14261 18499
rect 14591 18429 14625 18463
rect 15197 18465 15231 18499
rect 15457 18429 15491 18463
rect 15883 18465 15917 18499
rect 16247 18429 16281 18463
rect 16987 18465 17021 18499
rect 17351 18429 17385 18463
rect 18091 18465 18125 18499
rect 18455 18429 18489 18463
rect 19195 18465 19229 18499
rect 19559 18429 19593 18463
rect 20011 18469 20045 18503
rect 20119 18429 20153 18463
rect 5015 17857 5049 17891
rect 5123 17817 5157 17851
rect 5503 17821 5537 17855
rect 5606 17821 5640 17855
rect 5709 17821 5743 17855
rect 5817 17857 5851 17891
rect 5916 17857 5950 17891
rect 6015 17857 6049 17891
rect 6499 17821 6533 17855
rect 6863 17857 6897 17891
rect 7527 17821 7561 17855
rect 7637 17821 7671 17855
rect 7745 17857 7779 17891
rect 7855 17857 7889 17891
rect 8339 17821 8373 17855
rect 8703 17857 8737 17891
rect 9443 17821 9477 17855
rect 9807 17857 9841 17891
rect 10547 17821 10581 17855
rect 10911 17857 10945 17891
rect 11651 17821 11685 17855
rect 12015 17857 12049 17891
rect 12679 17821 12713 17855
rect 12789 17821 12823 17855
rect 12897 17857 12931 17891
rect 13007 17857 13041 17891
rect 13491 17821 13525 17855
rect 13855 17857 13889 17891
rect 14595 17821 14629 17855
rect 14959 17857 14993 17891
rect 15699 17821 15733 17855
rect 16063 17857 16097 17891
rect 16803 17821 16837 17855
rect 17167 17857 17201 17891
rect 18091 17821 18125 17855
rect 18455 17857 18489 17891
rect 19195 17821 19229 17855
rect 19559 17857 19593 17891
rect 20011 17817 20045 17851
rect 20119 17857 20153 17891
rect 5015 17341 5049 17375
rect 5123 17381 5157 17415
rect 5763 17377 5797 17411
rect 6127 17341 6161 17375
rect 6867 17377 6901 17411
rect 7231 17341 7265 17375
rect 7971 17377 8005 17411
rect 8335 17341 8369 17375
rect 9075 17377 9109 17411
rect 9439 17341 9473 17375
rect 10103 17377 10137 17411
rect 10213 17377 10247 17411
rect 10321 17341 10355 17375
rect 10431 17341 10465 17375
rect 10915 17377 10949 17411
rect 11279 17341 11313 17375
rect 12019 17377 12053 17411
rect 12383 17341 12417 17375
rect 13123 17377 13157 17411
rect 13487 17341 13521 17375
rect 14227 17377 14261 17411
rect 14591 17341 14625 17375
rect 15197 17377 15231 17411
rect 15457 17341 15491 17375
rect 15883 17377 15917 17411
rect 16247 17341 16281 17375
rect 16987 17377 17021 17411
rect 17351 17341 17385 17375
rect 18091 17377 18125 17411
rect 18455 17341 18489 17375
rect 19195 17377 19229 17411
rect 19559 17341 19593 17375
rect 20011 17381 20045 17415
rect 20119 17341 20153 17375
rect 5015 16769 5049 16803
rect 5123 16729 5157 16763
rect 5503 16733 5537 16767
rect 5606 16733 5640 16767
rect 5709 16733 5743 16767
rect 5817 16769 5851 16803
rect 5916 16769 5950 16803
rect 6015 16769 6049 16803
rect 6499 16733 6533 16767
rect 6863 16769 6897 16803
rect 7527 16733 7561 16767
rect 7637 16733 7671 16767
rect 7745 16769 7779 16803
rect 7855 16769 7889 16803
rect 8339 16733 8373 16767
rect 8703 16769 8737 16803
rect 9443 16733 9477 16767
rect 9807 16769 9841 16803
rect 10547 16733 10581 16767
rect 10911 16769 10945 16803
rect 11651 16733 11685 16767
rect 12015 16769 12049 16803
rect 12679 16733 12713 16767
rect 12789 16733 12823 16767
rect 12897 16769 12931 16803
rect 13007 16769 13041 16803
rect 13491 16733 13525 16767
rect 13855 16769 13889 16803
rect 14595 16733 14629 16767
rect 14959 16769 14993 16803
rect 15699 16733 15733 16767
rect 16063 16769 16097 16803
rect 16803 16733 16837 16767
rect 17167 16769 17201 16803
rect 18091 16733 18125 16767
rect 18455 16769 18489 16803
rect 19195 16733 19229 16767
rect 19559 16769 19593 16803
rect 20011 16729 20045 16763
rect 20119 16769 20153 16803
rect 5015 16253 5049 16287
rect 5123 16293 5157 16327
rect 5763 16289 5797 16323
rect 6127 16253 6161 16287
rect 6867 16289 6901 16323
rect 7231 16253 7265 16287
rect 7971 16289 8005 16323
rect 8335 16253 8369 16287
rect 9075 16289 9109 16323
rect 9439 16253 9473 16287
rect 10103 16289 10137 16323
rect 10213 16289 10247 16323
rect 10321 16253 10355 16287
rect 10431 16253 10465 16287
rect 10915 16289 10949 16323
rect 11279 16253 11313 16287
rect 12019 16289 12053 16323
rect 12383 16253 12417 16287
rect 13123 16289 13157 16323
rect 13487 16253 13521 16287
rect 14227 16289 14261 16323
rect 14591 16253 14625 16287
rect 15197 16289 15231 16323
rect 15457 16253 15491 16287
rect 15883 16289 15917 16323
rect 16247 16253 16281 16287
rect 16987 16289 17021 16323
rect 17351 16253 17385 16287
rect 18091 16289 18125 16323
rect 18455 16253 18489 16287
rect 19195 16289 19229 16323
rect 19559 16253 19593 16287
rect 20011 16293 20045 16327
rect 20119 16253 20153 16287
rect 5015 15681 5049 15715
rect 5123 15641 5157 15675
rect 5503 15645 5537 15679
rect 5606 15645 5640 15679
rect 5709 15645 5743 15679
rect 5817 15681 5851 15715
rect 5916 15681 5950 15715
rect 6015 15681 6049 15715
rect 6499 15645 6533 15679
rect 6863 15681 6897 15715
rect 7527 15645 7561 15679
rect 7637 15645 7671 15679
rect 7745 15681 7779 15715
rect 7855 15681 7889 15715
rect 8339 15645 8373 15679
rect 8703 15681 8737 15715
rect 9443 15645 9477 15679
rect 9807 15681 9841 15715
rect 10547 15645 10581 15679
rect 10911 15681 10945 15715
rect 11651 15645 11685 15679
rect 12015 15681 12049 15715
rect 12679 15645 12713 15679
rect 12789 15645 12823 15679
rect 12897 15681 12931 15715
rect 13007 15681 13041 15715
rect 13491 15645 13525 15679
rect 13855 15681 13889 15715
rect 14595 15645 14629 15679
rect 14959 15681 14993 15715
rect 15699 15645 15733 15679
rect 16063 15681 16097 15715
rect 16803 15645 16837 15679
rect 17167 15681 17201 15715
rect 18091 15645 18125 15679
rect 18455 15681 18489 15715
rect 19195 15645 19229 15679
rect 19559 15681 19593 15715
rect 20011 15641 20045 15675
rect 20119 15681 20153 15715
rect 5015 15165 5049 15199
rect 5123 15205 5157 15239
rect 5763 15201 5797 15235
rect 6127 15165 6161 15199
rect 6867 15201 6901 15235
rect 7231 15165 7265 15199
rect 7971 15201 8005 15235
rect 8335 15165 8369 15199
rect 9075 15201 9109 15235
rect 9439 15165 9473 15199
rect 10103 15201 10137 15235
rect 10213 15201 10247 15235
rect 10321 15165 10355 15199
rect 10431 15165 10465 15199
rect 10915 15201 10949 15235
rect 11279 15165 11313 15199
rect 12019 15201 12053 15235
rect 12383 15165 12417 15199
rect 12849 15191 12883 15225
rect 12963 15191 12997 15225
rect 13167 15191 13201 15225
rect 13363 15191 13397 15225
rect 13541 15201 13575 15235
rect 13801 15165 13835 15199
rect 14227 15201 14261 15235
rect 14591 15165 14625 15199
rect 15135 15205 15169 15239
rect 15243 15165 15277 15199
rect 15425 15191 15459 15225
rect 15539 15191 15573 15225
rect 15743 15191 15777 15225
rect 15939 15191 15973 15225
rect 16175 15201 16209 15235
rect 16285 15201 16319 15235
rect 16393 15165 16427 15199
rect 16503 15165 16537 15199
rect 16987 15201 17021 15235
rect 17351 15165 17385 15199
rect 18091 15201 18125 15235
rect 18455 15165 18489 15199
rect 19195 15201 19229 15235
rect 19559 15165 19593 15199
rect 20011 15205 20045 15239
rect 20119 15165 20153 15199
rect 5015 14593 5049 14627
rect 5123 14553 5157 14587
rect 5503 14557 5537 14591
rect 5606 14557 5640 14591
rect 5709 14557 5743 14591
rect 5817 14593 5851 14627
rect 5916 14593 5950 14627
rect 6015 14593 6049 14627
rect 6499 14557 6533 14591
rect 6863 14593 6897 14627
rect 7695 14557 7729 14591
rect 8059 14593 8093 14627
rect 8799 14557 8833 14591
rect 9163 14593 9197 14627
rect 9903 14557 9937 14591
rect 10267 14593 10301 14627
rect 10787 14644 10821 14678
rect 10955 14644 10989 14678
rect 10865 14531 10899 14565
rect 11027 14531 11061 14565
rect 11123 14531 11157 14565
rect 11264 14567 11298 14601
rect 11360 14567 11394 14601
rect 11759 14557 11793 14591
rect 11862 14557 11896 14591
rect 11965 14557 11999 14591
rect 12073 14593 12107 14627
rect 12172 14593 12206 14627
rect 12271 14593 12305 14627
rect 12811 14644 12845 14678
rect 12979 14644 13013 14678
rect 12889 14531 12923 14565
rect 13051 14531 13085 14565
rect 13147 14531 13181 14565
rect 13288 14567 13322 14601
rect 13384 14567 13418 14601
rect 13599 14557 13633 14591
rect 13702 14557 13736 14591
rect 13805 14557 13839 14591
rect 13913 14593 13947 14627
rect 14012 14593 14046 14627
rect 14111 14593 14145 14627
rect 14808 14667 14842 14701
rect 14277 14567 14311 14601
rect 14397 14580 14431 14614
rect 14610 14567 14644 14601
rect 14885 14559 14919 14593
rect 15086 14683 15120 14717
rect 14981 14531 15015 14565
rect 15125 14557 15159 14591
rect 15369 14569 15403 14603
rect 15551 14657 15585 14691
rect 15221 14509 15255 14543
rect 15465 14521 15499 14555
rect 15800 14683 15834 14717
rect 15981 14628 16015 14662
rect 15720 14515 15754 14549
rect 15822 14521 15856 14555
rect 16188 14582 16222 14616
rect 16290 14567 16324 14601
rect 16803 14557 16837 14591
rect 17167 14593 17201 14627
rect 18091 14557 18125 14591
rect 18455 14593 18489 14627
rect 19195 14557 19229 14591
rect 19559 14593 19593 14627
rect 20011 14553 20045 14587
rect 20119 14593 20153 14627
rect 5015 14077 5049 14111
rect 5123 14117 5157 14151
rect 5763 14113 5797 14147
rect 6127 14077 6161 14111
rect 6867 14113 6901 14147
rect 7231 14077 7265 14111
rect 7971 14113 8005 14147
rect 8335 14077 8369 14111
rect 9075 14113 9109 14147
rect 9439 14077 9473 14111
rect 10194 14103 10228 14137
rect 10469 14111 10503 14145
rect 10565 14139 10599 14173
rect 10392 14003 10426 14037
rect 10709 14113 10743 14147
rect 10805 14161 10839 14195
rect 10670 13987 10704 14021
rect 10953 14101 10987 14135
rect 11049 14149 11083 14183
rect 11304 14155 11338 14189
rect 11406 14149 11440 14183
rect 11135 14013 11169 14047
rect 11565 14042 11599 14076
rect 11384 13987 11418 14021
rect 11772 14088 11806 14122
rect 11874 14103 11908 14137
rect 12025 14090 12059 14124
rect 12145 14103 12179 14137
rect 12538 14103 12572 14137
rect 12606 14103 12640 14137
rect 12674 14103 12708 14137
rect 12742 14103 12776 14137
rect 12810 14103 12844 14137
rect 12878 14103 12912 14137
rect 12946 14103 12980 14137
rect 13014 14103 13048 14137
rect 13082 14103 13116 14137
rect 13150 14103 13184 14137
rect 13218 14103 13252 14137
rect 13286 14103 13320 14137
rect 13354 14103 13388 14137
rect 13422 14103 13456 14137
rect 13490 14103 13524 14137
rect 13558 14103 13592 14137
rect 13985 14103 14019 14137
rect 14321 14103 14355 14137
rect 14435 14103 14469 14137
rect 14639 14103 14673 14137
rect 14835 14103 14869 14137
rect 15246 14103 15280 14137
rect 15342 14103 15376 14137
rect 15483 14139 15517 14173
rect 15579 14139 15613 14173
rect 15741 14139 15775 14173
rect 15651 14026 15685 14060
rect 16073 14090 16107 14124
rect 16193 14103 16227 14137
rect 16349 14090 16383 14124
rect 15819 14026 15853 14060
rect 16469 14103 16503 14137
rect 16987 14113 17021 14147
rect 17351 14077 17385 14111
rect 18091 14113 18125 14147
rect 18455 14077 18489 14111
rect 19195 14113 19229 14147
rect 19559 14077 19593 14111
rect 20011 14117 20045 14151
rect 20119 14077 20153 14111
rect 5015 13505 5049 13539
rect 5123 13465 5157 13499
rect 5503 13469 5537 13503
rect 5606 13469 5640 13503
rect 5709 13469 5743 13503
rect 5817 13505 5851 13539
rect 5916 13505 5950 13539
rect 6015 13505 6049 13539
rect 6499 13469 6533 13503
rect 6863 13505 6897 13539
rect 7787 13469 7821 13503
rect 8151 13505 8185 13539
rect 8891 13469 8925 13503
rect 9255 13505 9289 13539
rect 9677 13479 9711 13513
rect 9797 13492 9831 13526
rect 10238 13479 10272 13513
rect 10306 13479 10340 13513
rect 10374 13479 10408 13513
rect 10442 13479 10476 13513
rect 10510 13479 10544 13513
rect 10578 13479 10612 13513
rect 10646 13479 10680 13513
rect 10714 13479 10748 13513
rect 10782 13479 10816 13513
rect 10850 13479 10884 13513
rect 10918 13479 10952 13513
rect 10986 13479 11020 13513
rect 11054 13479 11088 13513
rect 11122 13479 11156 13513
rect 11190 13479 11224 13513
rect 11258 13479 11292 13513
rect 11685 13479 11719 13513
rect 11943 13469 11977 13503
rect 12053 13469 12087 13503
rect 12161 13505 12195 13539
rect 12271 13505 12305 13539
rect 12577 13492 12611 13526
rect 13152 13579 13186 13613
rect 12697 13479 12731 13513
rect 12954 13479 12988 13513
rect 13229 13471 13263 13505
rect 13430 13595 13464 13629
rect 13325 13443 13359 13477
rect 13469 13469 13503 13503
rect 13713 13481 13747 13515
rect 13895 13569 13929 13603
rect 13565 13421 13599 13455
rect 13809 13433 13843 13467
rect 14144 13595 14178 13629
rect 14325 13540 14359 13574
rect 14064 13427 14098 13461
rect 14166 13433 14200 13467
rect 14532 13494 14566 13528
rect 14634 13479 14668 13513
rect 14737 13479 14771 13513
rect 15164 13479 15198 13513
rect 15232 13479 15266 13513
rect 15300 13479 15334 13513
rect 15368 13479 15402 13513
rect 15436 13479 15470 13513
rect 15504 13479 15538 13513
rect 15572 13479 15606 13513
rect 15640 13479 15674 13513
rect 15708 13479 15742 13513
rect 15776 13479 15810 13513
rect 15844 13479 15878 13513
rect 15912 13479 15946 13513
rect 15980 13479 16014 13513
rect 16048 13479 16082 13513
rect 16116 13479 16150 13513
rect 16184 13479 16218 13513
rect 16626 13479 16660 13513
rect 16722 13479 16756 13513
rect 17031 13556 17065 13590
rect 16863 13443 16897 13477
rect 17199 13556 17233 13590
rect 16959 13443 16993 13477
rect 17121 13443 17155 13477
rect 18091 13469 18125 13503
rect 18455 13505 18489 13539
rect 19195 13469 19229 13503
rect 19559 13505 19593 13539
rect 20011 13465 20045 13499
rect 20119 13505 20153 13539
rect 5015 12989 5049 13023
rect 5123 13029 5157 13063
rect 5319 13025 5353 13059
rect 5429 13025 5463 13059
rect 5537 12989 5571 13023
rect 5647 12989 5681 13023
rect 6131 13025 6165 13059
rect 6495 12989 6529 13023
rect 7235 13025 7269 13059
rect 7599 12989 7633 13023
rect 8339 13025 8373 13059
rect 8703 12989 8737 13023
rect 9169 13015 9203 13049
rect 9283 13015 9317 13049
rect 9487 13015 9521 13049
rect 9683 13015 9717 13049
rect 10045 13025 10079 13059
rect 10305 12989 10339 13023
rect 10470 13015 10504 13049
rect 10745 13023 10779 13057
rect 10841 13051 10875 13085
rect 10668 12915 10702 12949
rect 10985 13025 11019 13059
rect 11081 13073 11115 13107
rect 10946 12899 10980 12933
rect 11229 13013 11263 13047
rect 11325 13061 11359 13095
rect 11580 13067 11614 13101
rect 11682 13061 11716 13095
rect 11411 12925 11445 12959
rect 11841 12954 11875 12988
rect 11660 12899 11694 12933
rect 12048 13000 12082 13034
rect 12150 13015 12184 13049
rect 12248 13015 12282 13049
rect 12350 13000 12384 13034
rect 12716 13061 12750 13095
rect 12818 13067 12852 13101
rect 12557 12954 12591 12988
rect 12738 12899 12772 12933
rect 13073 13061 13107 13095
rect 13317 13073 13351 13107
rect 12987 12925 13021 12959
rect 13169 13013 13203 13047
rect 13413 13025 13447 13059
rect 13557 13051 13591 13085
rect 13452 12899 13486 12933
rect 13653 13023 13687 13057
rect 13928 13015 13962 13049
rect 14142 13015 14176 13049
rect 14238 13015 14272 13049
rect 14379 13051 14413 13085
rect 14475 13051 14509 13085
rect 14637 13051 14671 13085
rect 13730 12915 13764 12949
rect 14547 12938 14581 12972
rect 14715 12938 14749 12972
rect 15162 13015 15196 13049
rect 15437 13023 15471 13057
rect 15533 13051 15567 13085
rect 15360 12915 15394 12949
rect 15677 13025 15711 13059
rect 15773 13073 15807 13107
rect 15638 12899 15672 12933
rect 15921 13013 15955 13047
rect 16017 13061 16051 13095
rect 16272 13067 16306 13101
rect 16374 13061 16408 13095
rect 16103 12925 16137 12959
rect 16533 12954 16567 12988
rect 16352 12899 16386 12933
rect 16740 13000 16774 13034
rect 16842 13015 16876 13049
rect 17015 13015 17049 13049
rect 17211 13015 17245 13049
rect 17415 13015 17449 13049
rect 17529 13015 17563 13049
rect 18091 13025 18125 13059
rect 18455 12989 18489 13023
rect 19195 13025 19229 13059
rect 19559 12989 19593 13023
rect 20011 13029 20045 13063
rect 20119 12989 20153 13023
rect 5295 12626 5329 12660
rect 5295 12558 5329 12592
rect 5015 12417 5049 12451
rect 5123 12377 5157 12411
rect 5295 12291 5329 12325
rect 5295 12223 5329 12257
rect 5395 12626 5429 12660
rect 5395 12558 5429 12592
rect 5947 12381 5981 12415
rect 6311 12417 6345 12451
rect 6847 12391 6881 12425
rect 6915 12391 6949 12425
rect 6983 12391 7017 12425
rect 7129 12391 7163 12425
rect 5395 12295 5429 12329
rect 5395 12227 5429 12261
rect 7377 12381 7411 12415
rect 7637 12417 7671 12451
rect 8063 12381 8097 12415
rect 8427 12417 8461 12451
rect 8963 12391 8997 12425
rect 9031 12391 9065 12425
rect 9099 12391 9133 12425
rect 9245 12391 9279 12425
rect 9493 12381 9527 12415
rect 9753 12417 9787 12451
rect 10067 12391 10101 12425
rect 10135 12391 10169 12425
rect 10203 12391 10237 12425
rect 10349 12391 10383 12425
rect 10554 12391 10588 12425
rect 10650 12391 10684 12425
rect 10959 12468 10993 12502
rect 10791 12355 10825 12389
rect 11127 12468 11161 12502
rect 10887 12355 10921 12389
rect 11049 12355 11083 12389
rect 11523 12468 11557 12502
rect 11691 12468 11725 12502
rect 11601 12355 11635 12389
rect 11763 12355 11797 12389
rect 11859 12355 11893 12389
rect 12000 12391 12034 12425
rect 12096 12391 12130 12425
rect 12827 12391 12861 12425
rect 12895 12391 12929 12425
rect 12963 12391 12997 12425
rect 13109 12391 13143 12425
rect 13313 12391 13347 12425
rect 13459 12391 13493 12425
rect 13527 12391 13561 12425
rect 13595 12391 13629 12425
rect 13817 12391 13851 12425
rect 13937 12404 13971 12438
rect 14137 12391 14171 12425
rect 14251 12391 14285 12425
rect 14455 12391 14489 12425
rect 14651 12391 14685 12425
rect 15100 12391 15134 12425
rect 15202 12406 15236 12440
rect 15590 12507 15624 12541
rect 15409 12452 15443 12486
rect 15839 12481 15873 12515
rect 15568 12345 15602 12379
rect 15670 12339 15704 12373
rect 15925 12345 15959 12379
rect 16021 12393 16055 12427
rect 16304 12507 16338 12541
rect 16169 12333 16203 12367
rect 16265 12381 16299 12415
rect 16582 12491 16616 12525
rect 16409 12355 16443 12389
rect 16505 12383 16539 12417
rect 16780 12391 16814 12425
rect 17085 12391 17119 12425
rect 17231 12391 17265 12425
rect 17299 12391 17333 12425
rect 17367 12391 17401 12425
rect 17831 12381 17865 12415
rect 17941 12381 17975 12415
rect 18049 12417 18083 12451
rect 18159 12417 18193 12451
rect 18643 12381 18677 12415
rect 19007 12417 19041 12451
rect 19477 12391 19511 12425
rect 19623 12391 19657 12425
rect 19691 12391 19725 12425
rect 19759 12391 19793 12425
rect 20011 12377 20045 12411
rect 20119 12417 20153 12451
rect 29830 6797 29998 6831
rect 30210 6797 30378 6831
rect 30468 6797 30636 6831
rect 30850 6797 31018 6831
rect 31108 6797 31276 6831
rect 31366 6797 31534 6831
rect 31750 6797 31918 6831
rect 32008 6797 32176 6831
rect 32266 6797 32434 6831
rect 32524 6797 32692 6831
rect 32782 6797 32950 6831
rect 33040 6797 33208 6831
rect 33298 6797 33466 6831
rect 33556 6797 33724 6831
rect 33814 6797 33982 6831
rect 34072 6797 34240 6831
rect 34450 6797 34618 6831
rect 29830 6069 29998 6103
rect 30210 6069 30378 6103
rect 30468 6069 30636 6103
rect 30850 6069 31018 6103
rect 31108 6069 31276 6103
rect 31366 6069 31534 6103
rect 31750 6069 31918 6103
rect 32008 6069 32176 6103
rect 32266 6069 32434 6103
rect 32524 6069 32692 6103
rect 32782 6069 32950 6103
rect 33040 6069 33208 6103
rect 33298 6069 33466 6103
rect 33556 6069 33724 6103
rect 33814 6069 33982 6103
rect 34072 6069 34240 6103
rect 34450 6069 34618 6103
rect 30072 5777 30106 5811
rect 30392 5777 30426 5811
rect 30792 5777 30826 5811
rect 31092 5777 31126 5811
rect 30072 5049 30106 5083
rect 30296 5049 30330 5083
rect 30488 5049 30522 5083
rect 30696 5049 30730 5083
rect 30888 5049 30922 5083
rect 31092 5049 31126 5083
rect 1482 4277 1516 4311
rect 1995 4270 2029 4304
rect 2187 4270 2221 4304
rect 2379 4270 2413 4304
rect 2571 4270 2605 4304
rect 2763 4270 2797 4304
rect 2955 4270 2989 4304
rect 3182 4277 3216 4311
rect 1682 3877 1716 3911
rect 1482 3149 1516 3183
rect 1682 3149 1716 3183
rect 1899 3142 1933 3176
rect 2091 3142 2125 3176
rect 2283 3142 2317 3176
rect 2475 3142 2509 3176
rect 2667 3142 2701 3176
rect 2859 3142 2893 3176
rect 3182 3149 3216 3183
rect 4782 4277 4816 4311
rect 5295 4270 5329 4304
rect 5487 4270 5521 4304
rect 5679 4270 5713 4304
rect 5871 4270 5905 4304
rect 6063 4270 6097 4304
rect 6255 4270 6289 4304
rect 6482 4277 6516 4311
rect 4982 3877 5016 3911
rect 4782 3149 4816 3183
rect 4982 3149 5016 3183
rect 5199 3142 5233 3176
rect 5391 3142 5425 3176
rect 5583 3142 5617 3176
rect 5775 3142 5809 3176
rect 5967 3142 6001 3176
rect 6159 3142 6193 3176
rect 6482 3149 6516 3183
rect 8082 4277 8116 4311
rect 8595 4270 8629 4304
rect 8787 4270 8821 4304
rect 8979 4270 9013 4304
rect 9171 4270 9205 4304
rect 9363 4270 9397 4304
rect 9555 4270 9589 4304
rect 9782 4277 9816 4311
rect 8282 3877 8316 3911
rect 8082 3149 8116 3183
rect 8282 3149 8316 3183
rect 8499 3142 8533 3176
rect 8691 3142 8725 3176
rect 8883 3142 8917 3176
rect 9075 3142 9109 3176
rect 9267 3142 9301 3176
rect 9459 3142 9493 3176
rect 9782 3149 9816 3183
rect 11382 4277 11416 4311
rect 11895 4270 11929 4304
rect 12087 4270 12121 4304
rect 12279 4270 12313 4304
rect 12471 4270 12505 4304
rect 12663 4270 12697 4304
rect 12855 4270 12889 4304
rect 13082 4277 13116 4311
rect 11582 3877 11616 3911
rect 11382 3149 11416 3183
rect 11582 3149 11616 3183
rect 11799 3142 11833 3176
rect 11991 3142 12025 3176
rect 12183 3142 12217 3176
rect 12375 3142 12409 3176
rect 12567 3142 12601 3176
rect 12759 3142 12793 3176
rect 13082 3149 13116 3183
rect 14982 4277 15016 4311
rect 15495 4270 15529 4304
rect 15687 4270 15721 4304
rect 15879 4270 15913 4304
rect 16071 4270 16105 4304
rect 16263 4270 16297 4304
rect 16455 4270 16489 4304
rect 16682 4277 16716 4311
rect 15182 3877 15216 3911
rect 14982 3149 15016 3183
rect 15182 3149 15216 3183
rect 15399 3142 15433 3176
rect 15591 3142 15625 3176
rect 15783 3142 15817 3176
rect 15975 3142 16009 3176
rect 16167 3142 16201 3176
rect 16359 3142 16393 3176
rect 16682 3149 16716 3183
rect 18482 4277 18516 4311
rect 18995 4270 19029 4304
rect 19187 4270 19221 4304
rect 19379 4270 19413 4304
rect 19571 4270 19605 4304
rect 19763 4270 19797 4304
rect 19955 4270 19989 4304
rect 20182 4277 20216 4311
rect 18682 3877 18716 3911
rect 18482 3149 18516 3183
rect 18682 3149 18716 3183
rect 18899 3142 18933 3176
rect 19091 3142 19125 3176
rect 19283 3142 19317 3176
rect 19475 3142 19509 3176
rect 19667 3142 19701 3176
rect 19859 3142 19893 3176
rect 20182 3149 20216 3183
rect 22182 4277 22216 4311
rect 22695 4270 22729 4304
rect 22887 4270 22921 4304
rect 23079 4270 23113 4304
rect 23271 4270 23305 4304
rect 23463 4270 23497 4304
rect 23655 4270 23689 4304
rect 23882 4277 23916 4311
rect 22382 3877 22416 3911
rect 22182 3149 22216 3183
rect 22382 3149 22416 3183
rect 22599 3142 22633 3176
rect 22791 3142 22825 3176
rect 22983 3142 23017 3176
rect 23175 3142 23209 3176
rect 23367 3142 23401 3176
rect 23559 3142 23593 3176
rect 23882 3149 23916 3183
rect 25982 4277 26016 4311
rect 26495 4270 26529 4304
rect 26687 4270 26721 4304
rect 26879 4270 26913 4304
rect 27071 4270 27105 4304
rect 27263 4270 27297 4304
rect 27455 4270 27489 4304
rect 27682 4277 27716 4311
rect 26182 3877 26216 3911
rect 25982 3149 26016 3183
rect 26182 3149 26216 3183
rect 26399 3142 26433 3176
rect 26591 3142 26625 3176
rect 26783 3142 26817 3176
rect 26975 3142 27009 3176
rect 27167 3142 27201 3176
rect 27359 3142 27393 3176
rect 27682 3149 27716 3183
rect 29934 4596 30102 4630
rect 30314 4596 30482 4630
rect 30714 4596 30882 4630
rect 31094 4596 31262 4630
rect 31352 4596 31520 4630
rect 31610 4596 31778 4630
rect 31868 4596 32036 4630
rect 32126 4596 32294 4630
rect 32384 4596 32552 4630
rect 32642 4596 32810 4630
rect 32900 4596 33068 4630
rect 33158 4596 33326 4630
rect 33534 4596 33702 4630
rect 29934 4286 30102 4320
rect 30314 4286 30482 4320
rect 30714 4286 30882 4320
rect 31094 4286 31262 4320
rect 31352 4286 31520 4320
rect 31610 4286 31778 4320
rect 31868 4286 32036 4320
rect 32126 4286 32294 4320
rect 32384 4286 32552 4320
rect 32642 4286 32810 4320
rect 32900 4286 33068 4320
rect 33158 4286 33326 4320
rect 33534 4286 33702 4320
rect 1486 2746 1520 2780
rect 1686 2746 1720 2780
rect 1999 2739 2033 2773
rect 2191 2739 2225 2773
rect 2383 2739 2417 2773
rect 2575 2739 2609 2773
rect 2767 2739 2801 2773
rect 2959 2739 2993 2773
rect 3166 2746 3200 2780
rect 1686 2436 1720 2470
rect 1486 1636 1520 1670
rect 1903 1629 1937 1663
rect 2095 1629 2129 1663
rect 2287 1629 2321 1663
rect 2479 1629 2513 1663
rect 2671 1629 2705 1663
rect 2863 1629 2897 1663
rect 3166 1636 3200 1670
rect 4786 2746 4820 2780
rect 4986 2746 5020 2780
rect 5299 2739 5333 2773
rect 5491 2739 5525 2773
rect 5683 2739 5717 2773
rect 5875 2739 5909 2773
rect 6067 2739 6101 2773
rect 6259 2739 6293 2773
rect 6466 2746 6500 2780
rect 4986 2436 5020 2470
rect 4786 1636 4820 1670
rect 5203 1629 5237 1663
rect 5395 1629 5429 1663
rect 5587 1629 5621 1663
rect 5779 1629 5813 1663
rect 5971 1629 6005 1663
rect 6163 1629 6197 1663
rect 6466 1636 6500 1670
rect 8086 2746 8120 2780
rect 8286 2746 8320 2780
rect 8599 2739 8633 2773
rect 8791 2739 8825 2773
rect 8983 2739 9017 2773
rect 9175 2739 9209 2773
rect 9367 2739 9401 2773
rect 9559 2739 9593 2773
rect 9766 2746 9800 2780
rect 8286 2436 8320 2470
rect 8086 1636 8120 1670
rect 8503 1629 8537 1663
rect 8695 1629 8729 1663
rect 8887 1629 8921 1663
rect 9079 1629 9113 1663
rect 9271 1629 9305 1663
rect 9463 1629 9497 1663
rect 9766 1636 9800 1670
rect 11386 2746 11420 2780
rect 11586 2746 11620 2780
rect 11899 2739 11933 2773
rect 12091 2739 12125 2773
rect 12283 2739 12317 2773
rect 12475 2739 12509 2773
rect 12667 2739 12701 2773
rect 12859 2739 12893 2773
rect 13066 2746 13100 2780
rect 11586 2436 11620 2470
rect 11386 1636 11420 1670
rect 11803 1629 11837 1663
rect 11995 1629 12029 1663
rect 12187 1629 12221 1663
rect 12379 1629 12413 1663
rect 12571 1629 12605 1663
rect 12763 1629 12797 1663
rect 13066 1636 13100 1670
rect 14986 2746 15020 2780
rect 15186 2746 15220 2780
rect 15499 2739 15533 2773
rect 15691 2739 15725 2773
rect 15883 2739 15917 2773
rect 16075 2739 16109 2773
rect 16267 2739 16301 2773
rect 16459 2739 16493 2773
rect 16666 2746 16700 2780
rect 15186 2436 15220 2470
rect 14986 1636 15020 1670
rect 15403 1629 15437 1663
rect 15595 1629 15629 1663
rect 15787 1629 15821 1663
rect 15979 1629 16013 1663
rect 16171 1629 16205 1663
rect 16363 1629 16397 1663
rect 16666 1636 16700 1670
rect 18486 2746 18520 2780
rect 18686 2746 18720 2780
rect 18999 2739 19033 2773
rect 19191 2739 19225 2773
rect 19383 2739 19417 2773
rect 19575 2739 19609 2773
rect 19767 2739 19801 2773
rect 19959 2739 19993 2773
rect 20166 2746 20200 2780
rect 18686 2436 18720 2470
rect 18486 1636 18520 1670
rect 18903 1629 18937 1663
rect 19095 1629 19129 1663
rect 19287 1629 19321 1663
rect 19479 1629 19513 1663
rect 19671 1629 19705 1663
rect 19863 1629 19897 1663
rect 20166 1636 20200 1670
rect 22186 2746 22220 2780
rect 22386 2746 22420 2780
rect 22699 2739 22733 2773
rect 22891 2739 22925 2773
rect 23083 2739 23117 2773
rect 23275 2739 23309 2773
rect 23467 2739 23501 2773
rect 23659 2739 23693 2773
rect 23866 2746 23900 2780
rect 22386 2436 22420 2470
rect 22186 1636 22220 1670
rect 22603 1629 22637 1663
rect 22795 1629 22829 1663
rect 22987 1629 23021 1663
rect 23179 1629 23213 1663
rect 23371 1629 23405 1663
rect 23563 1629 23597 1663
rect 23866 1636 23900 1670
rect 25986 2746 26020 2780
rect 26186 2746 26220 2780
rect 26499 2739 26533 2773
rect 26691 2739 26725 2773
rect 26883 2739 26917 2773
rect 27075 2739 27109 2773
rect 27267 2739 27301 2773
rect 27459 2739 27493 2773
rect 27666 2746 27700 2780
rect 26186 2436 26220 2470
rect 25986 1636 26020 1670
rect 26403 1629 26437 1663
rect 26595 1629 26629 1663
rect 26787 1629 26821 1663
rect 26979 1629 27013 1663
rect 27171 1629 27205 1663
rect 27363 1629 27397 1663
rect 27666 1636 27700 1670
<< xpolycontact >>
rect 25846 8662 25916 9094
rect 25846 7146 25916 7578
rect 26164 8662 26234 9094
rect 26164 7146 26234 7578
rect 26482 8662 26552 9094
rect 26482 7146 26552 7578
rect 26800 8662 26870 9094
rect 26800 7146 26870 7578
rect 27118 8662 27188 9094
rect 27118 7146 27188 7578
rect 27436 8662 27506 9094
rect 27436 7146 27506 7578
rect 27754 8662 27824 9094
rect 27754 7146 27824 7578
rect 28072 8662 28142 9094
rect 28072 7146 28142 7578
rect 3516 5438 3586 5870
rect 3516 4806 3586 5238
rect 6816 5342 6886 5774
rect 6816 4806 6886 5238
rect 10116 5482 10186 5914
rect 10116 4806 10186 5238
rect 13416 5762 13486 6194
rect 13416 4806 13486 5238
rect 17016 6322 17086 6754
rect 17016 4806 17086 5238
rect 20216 6322 20286 6754
rect 20216 4806 20286 5238
rect 20534 6322 20604 6754
rect 20534 4806 20604 5238
rect 23316 6322 23386 6754
rect 23316 4806 23386 5238
rect 23634 6322 23704 6754
rect 23634 4806 23704 5238
rect 23952 6322 24022 6754
rect 23952 4806 24022 5238
rect 24270 6322 24340 6754
rect 24270 4806 24340 5238
rect 25816 6322 25886 6754
rect 25816 4806 25886 5238
rect 26134 6322 26204 6754
rect 26134 4806 26204 5238
rect 26452 6322 26522 6754
rect 26452 4806 26522 5238
rect 26770 6322 26840 6754
rect 26770 4806 26840 5238
rect 27088 6322 27158 6754
rect 27088 4806 27158 5238
rect 27406 6322 27476 6754
rect 27406 4806 27476 5238
rect 27724 6322 27794 6754
rect 27724 4806 27794 5238
rect 28042 6322 28112 6754
rect 28042 4806 28112 5238
<< ppolyres >>
rect 3516 5238 3586 5438
<< xpolyres >>
rect 25846 7578 25916 8662
rect 26164 7578 26234 8662
rect 26482 7578 26552 8662
rect 26800 7578 26870 8662
rect 27118 7578 27188 8662
rect 27436 7578 27506 8662
rect 27754 7578 27824 8662
rect 28072 7578 28142 8662
rect 6816 5238 6886 5342
rect 10116 5238 10186 5482
rect 13416 5238 13486 5762
rect 17016 5238 17086 6322
rect 20216 5238 20286 6322
rect 20534 5238 20604 6322
rect 23316 5238 23386 6322
rect 23634 5238 23704 6322
rect 23952 5238 24022 6322
rect 24270 5238 24340 6322
rect 25816 5238 25886 6322
rect 26134 5238 26204 6322
rect 26452 5238 26522 6322
rect 26770 5238 26840 6322
rect 27088 5238 27158 6322
rect 27406 5238 27476 6322
rect 27724 5238 27794 6322
rect 28042 5238 28112 6322
<< rmp >>
rect 5245 12408 5341 12417
rect 5383 12408 5479 12417
<< locali >>
rect 4948 27391 4977 27425
rect 5011 27391 5069 27425
rect 5103 27391 5161 27425
rect 5195 27391 5253 27425
rect 5287 27391 5345 27425
rect 5379 27391 5437 27425
rect 5471 27391 5529 27425
rect 5563 27391 5621 27425
rect 5655 27391 5713 27425
rect 5747 27391 5805 27425
rect 5839 27391 5897 27425
rect 5931 27391 5989 27425
rect 6023 27391 6081 27425
rect 6115 27391 6173 27425
rect 6207 27391 6265 27425
rect 6299 27391 6357 27425
rect 6391 27391 6449 27425
rect 6483 27391 6541 27425
rect 6575 27391 6633 27425
rect 6667 27391 6725 27425
rect 6759 27391 6817 27425
rect 6851 27391 6909 27425
rect 6943 27391 7001 27425
rect 7035 27391 7093 27425
rect 7127 27391 7185 27425
rect 7219 27391 7277 27425
rect 7311 27391 7369 27425
rect 7403 27391 7461 27425
rect 7495 27391 7553 27425
rect 7587 27391 7645 27425
rect 7679 27391 7737 27425
rect 7771 27391 7829 27425
rect 7863 27391 7921 27425
rect 7955 27391 8013 27425
rect 8047 27391 8105 27425
rect 8139 27391 8197 27425
rect 8231 27391 8289 27425
rect 8323 27391 8381 27425
rect 8415 27391 8473 27425
rect 8507 27391 8565 27425
rect 8599 27391 8657 27425
rect 8691 27391 8749 27425
rect 8783 27391 8841 27425
rect 8875 27391 8933 27425
rect 8967 27391 9025 27425
rect 9059 27391 9117 27425
rect 9151 27391 9209 27425
rect 9243 27391 9301 27425
rect 9335 27391 9393 27425
rect 9427 27391 9485 27425
rect 9519 27391 9577 27425
rect 9611 27391 9669 27425
rect 9703 27391 9761 27425
rect 9795 27391 9853 27425
rect 9887 27391 9945 27425
rect 9979 27391 10037 27425
rect 10071 27391 10129 27425
rect 10163 27391 10221 27425
rect 10255 27391 10313 27425
rect 10347 27391 10405 27425
rect 10439 27391 10497 27425
rect 10531 27391 10589 27425
rect 10623 27391 10681 27425
rect 10715 27391 10773 27425
rect 10807 27391 10865 27425
rect 10899 27391 10957 27425
rect 10991 27391 11049 27425
rect 11083 27391 11141 27425
rect 11175 27391 11233 27425
rect 11267 27391 11325 27425
rect 11359 27391 11417 27425
rect 11451 27391 11509 27425
rect 11543 27391 11601 27425
rect 11635 27391 11693 27425
rect 11727 27391 11785 27425
rect 11819 27391 11877 27425
rect 11911 27391 11969 27425
rect 12003 27391 12061 27425
rect 12095 27391 12153 27425
rect 12187 27391 12245 27425
rect 12279 27391 12337 27425
rect 12371 27391 12429 27425
rect 12463 27391 12521 27425
rect 12555 27391 12613 27425
rect 12647 27391 12705 27425
rect 12739 27391 12797 27425
rect 12831 27391 12889 27425
rect 12923 27391 12981 27425
rect 13015 27391 13073 27425
rect 13107 27391 13165 27425
rect 13199 27391 13257 27425
rect 13291 27391 13349 27425
rect 13383 27391 13441 27425
rect 13475 27391 13533 27425
rect 13567 27391 13625 27425
rect 13659 27391 13717 27425
rect 13751 27391 13809 27425
rect 13843 27391 13901 27425
rect 13935 27391 13993 27425
rect 14027 27391 14085 27425
rect 14119 27391 14177 27425
rect 14211 27391 14269 27425
rect 14303 27391 14361 27425
rect 14395 27391 14453 27425
rect 14487 27391 14545 27425
rect 14579 27391 14637 27425
rect 14671 27391 14729 27425
rect 14763 27391 14821 27425
rect 14855 27391 14913 27425
rect 14947 27391 15005 27425
rect 15039 27391 15097 27425
rect 15131 27391 15189 27425
rect 15223 27391 15281 27425
rect 15315 27391 15373 27425
rect 15407 27391 15465 27425
rect 15499 27391 15557 27425
rect 15591 27391 15649 27425
rect 15683 27391 15741 27425
rect 15775 27391 15833 27425
rect 15867 27391 15925 27425
rect 15959 27391 16017 27425
rect 16051 27391 16109 27425
rect 16143 27391 16201 27425
rect 16235 27391 16293 27425
rect 16327 27391 16385 27425
rect 16419 27391 16477 27425
rect 16511 27391 16569 27425
rect 16603 27391 16661 27425
rect 16695 27391 16753 27425
rect 16787 27391 16845 27425
rect 16879 27391 16937 27425
rect 16971 27391 17029 27425
rect 17063 27391 17121 27425
rect 17155 27391 17213 27425
rect 17247 27391 17305 27425
rect 17339 27391 17397 27425
rect 17431 27391 17489 27425
rect 17523 27391 17581 27425
rect 17615 27391 17673 27425
rect 17707 27391 17765 27425
rect 17799 27391 17857 27425
rect 17891 27391 17949 27425
rect 17983 27391 18041 27425
rect 18075 27391 18133 27425
rect 18167 27391 18225 27425
rect 18259 27391 18317 27425
rect 18351 27391 18409 27425
rect 18443 27391 18501 27425
rect 18535 27391 18593 27425
rect 18627 27391 18685 27425
rect 18719 27391 18777 27425
rect 18811 27391 18869 27425
rect 18903 27391 18961 27425
rect 18995 27391 19053 27425
rect 19087 27391 19145 27425
rect 19179 27391 19237 27425
rect 19271 27391 19329 27425
rect 19363 27391 19421 27425
rect 19455 27391 19513 27425
rect 19547 27391 19605 27425
rect 19639 27391 19697 27425
rect 19731 27391 19789 27425
rect 19823 27391 19881 27425
rect 19915 27391 19973 27425
rect 20007 27391 20065 27425
rect 20099 27391 20157 27425
rect 20191 27391 20220 27425
rect 4965 27328 5207 27391
rect 4965 27294 4983 27328
rect 5017 27294 5155 27328
rect 5189 27294 5207 27328
rect 4965 27241 5207 27294
rect 5241 27328 5483 27391
rect 5241 27294 5259 27328
rect 5293 27294 5431 27328
rect 5465 27294 5483 27328
rect 5529 27345 5585 27391
rect 5529 27311 5542 27345
rect 5576 27311 5585 27345
rect 5706 27345 5757 27391
rect 5529 27295 5585 27311
rect 5619 27323 5671 27339
rect 5241 27241 5483 27294
rect 5619 27289 5628 27323
rect 5662 27289 5671 27323
rect 5706 27311 5714 27345
rect 5748 27311 5757 27345
rect 5886 27345 5941 27391
rect 5706 27295 5757 27311
rect 5791 27323 5850 27339
rect 5619 27261 5671 27289
rect 5791 27289 5800 27323
rect 5834 27289 5850 27323
rect 5886 27311 5897 27345
rect 5931 27311 5941 27345
rect 5886 27295 5941 27311
rect 5975 27341 6035 27357
rect 5975 27307 5983 27341
rect 6017 27307 6035 27341
rect 5975 27291 6035 27307
rect 5791 27261 5850 27289
rect 4965 27167 5069 27241
rect 4965 27133 5015 27167
rect 5049 27133 5069 27167
rect 5103 27173 5123 27207
rect 5157 27173 5207 27207
rect 5103 27099 5207 27173
rect 4965 27052 5207 27099
rect 4965 27018 4983 27052
rect 5017 27018 5155 27052
rect 5189 27018 5207 27052
rect 4965 26957 5207 27018
rect 4965 26923 4983 26957
rect 5017 26923 5155 26957
rect 5189 26923 5207 26957
rect 4965 26881 5207 26923
rect 5241 27173 5291 27207
rect 5325 27173 5345 27207
rect 5241 27099 5345 27173
rect 5379 27167 5483 27241
rect 5379 27133 5399 27167
rect 5433 27133 5483 27167
rect 5520 27227 5850 27261
rect 5897 27255 5967 27257
rect 5520 27125 5601 27227
rect 5931 27221 5967 27255
rect 5897 27193 5967 27221
rect 5635 27159 5651 27193
rect 5685 27159 5719 27193
rect 5753 27159 5787 27193
rect 5821 27159 5863 27193
rect 5520 27101 5671 27125
rect 5241 27052 5483 27099
rect 5520 27091 5629 27101
rect 5619 27067 5629 27091
rect 5663 27067 5671 27101
rect 5829 27109 5863 27159
rect 5897 27159 5933 27193
rect 5897 27143 5967 27159
rect 6001 27109 6035 27291
rect 6162 27330 7231 27391
rect 6162 27296 6179 27330
rect 6213 27296 7179 27330
rect 7213 27296 7231 27330
rect 6162 27282 7231 27296
rect 7265 27297 7323 27391
rect 5829 27087 6035 27109
rect 5829 27075 5983 27087
rect 5241 27018 5259 27052
rect 5293 27018 5431 27052
rect 5465 27018 5483 27052
rect 5241 26957 5483 27018
rect 5241 26923 5259 26957
rect 5293 26923 5431 26957
rect 5465 26923 5483 26957
rect 5241 26881 5483 26923
rect 5528 27039 5585 27055
rect 5528 27005 5543 27039
rect 5577 27005 5585 27039
rect 5528 26971 5585 27005
rect 5528 26937 5543 26971
rect 5577 26937 5585 26971
rect 5528 26881 5585 26937
rect 5619 27041 5671 27067
rect 5973 27053 5983 27075
rect 6017 27053 6035 27087
rect 5619 27033 5843 27041
rect 5619 26999 5629 27033
rect 5663 27007 5843 27033
rect 5663 26999 5671 27007
rect 5619 26965 5671 26999
rect 5791 26992 5843 27007
rect 5619 26931 5629 26965
rect 5663 26931 5671 26965
rect 5619 26915 5671 26931
rect 5706 26957 5757 26973
rect 5706 26923 5715 26957
rect 5749 26923 5757 26957
rect 5706 26881 5757 26923
rect 5791 26958 5801 26992
rect 5835 26983 5843 26992
rect 5791 26949 5805 26958
rect 5839 26949 5843 26983
rect 5791 26915 5843 26949
rect 5877 27025 5939 27041
rect 5877 26991 5897 27025
rect 5931 26991 5939 27025
rect 5877 26957 5939 26991
rect 5877 26923 5897 26957
rect 5931 26923 5939 26957
rect 5877 26881 5939 26923
rect 5973 26965 6035 27053
rect 6480 27203 6550 27218
rect 6480 27169 6499 27203
rect 6533 27169 6550 27203
rect 6480 26968 6550 27169
rect 6846 27167 6914 27282
rect 7265 27263 7277 27297
rect 7311 27263 7323 27297
rect 7265 27246 7323 27263
rect 7357 27328 7599 27391
rect 7357 27294 7375 27328
rect 7409 27294 7547 27328
rect 7581 27294 7599 27328
rect 7357 27241 7599 27294
rect 7634 27330 8703 27391
rect 7634 27296 7651 27330
rect 7685 27296 8651 27330
rect 8685 27296 8703 27330
rect 7634 27282 8703 27296
rect 8738 27330 9807 27391
rect 8738 27296 8755 27330
rect 8789 27296 9755 27330
rect 9789 27296 9807 27330
rect 8738 27282 9807 27296
rect 9841 27297 9899 27391
rect 6846 27133 6863 27167
rect 6897 27133 6914 27167
rect 6846 27116 6914 27133
rect 7357 27173 7407 27207
rect 7441 27173 7461 27207
rect 7265 27079 7323 27114
rect 7265 27045 7277 27079
rect 7311 27045 7323 27079
rect 7265 26986 7323 27045
rect 5973 26931 5983 26965
rect 6017 26931 6035 26965
rect 5973 26915 6035 26931
rect 6162 26957 7231 26968
rect 6162 26923 6179 26957
rect 6213 26923 7179 26957
rect 7213 26923 7231 26957
rect 6162 26881 7231 26923
rect 7265 26952 7277 26986
rect 7311 26952 7323 26986
rect 7265 26881 7323 26952
rect 7357 27099 7461 27173
rect 7495 27167 7599 27241
rect 7495 27133 7515 27167
rect 7549 27133 7599 27167
rect 7952 27203 8022 27218
rect 7952 27169 7971 27203
rect 8005 27169 8022 27203
rect 7357 27052 7599 27099
rect 7357 27018 7375 27052
rect 7409 27018 7547 27052
rect 7581 27018 7599 27052
rect 7357 26957 7599 27018
rect 7952 26968 8022 27169
rect 8318 27167 8386 27282
rect 8318 27133 8335 27167
rect 8369 27133 8386 27167
rect 8318 27116 8386 27133
rect 9056 27203 9126 27218
rect 9056 27169 9075 27203
rect 9109 27169 9126 27203
rect 9056 26968 9126 27169
rect 9422 27167 9490 27282
rect 9841 27263 9853 27297
rect 9887 27263 9899 27297
rect 9841 27246 9899 27263
rect 10135 27336 10169 27357
rect 10205 27349 10271 27391
rect 10205 27315 10221 27349
rect 10255 27315 10271 27349
rect 10307 27319 10359 27357
rect 10135 27281 10169 27302
rect 10341 27285 10359 27319
rect 10135 27247 10268 27281
rect 10307 27256 10359 27285
rect 9422 27133 9439 27167
rect 9473 27133 9490 27167
rect 10121 27193 10189 27211
rect 10121 27187 10137 27193
rect 10121 27153 10129 27187
rect 10171 27159 10189 27193
rect 10163 27153 10189 27159
rect 10121 27137 10189 27153
rect 10234 27196 10268 27247
rect 10234 27180 10289 27196
rect 10234 27146 10255 27180
rect 9422 27116 9490 27133
rect 10234 27130 10289 27146
rect 9841 27079 9899 27114
rect 10234 27101 10268 27130
rect 9841 27045 9853 27079
rect 9887 27045 9899 27079
rect 9841 26986 9899 27045
rect 7357 26923 7375 26957
rect 7409 26923 7547 26957
rect 7581 26923 7599 26957
rect 7357 26881 7599 26923
rect 7634 26957 8703 26968
rect 7634 26923 7651 26957
rect 7685 26923 8651 26957
rect 8685 26923 8703 26957
rect 7634 26881 8703 26923
rect 8738 26957 9807 26968
rect 8738 26923 8755 26957
rect 8789 26923 9755 26957
rect 9789 26923 9807 26957
rect 8738 26881 9807 26923
rect 9841 26952 9853 26986
rect 9887 26952 9899 26986
rect 9841 26881 9899 26952
rect 10133 27067 10268 27101
rect 10323 27096 10359 27256
rect 10577 27330 11279 27391
rect 10577 27296 10595 27330
rect 10629 27296 11227 27330
rect 11261 27296 11279 27330
rect 10577 27237 11279 27296
rect 11314 27330 12383 27391
rect 11314 27296 11331 27330
rect 11365 27296 12331 27330
rect 12365 27296 12383 27330
rect 11314 27282 12383 27296
rect 12417 27297 12475 27391
rect 10133 27033 10169 27067
rect 10305 27046 10359 27096
rect 10133 26999 10135 27033
rect 10133 26965 10169 26999
rect 10133 26931 10135 26965
rect 10133 26915 10169 26931
rect 10205 26999 10221 27033
rect 10255 26999 10271 27033
rect 10205 26965 10271 26999
rect 10205 26931 10221 26965
rect 10255 26931 10271 26965
rect 10205 26881 10271 26931
rect 10305 27012 10307 27046
rect 10341 27012 10359 27046
rect 10305 26983 10359 27012
rect 10305 26965 10313 26983
rect 10305 26931 10307 26965
rect 10347 26949 10359 26983
rect 10341 26931 10359 26949
rect 10305 26915 10359 26931
rect 10577 27169 10655 27203
rect 10689 27169 10758 27203
rect 10792 27169 10861 27203
rect 10895 27169 10915 27203
rect 10577 27099 10915 27169
rect 10949 27167 11279 27237
rect 10949 27133 10969 27167
rect 11003 27133 11068 27167
rect 11102 27133 11167 27167
rect 11201 27133 11279 27167
rect 11632 27203 11702 27218
rect 11632 27169 11651 27203
rect 11685 27169 11702 27203
rect 10577 27059 11279 27099
rect 10577 27025 10595 27059
rect 10629 27025 11227 27059
rect 11261 27025 11279 27059
rect 10577 26957 11279 27025
rect 11632 26968 11702 27169
rect 11998 27167 12066 27282
rect 12417 27263 12429 27297
rect 12463 27263 12475 27297
rect 12417 27246 12475 27263
rect 12509 27328 12751 27391
rect 12509 27294 12527 27328
rect 12561 27294 12699 27328
rect 12733 27294 12751 27328
rect 12509 27241 12751 27294
rect 12786 27330 13855 27391
rect 12786 27296 12803 27330
rect 12837 27296 13803 27330
rect 13837 27296 13855 27330
rect 12786 27282 13855 27296
rect 13890 27330 14959 27391
rect 13890 27296 13907 27330
rect 13941 27296 14907 27330
rect 14941 27296 14959 27330
rect 13890 27282 14959 27296
rect 14993 27297 15051 27391
rect 11998 27133 12015 27167
rect 12049 27133 12066 27167
rect 11998 27116 12066 27133
rect 12509 27173 12559 27207
rect 12593 27173 12613 27207
rect 12417 27079 12475 27114
rect 12417 27045 12429 27079
rect 12463 27045 12475 27079
rect 12417 26986 12475 27045
rect 10577 26923 10595 26957
rect 10629 26923 11227 26957
rect 11261 26923 11279 26957
rect 10577 26881 11279 26923
rect 11314 26957 12383 26968
rect 11314 26923 11331 26957
rect 11365 26923 12331 26957
rect 12365 26923 12383 26957
rect 11314 26881 12383 26923
rect 12417 26952 12429 26986
rect 12463 26952 12475 26986
rect 12417 26881 12475 26952
rect 12509 27099 12613 27173
rect 12647 27167 12751 27241
rect 12647 27133 12667 27167
rect 12701 27133 12751 27167
rect 13104 27203 13174 27218
rect 13104 27169 13123 27203
rect 13157 27169 13174 27203
rect 12509 27052 12751 27099
rect 12509 27018 12527 27052
rect 12561 27018 12699 27052
rect 12733 27018 12751 27052
rect 12509 26957 12751 27018
rect 13104 26968 13174 27169
rect 13470 27167 13538 27282
rect 13470 27133 13487 27167
rect 13521 27133 13538 27167
rect 13470 27116 13538 27133
rect 14208 27203 14278 27218
rect 14208 27169 14227 27203
rect 14261 27169 14278 27203
rect 14208 26968 14278 27169
rect 14574 27167 14642 27282
rect 14993 27263 15005 27297
rect 15039 27263 15051 27297
rect 14993 27246 15051 27263
rect 15085 27328 15327 27391
rect 15085 27294 15103 27328
rect 15137 27294 15275 27328
rect 15309 27294 15327 27328
rect 15085 27241 15327 27294
rect 15362 27330 16431 27391
rect 15362 27296 15379 27330
rect 15413 27296 16379 27330
rect 16413 27296 16431 27330
rect 15362 27282 16431 27296
rect 16466 27330 17535 27391
rect 16466 27296 16483 27330
rect 16517 27296 17483 27330
rect 17517 27296 17535 27330
rect 16466 27282 17535 27296
rect 17569 27297 17627 27391
rect 14574 27133 14591 27167
rect 14625 27133 14642 27167
rect 14574 27116 14642 27133
rect 15085 27173 15135 27207
rect 15169 27173 15189 27207
rect 14993 27079 15051 27114
rect 14993 27045 15005 27079
rect 15039 27045 15051 27079
rect 14993 26986 15051 27045
rect 12509 26923 12527 26957
rect 12561 26923 12699 26957
rect 12733 26923 12751 26957
rect 12509 26881 12751 26923
rect 12786 26957 13855 26968
rect 12786 26923 12803 26957
rect 12837 26923 13803 26957
rect 13837 26923 13855 26957
rect 12786 26881 13855 26923
rect 13890 26957 14959 26968
rect 13890 26923 13907 26957
rect 13941 26923 14907 26957
rect 14941 26923 14959 26957
rect 13890 26881 14959 26923
rect 14993 26952 15005 26986
rect 15039 26952 15051 26986
rect 14993 26881 15051 26952
rect 15085 27099 15189 27173
rect 15223 27167 15327 27241
rect 15223 27133 15243 27167
rect 15277 27133 15327 27167
rect 15680 27203 15750 27218
rect 15680 27169 15699 27203
rect 15733 27169 15750 27203
rect 15085 27052 15327 27099
rect 15085 27018 15103 27052
rect 15137 27018 15275 27052
rect 15309 27018 15327 27052
rect 15085 26957 15327 27018
rect 15680 26968 15750 27169
rect 16046 27167 16114 27282
rect 16046 27133 16063 27167
rect 16097 27133 16114 27167
rect 16046 27116 16114 27133
rect 16784 27203 16854 27218
rect 16784 27169 16803 27203
rect 16837 27169 16854 27203
rect 16784 26968 16854 27169
rect 17150 27167 17218 27282
rect 17569 27263 17581 27297
rect 17615 27263 17627 27297
rect 17569 27246 17627 27263
rect 17753 27330 18455 27391
rect 17753 27296 17771 27330
rect 17805 27296 18403 27330
rect 18437 27296 18455 27330
rect 17753 27237 18455 27296
rect 18501 27345 18557 27391
rect 18501 27311 18514 27345
rect 18548 27311 18557 27345
rect 18678 27345 18729 27391
rect 18501 27295 18557 27311
rect 18591 27323 18643 27339
rect 18591 27289 18600 27323
rect 18634 27289 18643 27323
rect 18678 27311 18686 27345
rect 18720 27311 18729 27345
rect 18858 27345 18913 27391
rect 18678 27295 18729 27311
rect 18763 27323 18822 27339
rect 18591 27261 18643 27289
rect 18763 27289 18772 27323
rect 18806 27289 18822 27323
rect 18858 27311 18869 27345
rect 18903 27311 18913 27345
rect 18858 27295 18913 27311
rect 18947 27341 19007 27357
rect 18947 27307 18955 27341
rect 18989 27307 19007 27341
rect 18947 27291 19007 27307
rect 18763 27261 18822 27289
rect 17150 27133 17167 27167
rect 17201 27133 17218 27167
rect 17150 27116 17218 27133
rect 17753 27169 17831 27203
rect 17865 27169 17934 27203
rect 17968 27169 18037 27203
rect 18071 27169 18091 27203
rect 17569 27079 17627 27114
rect 17569 27045 17581 27079
rect 17615 27045 17627 27079
rect 17569 26986 17627 27045
rect 15085 26923 15103 26957
rect 15137 26923 15275 26957
rect 15309 26923 15327 26957
rect 15085 26881 15327 26923
rect 15362 26957 16431 26968
rect 15362 26923 15379 26957
rect 15413 26923 16379 26957
rect 16413 26923 16431 26957
rect 15362 26881 16431 26923
rect 16466 26957 17535 26968
rect 16466 26923 16483 26957
rect 16517 26923 17483 26957
rect 17517 26923 17535 26957
rect 16466 26881 17535 26923
rect 17569 26952 17581 26986
rect 17615 26952 17627 26986
rect 17569 26881 17627 26952
rect 17753 27099 18091 27169
rect 18125 27167 18455 27237
rect 18125 27133 18145 27167
rect 18179 27133 18244 27167
rect 18278 27133 18343 27167
rect 18377 27133 18455 27167
rect 18492 27227 18822 27261
rect 18869 27255 18939 27257
rect 18492 27125 18573 27227
rect 18903 27221 18939 27255
rect 18869 27193 18939 27221
rect 18607 27159 18623 27193
rect 18657 27159 18691 27193
rect 18725 27159 18759 27193
rect 18793 27159 18835 27193
rect 18492 27101 18643 27125
rect 17753 27059 18455 27099
rect 18492 27091 18601 27101
rect 17753 27025 17771 27059
rect 17805 27025 18403 27059
rect 18437 27025 18455 27059
rect 18591 27067 18601 27091
rect 18635 27067 18643 27101
rect 18801 27109 18835 27159
rect 18869 27159 18905 27193
rect 18869 27143 18939 27159
rect 18973 27109 19007 27291
rect 19225 27330 19927 27391
rect 19225 27296 19243 27330
rect 19277 27296 19875 27330
rect 19909 27296 19927 27330
rect 19225 27237 19927 27296
rect 19961 27328 20203 27391
rect 19961 27294 19979 27328
rect 20013 27294 20151 27328
rect 20185 27294 20203 27328
rect 19961 27241 20203 27294
rect 18801 27087 19007 27109
rect 18801 27075 18955 27087
rect 17753 26957 18455 27025
rect 17753 26923 17771 26957
rect 17805 26923 18403 26957
rect 18437 26923 18455 26957
rect 17753 26881 18455 26923
rect 18500 27039 18557 27055
rect 18500 27005 18515 27039
rect 18549 27005 18557 27039
rect 18500 26971 18557 27005
rect 18500 26937 18515 26971
rect 18549 26937 18557 26971
rect 18500 26881 18557 26937
rect 18591 27041 18643 27067
rect 18945 27053 18955 27075
rect 18989 27053 19007 27087
rect 18591 27033 18815 27041
rect 18591 26999 18601 27033
rect 18635 27007 18815 27033
rect 18635 26999 18643 27007
rect 18591 26965 18643 26999
rect 18763 26992 18815 27007
rect 18591 26931 18601 26965
rect 18635 26931 18643 26965
rect 18591 26915 18643 26931
rect 18678 26957 18729 26973
rect 18678 26923 18687 26957
rect 18721 26923 18729 26957
rect 18678 26881 18729 26923
rect 18763 26958 18773 26992
rect 18807 26983 18815 26992
rect 18763 26949 18777 26958
rect 18811 26949 18815 26983
rect 18763 26915 18815 26949
rect 18849 27025 18911 27041
rect 18849 26991 18869 27025
rect 18903 26991 18911 27025
rect 18849 26957 18911 26991
rect 18849 26923 18869 26957
rect 18903 26923 18911 26957
rect 18849 26881 18911 26923
rect 18945 26965 19007 27053
rect 18945 26931 18955 26965
rect 18989 26931 19007 26965
rect 18945 26915 19007 26931
rect 19225 27169 19303 27203
rect 19337 27169 19406 27203
rect 19440 27169 19509 27203
rect 19543 27169 19563 27203
rect 19225 27099 19563 27169
rect 19597 27167 19927 27237
rect 19597 27133 19617 27167
rect 19651 27133 19716 27167
rect 19750 27133 19815 27167
rect 19849 27133 19927 27167
rect 19961 27173 20011 27207
rect 20045 27173 20065 27207
rect 19961 27099 20065 27173
rect 20099 27167 20203 27241
rect 20099 27133 20119 27167
rect 20153 27133 20203 27167
rect 19225 27059 19927 27099
rect 19225 27025 19243 27059
rect 19277 27025 19875 27059
rect 19909 27025 19927 27059
rect 19225 26957 19927 27025
rect 19225 26923 19243 26957
rect 19277 26923 19875 26957
rect 19909 26923 19927 26957
rect 19225 26881 19927 26923
rect 19961 27052 20203 27099
rect 19961 27018 19979 27052
rect 20013 27018 20151 27052
rect 20185 27018 20203 27052
rect 19961 26957 20203 27018
rect 19961 26923 19979 26957
rect 20013 26923 20151 26957
rect 20185 26923 20203 26957
rect 19961 26881 20203 26923
rect 4948 26847 4977 26881
rect 5011 26847 5069 26881
rect 5103 26847 5161 26881
rect 5195 26847 5253 26881
rect 5287 26847 5345 26881
rect 5379 26847 5437 26881
rect 5471 26847 5529 26881
rect 5563 26847 5621 26881
rect 5655 26847 5713 26881
rect 5747 26847 5805 26881
rect 5839 26847 5897 26881
rect 5931 26847 5989 26881
rect 6023 26847 6081 26881
rect 6115 26847 6173 26881
rect 6207 26847 6265 26881
rect 6299 26847 6357 26881
rect 6391 26847 6449 26881
rect 6483 26847 6541 26881
rect 6575 26847 6633 26881
rect 6667 26847 6725 26881
rect 6759 26847 6817 26881
rect 6851 26847 6909 26881
rect 6943 26847 7001 26881
rect 7035 26847 7093 26881
rect 7127 26847 7185 26881
rect 7219 26847 7277 26881
rect 7311 26847 7369 26881
rect 7403 26847 7461 26881
rect 7495 26847 7553 26881
rect 7587 26847 7645 26881
rect 7679 26847 7737 26881
rect 7771 26847 7829 26881
rect 7863 26847 7921 26881
rect 7955 26847 8013 26881
rect 8047 26847 8105 26881
rect 8139 26847 8197 26881
rect 8231 26847 8289 26881
rect 8323 26847 8381 26881
rect 8415 26847 8473 26881
rect 8507 26847 8565 26881
rect 8599 26847 8657 26881
rect 8691 26847 8749 26881
rect 8783 26847 8841 26881
rect 8875 26847 8933 26881
rect 8967 26847 9025 26881
rect 9059 26847 9117 26881
rect 9151 26847 9209 26881
rect 9243 26847 9301 26881
rect 9335 26847 9393 26881
rect 9427 26847 9485 26881
rect 9519 26847 9577 26881
rect 9611 26847 9669 26881
rect 9703 26847 9761 26881
rect 9795 26847 9853 26881
rect 9887 26847 9945 26881
rect 9979 26847 10037 26881
rect 10071 26847 10129 26881
rect 10163 26847 10221 26881
rect 10255 26847 10313 26881
rect 10347 26847 10405 26881
rect 10439 26847 10497 26881
rect 10531 26847 10589 26881
rect 10623 26847 10681 26881
rect 10715 26847 10773 26881
rect 10807 26847 10865 26881
rect 10899 26847 10957 26881
rect 10991 26847 11049 26881
rect 11083 26847 11141 26881
rect 11175 26847 11233 26881
rect 11267 26847 11325 26881
rect 11359 26847 11417 26881
rect 11451 26847 11509 26881
rect 11543 26847 11601 26881
rect 11635 26847 11693 26881
rect 11727 26847 11785 26881
rect 11819 26847 11877 26881
rect 11911 26847 11969 26881
rect 12003 26847 12061 26881
rect 12095 26847 12153 26881
rect 12187 26847 12245 26881
rect 12279 26847 12337 26881
rect 12371 26847 12429 26881
rect 12463 26847 12521 26881
rect 12555 26847 12613 26881
rect 12647 26847 12705 26881
rect 12739 26847 12797 26881
rect 12831 26847 12889 26881
rect 12923 26847 12981 26881
rect 13015 26847 13073 26881
rect 13107 26847 13165 26881
rect 13199 26847 13257 26881
rect 13291 26847 13349 26881
rect 13383 26847 13441 26881
rect 13475 26847 13533 26881
rect 13567 26847 13625 26881
rect 13659 26847 13717 26881
rect 13751 26847 13809 26881
rect 13843 26847 13901 26881
rect 13935 26847 13993 26881
rect 14027 26847 14085 26881
rect 14119 26847 14177 26881
rect 14211 26847 14269 26881
rect 14303 26847 14361 26881
rect 14395 26847 14453 26881
rect 14487 26847 14545 26881
rect 14579 26847 14637 26881
rect 14671 26847 14729 26881
rect 14763 26847 14821 26881
rect 14855 26847 14913 26881
rect 14947 26847 15005 26881
rect 15039 26847 15097 26881
rect 15131 26847 15189 26881
rect 15223 26847 15281 26881
rect 15315 26847 15373 26881
rect 15407 26847 15465 26881
rect 15499 26847 15557 26881
rect 15591 26847 15649 26881
rect 15683 26847 15741 26881
rect 15775 26847 15833 26881
rect 15867 26847 15925 26881
rect 15959 26847 16017 26881
rect 16051 26847 16109 26881
rect 16143 26847 16201 26881
rect 16235 26847 16293 26881
rect 16327 26847 16385 26881
rect 16419 26847 16477 26881
rect 16511 26847 16569 26881
rect 16603 26847 16661 26881
rect 16695 26847 16753 26881
rect 16787 26847 16845 26881
rect 16879 26847 16937 26881
rect 16971 26847 17029 26881
rect 17063 26847 17121 26881
rect 17155 26847 17213 26881
rect 17247 26847 17305 26881
rect 17339 26847 17397 26881
rect 17431 26847 17489 26881
rect 17523 26847 17581 26881
rect 17615 26847 17673 26881
rect 17707 26847 17765 26881
rect 17799 26847 17857 26881
rect 17891 26847 17949 26881
rect 17983 26847 18041 26881
rect 18075 26847 18133 26881
rect 18167 26847 18225 26881
rect 18259 26847 18317 26881
rect 18351 26847 18409 26881
rect 18443 26847 18501 26881
rect 18535 26847 18593 26881
rect 18627 26847 18685 26881
rect 18719 26847 18777 26881
rect 18811 26847 18869 26881
rect 18903 26847 18961 26881
rect 18995 26847 19053 26881
rect 19087 26847 19145 26881
rect 19179 26847 19237 26881
rect 19271 26847 19329 26881
rect 19363 26847 19421 26881
rect 19455 26847 19513 26881
rect 19547 26847 19605 26881
rect 19639 26847 19697 26881
rect 19731 26847 19789 26881
rect 19823 26847 19881 26881
rect 19915 26847 19973 26881
rect 20007 26847 20065 26881
rect 20099 26847 20157 26881
rect 20191 26847 20220 26881
rect 4965 26805 5207 26847
rect 4965 26771 4983 26805
rect 5017 26771 5155 26805
rect 5189 26771 5207 26805
rect 4965 26710 5207 26771
rect 4965 26676 4983 26710
rect 5017 26676 5155 26710
rect 5189 26676 5207 26710
rect 4965 26629 5207 26676
rect 4965 26561 5015 26595
rect 5049 26561 5069 26595
rect 4965 26487 5069 26561
rect 5103 26555 5207 26629
rect 5103 26521 5123 26555
rect 5157 26521 5207 26555
rect 5425 26805 6127 26847
rect 5425 26771 5443 26805
rect 5477 26771 6075 26805
rect 6109 26771 6127 26805
rect 5425 26703 6127 26771
rect 6162 26805 7231 26847
rect 6162 26771 6179 26805
rect 6213 26771 7179 26805
rect 7213 26771 7231 26805
rect 6162 26760 7231 26771
rect 7265 26776 7323 26847
rect 5425 26669 5443 26703
rect 5477 26669 6075 26703
rect 6109 26669 6127 26703
rect 5425 26629 6127 26669
rect 5425 26559 5763 26629
rect 5425 26525 5503 26559
rect 5537 26525 5606 26559
rect 5640 26525 5709 26559
rect 5743 26525 5763 26559
rect 5797 26561 5817 26595
rect 5851 26561 5916 26595
rect 5950 26561 6015 26595
rect 6049 26561 6127 26595
rect 5797 26491 6127 26561
rect 6480 26559 6550 26760
rect 7265 26742 7277 26776
rect 7311 26742 7323 26776
rect 7265 26683 7323 26742
rect 7265 26649 7277 26683
rect 7311 26649 7323 26683
rect 7265 26614 7323 26649
rect 7449 26805 7967 26847
rect 7449 26771 7467 26805
rect 7501 26771 7915 26805
rect 7949 26771 7967 26805
rect 7449 26703 7967 26771
rect 8002 26805 9071 26847
rect 8002 26771 8019 26805
rect 8053 26771 9019 26805
rect 9053 26771 9071 26805
rect 8002 26760 9071 26771
rect 9106 26805 10175 26847
rect 9106 26771 9123 26805
rect 9157 26771 10123 26805
rect 10157 26771 10175 26805
rect 9106 26760 10175 26771
rect 10210 26805 11279 26847
rect 10210 26771 10227 26805
rect 10261 26771 11227 26805
rect 11261 26771 11279 26805
rect 10210 26760 11279 26771
rect 11314 26805 12383 26847
rect 11314 26771 11331 26805
rect 11365 26771 12331 26805
rect 12365 26771 12383 26805
rect 11314 26760 12383 26771
rect 12417 26776 12475 26847
rect 7449 26669 7467 26703
rect 7501 26669 7915 26703
rect 7949 26669 7967 26703
rect 7449 26629 7967 26669
rect 6480 26525 6499 26559
rect 6533 26525 6550 26559
rect 6480 26510 6550 26525
rect 6846 26595 6914 26612
rect 6846 26561 6863 26595
rect 6897 26561 6914 26595
rect 4965 26434 5207 26487
rect 4965 26400 4983 26434
rect 5017 26400 5155 26434
rect 5189 26400 5207 26434
rect 4965 26337 5207 26400
rect 5425 26432 6127 26491
rect 6846 26446 6914 26561
rect 7449 26559 7691 26629
rect 7449 26525 7527 26559
rect 7561 26525 7637 26559
rect 7671 26525 7691 26559
rect 7725 26561 7745 26595
rect 7779 26561 7855 26595
rect 7889 26561 7967 26595
rect 7725 26491 7967 26561
rect 8320 26559 8390 26760
rect 8320 26525 8339 26559
rect 8373 26525 8390 26559
rect 8320 26510 8390 26525
rect 8686 26595 8754 26612
rect 8686 26561 8703 26595
rect 8737 26561 8754 26595
rect 7265 26465 7323 26482
rect 5425 26398 5443 26432
rect 5477 26398 6075 26432
rect 6109 26398 6127 26432
rect 5425 26337 6127 26398
rect 6162 26432 7231 26446
rect 6162 26398 6179 26432
rect 6213 26398 7179 26432
rect 7213 26398 7231 26432
rect 6162 26337 7231 26398
rect 7265 26431 7277 26465
rect 7311 26431 7323 26465
rect 7265 26337 7323 26431
rect 7449 26432 7967 26491
rect 8686 26446 8754 26561
rect 9424 26559 9494 26760
rect 9424 26525 9443 26559
rect 9477 26525 9494 26559
rect 9424 26510 9494 26525
rect 9790 26595 9858 26612
rect 9790 26561 9807 26595
rect 9841 26561 9858 26595
rect 9790 26446 9858 26561
rect 10528 26559 10598 26760
rect 10528 26525 10547 26559
rect 10581 26525 10598 26559
rect 10528 26510 10598 26525
rect 10894 26595 10962 26612
rect 10894 26561 10911 26595
rect 10945 26561 10962 26595
rect 10894 26446 10962 26561
rect 11632 26559 11702 26760
rect 12417 26742 12429 26776
rect 12463 26742 12475 26776
rect 12417 26683 12475 26742
rect 12417 26649 12429 26683
rect 12463 26649 12475 26683
rect 12417 26614 12475 26649
rect 12601 26805 13119 26847
rect 12601 26771 12619 26805
rect 12653 26771 13067 26805
rect 13101 26771 13119 26805
rect 12601 26703 13119 26771
rect 13154 26805 14223 26847
rect 13154 26771 13171 26805
rect 13205 26771 14171 26805
rect 14205 26771 14223 26805
rect 13154 26760 14223 26771
rect 14258 26805 15327 26847
rect 14258 26771 14275 26805
rect 14309 26771 15275 26805
rect 15309 26771 15327 26805
rect 14258 26760 15327 26771
rect 15362 26805 16431 26847
rect 15362 26771 15379 26805
rect 15413 26771 16379 26805
rect 16413 26771 16431 26805
rect 15362 26760 16431 26771
rect 16466 26805 17535 26847
rect 16466 26771 16483 26805
rect 16517 26771 17483 26805
rect 17517 26771 17535 26805
rect 16466 26760 17535 26771
rect 17569 26776 17627 26847
rect 12601 26669 12619 26703
rect 12653 26669 13067 26703
rect 13101 26669 13119 26703
rect 12601 26629 13119 26669
rect 11632 26525 11651 26559
rect 11685 26525 11702 26559
rect 11632 26510 11702 26525
rect 11998 26595 12066 26612
rect 11998 26561 12015 26595
rect 12049 26561 12066 26595
rect 11998 26446 12066 26561
rect 12601 26559 12843 26629
rect 12601 26525 12679 26559
rect 12713 26525 12789 26559
rect 12823 26525 12843 26559
rect 12877 26561 12897 26595
rect 12931 26561 13007 26595
rect 13041 26561 13119 26595
rect 12877 26491 13119 26561
rect 13472 26559 13542 26760
rect 13472 26525 13491 26559
rect 13525 26525 13542 26559
rect 13472 26510 13542 26525
rect 13838 26595 13906 26612
rect 13838 26561 13855 26595
rect 13889 26561 13906 26595
rect 12417 26465 12475 26482
rect 7449 26398 7467 26432
rect 7501 26398 7915 26432
rect 7949 26398 7967 26432
rect 7449 26337 7967 26398
rect 8002 26432 9071 26446
rect 8002 26398 8019 26432
rect 8053 26398 9019 26432
rect 9053 26398 9071 26432
rect 8002 26337 9071 26398
rect 9106 26432 10175 26446
rect 9106 26398 9123 26432
rect 9157 26398 10123 26432
rect 10157 26398 10175 26432
rect 9106 26337 10175 26398
rect 10210 26432 11279 26446
rect 10210 26398 10227 26432
rect 10261 26398 11227 26432
rect 11261 26398 11279 26432
rect 10210 26337 11279 26398
rect 11314 26432 12383 26446
rect 11314 26398 11331 26432
rect 11365 26398 12331 26432
rect 12365 26398 12383 26432
rect 11314 26337 12383 26398
rect 12417 26431 12429 26465
rect 12463 26431 12475 26465
rect 12417 26337 12475 26431
rect 12601 26432 13119 26491
rect 13838 26446 13906 26561
rect 14576 26559 14646 26760
rect 14576 26525 14595 26559
rect 14629 26525 14646 26559
rect 14576 26510 14646 26525
rect 14942 26595 15010 26612
rect 14942 26561 14959 26595
rect 14993 26561 15010 26595
rect 14942 26446 15010 26561
rect 15680 26559 15750 26760
rect 15680 26525 15699 26559
rect 15733 26525 15750 26559
rect 15680 26510 15750 26525
rect 16046 26595 16114 26612
rect 16046 26561 16063 26595
rect 16097 26561 16114 26595
rect 16046 26446 16114 26561
rect 16784 26559 16854 26760
rect 17569 26742 17581 26776
rect 17615 26742 17627 26776
rect 17754 26805 18823 26847
rect 17754 26771 17771 26805
rect 17805 26771 18771 26805
rect 18805 26771 18823 26805
rect 17754 26760 18823 26771
rect 18858 26805 19927 26847
rect 18858 26771 18875 26805
rect 18909 26771 19875 26805
rect 19909 26771 19927 26805
rect 18858 26760 19927 26771
rect 19961 26805 20203 26847
rect 19961 26771 19979 26805
rect 20013 26771 20151 26805
rect 20185 26771 20203 26805
rect 17569 26683 17627 26742
rect 17569 26649 17581 26683
rect 17615 26649 17627 26683
rect 17569 26614 17627 26649
rect 16784 26525 16803 26559
rect 16837 26525 16854 26559
rect 16784 26510 16854 26525
rect 17150 26595 17218 26612
rect 17150 26561 17167 26595
rect 17201 26561 17218 26595
rect 17150 26446 17218 26561
rect 18072 26559 18142 26760
rect 18072 26525 18091 26559
rect 18125 26525 18142 26559
rect 18072 26510 18142 26525
rect 18438 26595 18506 26612
rect 18438 26561 18455 26595
rect 18489 26561 18506 26595
rect 17569 26465 17627 26482
rect 12601 26398 12619 26432
rect 12653 26398 13067 26432
rect 13101 26398 13119 26432
rect 12601 26337 13119 26398
rect 13154 26432 14223 26446
rect 13154 26398 13171 26432
rect 13205 26398 14171 26432
rect 14205 26398 14223 26432
rect 13154 26337 14223 26398
rect 14258 26432 15327 26446
rect 14258 26398 14275 26432
rect 14309 26398 15275 26432
rect 15309 26398 15327 26432
rect 14258 26337 15327 26398
rect 15362 26432 16431 26446
rect 15362 26398 15379 26432
rect 15413 26398 16379 26432
rect 16413 26398 16431 26432
rect 15362 26337 16431 26398
rect 16466 26432 17535 26446
rect 16466 26398 16483 26432
rect 16517 26398 17483 26432
rect 17517 26398 17535 26432
rect 16466 26337 17535 26398
rect 17569 26431 17581 26465
rect 17615 26431 17627 26465
rect 18438 26446 18506 26561
rect 19176 26559 19246 26760
rect 19961 26710 20203 26771
rect 19961 26676 19979 26710
rect 20013 26676 20151 26710
rect 20185 26676 20203 26710
rect 19961 26629 20203 26676
rect 19176 26525 19195 26559
rect 19229 26525 19246 26559
rect 19176 26510 19246 26525
rect 19542 26595 19610 26612
rect 19542 26561 19559 26595
rect 19593 26561 19610 26595
rect 19542 26446 19610 26561
rect 19961 26555 20065 26629
rect 19961 26521 20011 26555
rect 20045 26521 20065 26555
rect 20099 26561 20119 26595
rect 20153 26561 20203 26595
rect 20099 26487 20203 26561
rect 17569 26337 17627 26431
rect 17754 26432 18823 26446
rect 17754 26398 17771 26432
rect 17805 26398 18771 26432
rect 18805 26398 18823 26432
rect 17754 26337 18823 26398
rect 18858 26432 19927 26446
rect 18858 26398 18875 26432
rect 18909 26398 19875 26432
rect 19909 26398 19927 26432
rect 18858 26337 19927 26398
rect 19961 26434 20203 26487
rect 19961 26400 19979 26434
rect 20013 26400 20151 26434
rect 20185 26400 20203 26434
rect 19961 26337 20203 26400
rect 4948 26303 4977 26337
rect 5011 26303 5069 26337
rect 5103 26303 5161 26337
rect 5195 26303 5253 26337
rect 5287 26303 5345 26337
rect 5379 26303 5437 26337
rect 5471 26303 5529 26337
rect 5563 26303 5621 26337
rect 5655 26303 5713 26337
rect 5747 26303 5805 26337
rect 5839 26303 5897 26337
rect 5931 26303 5989 26337
rect 6023 26303 6081 26337
rect 6115 26303 6173 26337
rect 6207 26303 6265 26337
rect 6299 26303 6357 26337
rect 6391 26303 6449 26337
rect 6483 26303 6541 26337
rect 6575 26303 6633 26337
rect 6667 26303 6725 26337
rect 6759 26303 6817 26337
rect 6851 26303 6909 26337
rect 6943 26303 7001 26337
rect 7035 26303 7093 26337
rect 7127 26303 7185 26337
rect 7219 26303 7277 26337
rect 7311 26303 7369 26337
rect 7403 26303 7461 26337
rect 7495 26303 7553 26337
rect 7587 26303 7645 26337
rect 7679 26303 7737 26337
rect 7771 26303 7829 26337
rect 7863 26303 7921 26337
rect 7955 26303 8013 26337
rect 8047 26303 8105 26337
rect 8139 26303 8197 26337
rect 8231 26303 8289 26337
rect 8323 26303 8381 26337
rect 8415 26303 8473 26337
rect 8507 26303 8565 26337
rect 8599 26303 8657 26337
rect 8691 26303 8749 26337
rect 8783 26303 8841 26337
rect 8875 26303 8933 26337
rect 8967 26303 9025 26337
rect 9059 26303 9117 26337
rect 9151 26303 9209 26337
rect 9243 26303 9301 26337
rect 9335 26303 9393 26337
rect 9427 26303 9485 26337
rect 9519 26303 9577 26337
rect 9611 26303 9669 26337
rect 9703 26303 9761 26337
rect 9795 26303 9853 26337
rect 9887 26303 9945 26337
rect 9979 26303 10037 26337
rect 10071 26303 10129 26337
rect 10163 26303 10221 26337
rect 10255 26303 10313 26337
rect 10347 26303 10405 26337
rect 10439 26303 10497 26337
rect 10531 26303 10589 26337
rect 10623 26303 10681 26337
rect 10715 26303 10773 26337
rect 10807 26303 10865 26337
rect 10899 26303 10957 26337
rect 10991 26303 11049 26337
rect 11083 26303 11141 26337
rect 11175 26303 11233 26337
rect 11267 26303 11325 26337
rect 11359 26303 11417 26337
rect 11451 26303 11509 26337
rect 11543 26303 11601 26337
rect 11635 26303 11693 26337
rect 11727 26303 11785 26337
rect 11819 26303 11877 26337
rect 11911 26303 11969 26337
rect 12003 26303 12061 26337
rect 12095 26303 12153 26337
rect 12187 26303 12245 26337
rect 12279 26303 12337 26337
rect 12371 26303 12429 26337
rect 12463 26303 12521 26337
rect 12555 26303 12613 26337
rect 12647 26303 12705 26337
rect 12739 26303 12797 26337
rect 12831 26303 12889 26337
rect 12923 26303 12981 26337
rect 13015 26303 13073 26337
rect 13107 26303 13165 26337
rect 13199 26303 13257 26337
rect 13291 26303 13349 26337
rect 13383 26303 13441 26337
rect 13475 26303 13533 26337
rect 13567 26303 13625 26337
rect 13659 26303 13717 26337
rect 13751 26303 13809 26337
rect 13843 26303 13901 26337
rect 13935 26303 13993 26337
rect 14027 26303 14085 26337
rect 14119 26303 14177 26337
rect 14211 26303 14269 26337
rect 14303 26303 14361 26337
rect 14395 26303 14453 26337
rect 14487 26303 14545 26337
rect 14579 26303 14637 26337
rect 14671 26303 14729 26337
rect 14763 26303 14821 26337
rect 14855 26303 14913 26337
rect 14947 26303 15005 26337
rect 15039 26303 15097 26337
rect 15131 26303 15189 26337
rect 15223 26303 15281 26337
rect 15315 26303 15373 26337
rect 15407 26303 15465 26337
rect 15499 26303 15557 26337
rect 15591 26303 15649 26337
rect 15683 26303 15741 26337
rect 15775 26303 15833 26337
rect 15867 26303 15925 26337
rect 15959 26303 16017 26337
rect 16051 26303 16109 26337
rect 16143 26303 16201 26337
rect 16235 26303 16293 26337
rect 16327 26303 16385 26337
rect 16419 26303 16477 26337
rect 16511 26303 16569 26337
rect 16603 26303 16661 26337
rect 16695 26303 16753 26337
rect 16787 26303 16845 26337
rect 16879 26303 16937 26337
rect 16971 26303 17029 26337
rect 17063 26303 17121 26337
rect 17155 26303 17213 26337
rect 17247 26303 17305 26337
rect 17339 26303 17397 26337
rect 17431 26303 17489 26337
rect 17523 26303 17581 26337
rect 17615 26303 17673 26337
rect 17707 26303 17765 26337
rect 17799 26303 17857 26337
rect 17891 26303 17949 26337
rect 17983 26303 18041 26337
rect 18075 26303 18133 26337
rect 18167 26303 18225 26337
rect 18259 26303 18317 26337
rect 18351 26303 18409 26337
rect 18443 26303 18501 26337
rect 18535 26303 18593 26337
rect 18627 26303 18685 26337
rect 18719 26303 18777 26337
rect 18811 26303 18869 26337
rect 18903 26303 18961 26337
rect 18995 26303 19053 26337
rect 19087 26303 19145 26337
rect 19179 26303 19237 26337
rect 19271 26303 19329 26337
rect 19363 26303 19421 26337
rect 19455 26303 19513 26337
rect 19547 26303 19605 26337
rect 19639 26303 19697 26337
rect 19731 26303 19789 26337
rect 19823 26303 19881 26337
rect 19915 26303 19973 26337
rect 20007 26303 20065 26337
rect 20099 26303 20157 26337
rect 20191 26303 20220 26337
rect 4965 26240 5207 26303
rect 4965 26206 4983 26240
rect 5017 26206 5155 26240
rect 5189 26206 5207 26240
rect 4965 26153 5207 26206
rect 5426 26242 6495 26303
rect 5426 26208 5443 26242
rect 5477 26208 6443 26242
rect 6477 26208 6495 26242
rect 5426 26194 6495 26208
rect 6530 26242 7599 26303
rect 6530 26208 6547 26242
rect 6581 26208 7547 26242
rect 7581 26208 7599 26242
rect 6530 26194 7599 26208
rect 7634 26242 8703 26303
rect 7634 26208 7651 26242
rect 7685 26208 8651 26242
rect 8685 26208 8703 26242
rect 7634 26194 8703 26208
rect 8738 26242 9807 26303
rect 8738 26208 8755 26242
rect 8789 26208 9755 26242
rect 9789 26208 9807 26242
rect 8738 26194 9807 26208
rect 9841 26209 9899 26303
rect 4965 26079 5069 26153
rect 4965 26045 5015 26079
rect 5049 26045 5069 26079
rect 5103 26085 5123 26119
rect 5157 26085 5207 26119
rect 5103 26011 5207 26085
rect 4965 25964 5207 26011
rect 4965 25930 4983 25964
rect 5017 25930 5155 25964
rect 5189 25930 5207 25964
rect 4965 25869 5207 25930
rect 5744 26115 5814 26130
rect 5744 26081 5763 26115
rect 5797 26081 5814 26115
rect 5744 25880 5814 26081
rect 6110 26079 6178 26194
rect 6110 26045 6127 26079
rect 6161 26045 6178 26079
rect 6110 26028 6178 26045
rect 6848 26115 6918 26130
rect 6848 26081 6867 26115
rect 6901 26081 6918 26115
rect 6848 25880 6918 26081
rect 7214 26079 7282 26194
rect 7214 26045 7231 26079
rect 7265 26045 7282 26079
rect 7214 26028 7282 26045
rect 7952 26115 8022 26130
rect 7952 26081 7971 26115
rect 8005 26081 8022 26115
rect 7952 25880 8022 26081
rect 8318 26079 8386 26194
rect 8318 26045 8335 26079
rect 8369 26045 8386 26079
rect 8318 26028 8386 26045
rect 9056 26115 9126 26130
rect 9056 26081 9075 26115
rect 9109 26081 9126 26115
rect 9056 25880 9126 26081
rect 9422 26079 9490 26194
rect 9841 26175 9853 26209
rect 9887 26175 9899 26209
rect 9841 26158 9899 26175
rect 10025 26242 10543 26303
rect 10025 26208 10043 26242
rect 10077 26208 10491 26242
rect 10525 26208 10543 26242
rect 10025 26149 10543 26208
rect 10578 26242 11647 26303
rect 10578 26208 10595 26242
rect 10629 26208 11595 26242
rect 11629 26208 11647 26242
rect 10578 26194 11647 26208
rect 11682 26242 12751 26303
rect 11682 26208 11699 26242
rect 11733 26208 12699 26242
rect 12733 26208 12751 26242
rect 11682 26194 12751 26208
rect 12786 26242 13855 26303
rect 12786 26208 12803 26242
rect 12837 26208 13803 26242
rect 13837 26208 13855 26242
rect 12786 26194 13855 26208
rect 13890 26242 14959 26303
rect 13890 26208 13907 26242
rect 13941 26208 14907 26242
rect 14941 26208 14959 26242
rect 13890 26194 14959 26208
rect 14993 26209 15051 26303
rect 9422 26045 9439 26079
rect 9473 26045 9490 26079
rect 9422 26028 9490 26045
rect 10025 26081 10103 26115
rect 10137 26081 10213 26115
rect 10247 26081 10267 26115
rect 9841 25991 9899 26026
rect 9841 25957 9853 25991
rect 9887 25957 9899 25991
rect 9841 25898 9899 25957
rect 4965 25835 4983 25869
rect 5017 25835 5155 25869
rect 5189 25835 5207 25869
rect 4965 25793 5207 25835
rect 5426 25869 6495 25880
rect 5426 25835 5443 25869
rect 5477 25835 6443 25869
rect 6477 25835 6495 25869
rect 5426 25793 6495 25835
rect 6530 25869 7599 25880
rect 6530 25835 6547 25869
rect 6581 25835 7547 25869
rect 7581 25835 7599 25869
rect 6530 25793 7599 25835
rect 7634 25869 8703 25880
rect 7634 25835 7651 25869
rect 7685 25835 8651 25869
rect 8685 25835 8703 25869
rect 7634 25793 8703 25835
rect 8738 25869 9807 25880
rect 8738 25835 8755 25869
rect 8789 25835 9755 25869
rect 9789 25835 9807 25869
rect 8738 25793 9807 25835
rect 9841 25864 9853 25898
rect 9887 25864 9899 25898
rect 9841 25793 9899 25864
rect 10025 26011 10267 26081
rect 10301 26079 10543 26149
rect 10301 26045 10321 26079
rect 10355 26045 10431 26079
rect 10465 26045 10543 26079
rect 10896 26115 10966 26130
rect 10896 26081 10915 26115
rect 10949 26081 10966 26115
rect 10025 25971 10543 26011
rect 10025 25937 10043 25971
rect 10077 25937 10491 25971
rect 10525 25937 10543 25971
rect 10025 25869 10543 25937
rect 10896 25880 10966 26081
rect 11262 26079 11330 26194
rect 11262 26045 11279 26079
rect 11313 26045 11330 26079
rect 11262 26028 11330 26045
rect 12000 26115 12070 26130
rect 12000 26081 12019 26115
rect 12053 26081 12070 26115
rect 12000 25880 12070 26081
rect 12366 26079 12434 26194
rect 12366 26045 12383 26079
rect 12417 26045 12434 26079
rect 12366 26028 12434 26045
rect 13104 26115 13174 26130
rect 13104 26081 13123 26115
rect 13157 26081 13174 26115
rect 13104 25880 13174 26081
rect 13470 26079 13538 26194
rect 13470 26045 13487 26079
rect 13521 26045 13538 26079
rect 13470 26028 13538 26045
rect 14208 26115 14278 26130
rect 14208 26081 14227 26115
rect 14261 26081 14278 26115
rect 14208 25880 14278 26081
rect 14574 26079 14642 26194
rect 14993 26175 15005 26209
rect 15039 26175 15051 26209
rect 14993 26158 15051 26175
rect 15177 26235 15511 26303
rect 15177 26201 15195 26235
rect 15229 26201 15459 26235
rect 15493 26201 15511 26235
rect 15177 26149 15511 26201
rect 15546 26242 16615 26303
rect 15546 26208 15563 26242
rect 15597 26208 16563 26242
rect 16597 26208 16615 26242
rect 15546 26194 16615 26208
rect 16650 26242 17719 26303
rect 16650 26208 16667 26242
rect 16701 26208 17667 26242
rect 17701 26208 17719 26242
rect 16650 26194 17719 26208
rect 17754 26242 18823 26303
rect 17754 26208 17771 26242
rect 17805 26208 18771 26242
rect 18805 26208 18823 26242
rect 17754 26194 18823 26208
rect 18858 26242 19927 26303
rect 18858 26208 18875 26242
rect 18909 26208 19875 26242
rect 19909 26208 19927 26242
rect 18858 26194 19927 26208
rect 19961 26240 20203 26303
rect 19961 26206 19979 26240
rect 20013 26206 20151 26240
rect 20185 26206 20203 26240
rect 14574 26045 14591 26079
rect 14625 26045 14642 26079
rect 14574 26028 14642 26045
rect 15177 26081 15197 26115
rect 15231 26081 15327 26115
rect 14993 25991 15051 26026
rect 14993 25957 15005 25991
rect 15039 25957 15051 25991
rect 14993 25898 15051 25957
rect 10025 25835 10043 25869
rect 10077 25835 10491 25869
rect 10525 25835 10543 25869
rect 10025 25793 10543 25835
rect 10578 25869 11647 25880
rect 10578 25835 10595 25869
rect 10629 25835 11595 25869
rect 11629 25835 11647 25869
rect 10578 25793 11647 25835
rect 11682 25869 12751 25880
rect 11682 25835 11699 25869
rect 11733 25835 12699 25869
rect 12733 25835 12751 25869
rect 11682 25793 12751 25835
rect 12786 25869 13855 25880
rect 12786 25835 12803 25869
rect 12837 25835 13803 25869
rect 13837 25835 13855 25869
rect 12786 25793 13855 25835
rect 13890 25869 14959 25880
rect 13890 25835 13907 25869
rect 13941 25835 14907 25869
rect 14941 25835 14959 25869
rect 13890 25793 14959 25835
rect 14993 25864 15005 25898
rect 15039 25864 15051 25898
rect 14993 25793 15051 25864
rect 15177 26011 15327 26081
rect 15361 26079 15511 26149
rect 15361 26045 15457 26079
rect 15491 26045 15511 26079
rect 15864 26115 15934 26130
rect 15864 26081 15883 26115
rect 15917 26081 15934 26115
rect 15177 25971 15511 26011
rect 15177 25937 15195 25971
rect 15229 25937 15459 25971
rect 15493 25937 15511 25971
rect 15177 25869 15511 25937
rect 15864 25880 15934 26081
rect 16230 26079 16298 26194
rect 16230 26045 16247 26079
rect 16281 26045 16298 26079
rect 16230 26028 16298 26045
rect 16968 26115 17038 26130
rect 16968 26081 16987 26115
rect 17021 26081 17038 26115
rect 16968 25880 17038 26081
rect 17334 26079 17402 26194
rect 17334 26045 17351 26079
rect 17385 26045 17402 26079
rect 17334 26028 17402 26045
rect 18072 26115 18142 26130
rect 18072 26081 18091 26115
rect 18125 26081 18142 26115
rect 18072 25880 18142 26081
rect 18438 26079 18506 26194
rect 18438 26045 18455 26079
rect 18489 26045 18506 26079
rect 18438 26028 18506 26045
rect 19176 26115 19246 26130
rect 19176 26081 19195 26115
rect 19229 26081 19246 26115
rect 19176 25880 19246 26081
rect 19542 26079 19610 26194
rect 19961 26153 20203 26206
rect 19542 26045 19559 26079
rect 19593 26045 19610 26079
rect 19542 26028 19610 26045
rect 19961 26085 20011 26119
rect 20045 26085 20065 26119
rect 19961 26011 20065 26085
rect 20099 26079 20203 26153
rect 20099 26045 20119 26079
rect 20153 26045 20203 26079
rect 19961 25964 20203 26011
rect 19961 25930 19979 25964
rect 20013 25930 20151 25964
rect 20185 25930 20203 25964
rect 15177 25835 15195 25869
rect 15229 25835 15459 25869
rect 15493 25835 15511 25869
rect 15177 25793 15511 25835
rect 15546 25869 16615 25880
rect 15546 25835 15563 25869
rect 15597 25835 16563 25869
rect 16597 25835 16615 25869
rect 15546 25793 16615 25835
rect 16650 25869 17719 25880
rect 16650 25835 16667 25869
rect 16701 25835 17667 25869
rect 17701 25835 17719 25869
rect 16650 25793 17719 25835
rect 17754 25869 18823 25880
rect 17754 25835 17771 25869
rect 17805 25835 18771 25869
rect 18805 25835 18823 25869
rect 17754 25793 18823 25835
rect 18858 25869 19927 25880
rect 18858 25835 18875 25869
rect 18909 25835 19875 25869
rect 19909 25835 19927 25869
rect 18858 25793 19927 25835
rect 19961 25869 20203 25930
rect 19961 25835 19979 25869
rect 20013 25835 20151 25869
rect 20185 25835 20203 25869
rect 19961 25793 20203 25835
rect 4948 25759 4977 25793
rect 5011 25759 5069 25793
rect 5103 25759 5161 25793
rect 5195 25759 5253 25793
rect 5287 25759 5345 25793
rect 5379 25759 5437 25793
rect 5471 25759 5529 25793
rect 5563 25759 5621 25793
rect 5655 25759 5713 25793
rect 5747 25759 5805 25793
rect 5839 25759 5897 25793
rect 5931 25759 5989 25793
rect 6023 25759 6081 25793
rect 6115 25759 6173 25793
rect 6207 25759 6265 25793
rect 6299 25759 6357 25793
rect 6391 25759 6449 25793
rect 6483 25759 6541 25793
rect 6575 25759 6633 25793
rect 6667 25759 6725 25793
rect 6759 25759 6817 25793
rect 6851 25759 6909 25793
rect 6943 25759 7001 25793
rect 7035 25759 7093 25793
rect 7127 25759 7185 25793
rect 7219 25759 7277 25793
rect 7311 25759 7369 25793
rect 7403 25759 7461 25793
rect 7495 25759 7553 25793
rect 7587 25759 7645 25793
rect 7679 25759 7737 25793
rect 7771 25759 7829 25793
rect 7863 25759 7921 25793
rect 7955 25759 8013 25793
rect 8047 25759 8105 25793
rect 8139 25759 8197 25793
rect 8231 25759 8289 25793
rect 8323 25759 8381 25793
rect 8415 25759 8473 25793
rect 8507 25759 8565 25793
rect 8599 25759 8657 25793
rect 8691 25759 8749 25793
rect 8783 25759 8841 25793
rect 8875 25759 8933 25793
rect 8967 25759 9025 25793
rect 9059 25759 9117 25793
rect 9151 25759 9209 25793
rect 9243 25759 9301 25793
rect 9335 25759 9393 25793
rect 9427 25759 9485 25793
rect 9519 25759 9577 25793
rect 9611 25759 9669 25793
rect 9703 25759 9761 25793
rect 9795 25759 9853 25793
rect 9887 25759 9945 25793
rect 9979 25759 10037 25793
rect 10071 25759 10129 25793
rect 10163 25759 10221 25793
rect 10255 25759 10313 25793
rect 10347 25759 10405 25793
rect 10439 25759 10497 25793
rect 10531 25759 10589 25793
rect 10623 25759 10681 25793
rect 10715 25759 10773 25793
rect 10807 25759 10865 25793
rect 10899 25759 10957 25793
rect 10991 25759 11049 25793
rect 11083 25759 11141 25793
rect 11175 25759 11233 25793
rect 11267 25759 11325 25793
rect 11359 25759 11417 25793
rect 11451 25759 11509 25793
rect 11543 25759 11601 25793
rect 11635 25759 11693 25793
rect 11727 25759 11785 25793
rect 11819 25759 11877 25793
rect 11911 25759 11969 25793
rect 12003 25759 12061 25793
rect 12095 25759 12153 25793
rect 12187 25759 12245 25793
rect 12279 25759 12337 25793
rect 12371 25759 12429 25793
rect 12463 25759 12521 25793
rect 12555 25759 12613 25793
rect 12647 25759 12705 25793
rect 12739 25759 12797 25793
rect 12831 25759 12889 25793
rect 12923 25759 12981 25793
rect 13015 25759 13073 25793
rect 13107 25759 13165 25793
rect 13199 25759 13257 25793
rect 13291 25759 13349 25793
rect 13383 25759 13441 25793
rect 13475 25759 13533 25793
rect 13567 25759 13625 25793
rect 13659 25759 13717 25793
rect 13751 25759 13809 25793
rect 13843 25759 13901 25793
rect 13935 25759 13993 25793
rect 14027 25759 14085 25793
rect 14119 25759 14177 25793
rect 14211 25759 14269 25793
rect 14303 25759 14361 25793
rect 14395 25759 14453 25793
rect 14487 25759 14545 25793
rect 14579 25759 14637 25793
rect 14671 25759 14729 25793
rect 14763 25759 14821 25793
rect 14855 25759 14913 25793
rect 14947 25759 15005 25793
rect 15039 25759 15097 25793
rect 15131 25759 15189 25793
rect 15223 25759 15281 25793
rect 15315 25759 15373 25793
rect 15407 25759 15465 25793
rect 15499 25759 15557 25793
rect 15591 25759 15649 25793
rect 15683 25759 15741 25793
rect 15775 25759 15833 25793
rect 15867 25759 15925 25793
rect 15959 25759 16017 25793
rect 16051 25759 16109 25793
rect 16143 25759 16201 25793
rect 16235 25759 16293 25793
rect 16327 25759 16385 25793
rect 16419 25759 16477 25793
rect 16511 25759 16569 25793
rect 16603 25759 16661 25793
rect 16695 25759 16753 25793
rect 16787 25759 16845 25793
rect 16879 25759 16937 25793
rect 16971 25759 17029 25793
rect 17063 25759 17121 25793
rect 17155 25759 17213 25793
rect 17247 25759 17305 25793
rect 17339 25759 17397 25793
rect 17431 25759 17489 25793
rect 17523 25759 17581 25793
rect 17615 25759 17673 25793
rect 17707 25759 17765 25793
rect 17799 25759 17857 25793
rect 17891 25759 17949 25793
rect 17983 25759 18041 25793
rect 18075 25759 18133 25793
rect 18167 25759 18225 25793
rect 18259 25759 18317 25793
rect 18351 25759 18409 25793
rect 18443 25759 18501 25793
rect 18535 25759 18593 25793
rect 18627 25759 18685 25793
rect 18719 25759 18777 25793
rect 18811 25759 18869 25793
rect 18903 25759 18961 25793
rect 18995 25759 19053 25793
rect 19087 25759 19145 25793
rect 19179 25759 19237 25793
rect 19271 25759 19329 25793
rect 19363 25759 19421 25793
rect 19455 25759 19513 25793
rect 19547 25759 19605 25793
rect 19639 25759 19697 25793
rect 19731 25759 19789 25793
rect 19823 25759 19881 25793
rect 19915 25759 19973 25793
rect 20007 25759 20065 25793
rect 20099 25759 20157 25793
rect 20191 25759 20220 25793
rect 4965 25717 5207 25759
rect 4965 25683 4983 25717
rect 5017 25683 5155 25717
rect 5189 25683 5207 25717
rect 4965 25622 5207 25683
rect 4965 25588 4983 25622
rect 5017 25588 5155 25622
rect 5189 25588 5207 25622
rect 4965 25541 5207 25588
rect 4965 25473 5015 25507
rect 5049 25473 5069 25507
rect 4965 25399 5069 25473
rect 5103 25467 5207 25541
rect 5103 25433 5123 25467
rect 5157 25433 5207 25467
rect 5425 25717 6127 25759
rect 5425 25683 5443 25717
rect 5477 25683 6075 25717
rect 6109 25683 6127 25717
rect 5425 25615 6127 25683
rect 6162 25717 7231 25759
rect 6162 25683 6179 25717
rect 6213 25683 7179 25717
rect 7213 25683 7231 25717
rect 6162 25672 7231 25683
rect 7265 25688 7323 25759
rect 5425 25581 5443 25615
rect 5477 25581 6075 25615
rect 6109 25581 6127 25615
rect 5425 25541 6127 25581
rect 5425 25471 5763 25541
rect 5425 25437 5503 25471
rect 5537 25437 5606 25471
rect 5640 25437 5709 25471
rect 5743 25437 5763 25471
rect 5797 25473 5817 25507
rect 5851 25473 5916 25507
rect 5950 25473 6015 25507
rect 6049 25473 6127 25507
rect 5797 25403 6127 25473
rect 6480 25471 6550 25672
rect 7265 25654 7277 25688
rect 7311 25654 7323 25688
rect 7265 25595 7323 25654
rect 7265 25561 7277 25595
rect 7311 25561 7323 25595
rect 7265 25526 7323 25561
rect 7449 25717 7967 25759
rect 7449 25683 7467 25717
rect 7501 25683 7915 25717
rect 7949 25683 7967 25717
rect 7449 25615 7967 25683
rect 8002 25717 9071 25759
rect 8002 25683 8019 25717
rect 8053 25683 9019 25717
rect 9053 25683 9071 25717
rect 8002 25672 9071 25683
rect 9106 25717 10175 25759
rect 9106 25683 9123 25717
rect 9157 25683 10123 25717
rect 10157 25683 10175 25717
rect 9106 25672 10175 25683
rect 10210 25717 11279 25759
rect 10210 25683 10227 25717
rect 10261 25683 11227 25717
rect 11261 25683 11279 25717
rect 10210 25672 11279 25683
rect 11314 25717 12383 25759
rect 11314 25683 11331 25717
rect 11365 25683 12331 25717
rect 12365 25683 12383 25717
rect 11314 25672 12383 25683
rect 12417 25688 12475 25759
rect 7449 25581 7467 25615
rect 7501 25581 7915 25615
rect 7949 25581 7967 25615
rect 7449 25541 7967 25581
rect 6480 25437 6499 25471
rect 6533 25437 6550 25471
rect 6480 25422 6550 25437
rect 6846 25507 6914 25524
rect 6846 25473 6863 25507
rect 6897 25473 6914 25507
rect 4965 25346 5207 25399
rect 4965 25312 4983 25346
rect 5017 25312 5155 25346
rect 5189 25312 5207 25346
rect 4965 25249 5207 25312
rect 5425 25344 6127 25403
rect 6846 25358 6914 25473
rect 7449 25471 7691 25541
rect 7449 25437 7527 25471
rect 7561 25437 7637 25471
rect 7671 25437 7691 25471
rect 7725 25473 7745 25507
rect 7779 25473 7855 25507
rect 7889 25473 7967 25507
rect 7725 25403 7967 25473
rect 8320 25471 8390 25672
rect 8320 25437 8339 25471
rect 8373 25437 8390 25471
rect 8320 25422 8390 25437
rect 8686 25507 8754 25524
rect 8686 25473 8703 25507
rect 8737 25473 8754 25507
rect 7265 25377 7323 25394
rect 5425 25310 5443 25344
rect 5477 25310 6075 25344
rect 6109 25310 6127 25344
rect 5425 25249 6127 25310
rect 6162 25344 7231 25358
rect 6162 25310 6179 25344
rect 6213 25310 7179 25344
rect 7213 25310 7231 25344
rect 6162 25249 7231 25310
rect 7265 25343 7277 25377
rect 7311 25343 7323 25377
rect 7265 25249 7323 25343
rect 7449 25344 7967 25403
rect 8686 25358 8754 25473
rect 9424 25471 9494 25672
rect 9424 25437 9443 25471
rect 9477 25437 9494 25471
rect 9424 25422 9494 25437
rect 9790 25507 9858 25524
rect 9790 25473 9807 25507
rect 9841 25473 9858 25507
rect 9790 25358 9858 25473
rect 10528 25471 10598 25672
rect 10528 25437 10547 25471
rect 10581 25437 10598 25471
rect 10528 25422 10598 25437
rect 10894 25507 10962 25524
rect 10894 25473 10911 25507
rect 10945 25473 10962 25507
rect 10894 25358 10962 25473
rect 11632 25471 11702 25672
rect 12417 25654 12429 25688
rect 12463 25654 12475 25688
rect 12417 25595 12475 25654
rect 12417 25561 12429 25595
rect 12463 25561 12475 25595
rect 12417 25526 12475 25561
rect 12601 25717 13119 25759
rect 12601 25683 12619 25717
rect 12653 25683 13067 25717
rect 13101 25683 13119 25717
rect 12601 25615 13119 25683
rect 13154 25717 14223 25759
rect 13154 25683 13171 25717
rect 13205 25683 14171 25717
rect 14205 25683 14223 25717
rect 13154 25672 14223 25683
rect 14258 25717 15327 25759
rect 14258 25683 14275 25717
rect 14309 25683 15275 25717
rect 15309 25683 15327 25717
rect 14258 25672 15327 25683
rect 15362 25717 16431 25759
rect 15362 25683 15379 25717
rect 15413 25683 16379 25717
rect 16413 25683 16431 25717
rect 15362 25672 16431 25683
rect 16466 25717 17535 25759
rect 16466 25683 16483 25717
rect 16517 25683 17483 25717
rect 17517 25683 17535 25717
rect 16466 25672 17535 25683
rect 17569 25688 17627 25759
rect 12601 25581 12619 25615
rect 12653 25581 13067 25615
rect 13101 25581 13119 25615
rect 12601 25541 13119 25581
rect 11632 25437 11651 25471
rect 11685 25437 11702 25471
rect 11632 25422 11702 25437
rect 11998 25507 12066 25524
rect 11998 25473 12015 25507
rect 12049 25473 12066 25507
rect 11998 25358 12066 25473
rect 12601 25471 12843 25541
rect 12601 25437 12679 25471
rect 12713 25437 12789 25471
rect 12823 25437 12843 25471
rect 12877 25473 12897 25507
rect 12931 25473 13007 25507
rect 13041 25473 13119 25507
rect 12877 25403 13119 25473
rect 13472 25471 13542 25672
rect 13472 25437 13491 25471
rect 13525 25437 13542 25471
rect 13472 25422 13542 25437
rect 13838 25507 13906 25524
rect 13838 25473 13855 25507
rect 13889 25473 13906 25507
rect 12417 25377 12475 25394
rect 7449 25310 7467 25344
rect 7501 25310 7915 25344
rect 7949 25310 7967 25344
rect 7449 25249 7967 25310
rect 8002 25344 9071 25358
rect 8002 25310 8019 25344
rect 8053 25310 9019 25344
rect 9053 25310 9071 25344
rect 8002 25249 9071 25310
rect 9106 25344 10175 25358
rect 9106 25310 9123 25344
rect 9157 25310 10123 25344
rect 10157 25310 10175 25344
rect 9106 25249 10175 25310
rect 10210 25344 11279 25358
rect 10210 25310 10227 25344
rect 10261 25310 11227 25344
rect 11261 25310 11279 25344
rect 10210 25249 11279 25310
rect 11314 25344 12383 25358
rect 11314 25310 11331 25344
rect 11365 25310 12331 25344
rect 12365 25310 12383 25344
rect 11314 25249 12383 25310
rect 12417 25343 12429 25377
rect 12463 25343 12475 25377
rect 12417 25249 12475 25343
rect 12601 25344 13119 25403
rect 13838 25358 13906 25473
rect 14576 25471 14646 25672
rect 14576 25437 14595 25471
rect 14629 25437 14646 25471
rect 14576 25422 14646 25437
rect 14942 25507 15010 25524
rect 14942 25473 14959 25507
rect 14993 25473 15010 25507
rect 14942 25358 15010 25473
rect 15680 25471 15750 25672
rect 15680 25437 15699 25471
rect 15733 25437 15750 25471
rect 15680 25422 15750 25437
rect 16046 25507 16114 25524
rect 16046 25473 16063 25507
rect 16097 25473 16114 25507
rect 16046 25358 16114 25473
rect 16784 25471 16854 25672
rect 17569 25654 17581 25688
rect 17615 25654 17627 25688
rect 17754 25717 18823 25759
rect 17754 25683 17771 25717
rect 17805 25683 18771 25717
rect 18805 25683 18823 25717
rect 17754 25672 18823 25683
rect 18858 25717 19927 25759
rect 18858 25683 18875 25717
rect 18909 25683 19875 25717
rect 19909 25683 19927 25717
rect 18858 25672 19927 25683
rect 19961 25717 20203 25759
rect 19961 25683 19979 25717
rect 20013 25683 20151 25717
rect 20185 25683 20203 25717
rect 17569 25595 17627 25654
rect 17569 25561 17581 25595
rect 17615 25561 17627 25595
rect 17569 25526 17627 25561
rect 16784 25437 16803 25471
rect 16837 25437 16854 25471
rect 16784 25422 16854 25437
rect 17150 25507 17218 25524
rect 17150 25473 17167 25507
rect 17201 25473 17218 25507
rect 17150 25358 17218 25473
rect 18072 25471 18142 25672
rect 18072 25437 18091 25471
rect 18125 25437 18142 25471
rect 18072 25422 18142 25437
rect 18438 25507 18506 25524
rect 18438 25473 18455 25507
rect 18489 25473 18506 25507
rect 17569 25377 17627 25394
rect 12601 25310 12619 25344
rect 12653 25310 13067 25344
rect 13101 25310 13119 25344
rect 12601 25249 13119 25310
rect 13154 25344 14223 25358
rect 13154 25310 13171 25344
rect 13205 25310 14171 25344
rect 14205 25310 14223 25344
rect 13154 25249 14223 25310
rect 14258 25344 15327 25358
rect 14258 25310 14275 25344
rect 14309 25310 15275 25344
rect 15309 25310 15327 25344
rect 14258 25249 15327 25310
rect 15362 25344 16431 25358
rect 15362 25310 15379 25344
rect 15413 25310 16379 25344
rect 16413 25310 16431 25344
rect 15362 25249 16431 25310
rect 16466 25344 17535 25358
rect 16466 25310 16483 25344
rect 16517 25310 17483 25344
rect 17517 25310 17535 25344
rect 16466 25249 17535 25310
rect 17569 25343 17581 25377
rect 17615 25343 17627 25377
rect 18438 25358 18506 25473
rect 19176 25471 19246 25672
rect 19961 25622 20203 25683
rect 19961 25588 19979 25622
rect 20013 25588 20151 25622
rect 20185 25588 20203 25622
rect 19961 25541 20203 25588
rect 19176 25437 19195 25471
rect 19229 25437 19246 25471
rect 19176 25422 19246 25437
rect 19542 25507 19610 25524
rect 19542 25473 19559 25507
rect 19593 25473 19610 25507
rect 19542 25358 19610 25473
rect 19961 25467 20065 25541
rect 19961 25433 20011 25467
rect 20045 25433 20065 25467
rect 20099 25473 20119 25507
rect 20153 25473 20203 25507
rect 20099 25399 20203 25473
rect 17569 25249 17627 25343
rect 17754 25344 18823 25358
rect 17754 25310 17771 25344
rect 17805 25310 18771 25344
rect 18805 25310 18823 25344
rect 17754 25249 18823 25310
rect 18858 25344 19927 25358
rect 18858 25310 18875 25344
rect 18909 25310 19875 25344
rect 19909 25310 19927 25344
rect 18858 25249 19927 25310
rect 19961 25346 20203 25399
rect 19961 25312 19979 25346
rect 20013 25312 20151 25346
rect 20185 25312 20203 25346
rect 19961 25249 20203 25312
rect 4948 25215 4977 25249
rect 5011 25215 5069 25249
rect 5103 25215 5161 25249
rect 5195 25215 5253 25249
rect 5287 25215 5345 25249
rect 5379 25215 5437 25249
rect 5471 25215 5529 25249
rect 5563 25215 5621 25249
rect 5655 25215 5713 25249
rect 5747 25215 5805 25249
rect 5839 25215 5897 25249
rect 5931 25215 5989 25249
rect 6023 25215 6081 25249
rect 6115 25215 6173 25249
rect 6207 25215 6265 25249
rect 6299 25215 6357 25249
rect 6391 25215 6449 25249
rect 6483 25215 6541 25249
rect 6575 25215 6633 25249
rect 6667 25215 6725 25249
rect 6759 25215 6817 25249
rect 6851 25215 6909 25249
rect 6943 25215 7001 25249
rect 7035 25215 7093 25249
rect 7127 25215 7185 25249
rect 7219 25215 7277 25249
rect 7311 25215 7369 25249
rect 7403 25215 7461 25249
rect 7495 25215 7553 25249
rect 7587 25215 7645 25249
rect 7679 25215 7737 25249
rect 7771 25215 7829 25249
rect 7863 25215 7921 25249
rect 7955 25215 8013 25249
rect 8047 25215 8105 25249
rect 8139 25215 8197 25249
rect 8231 25215 8289 25249
rect 8323 25215 8381 25249
rect 8415 25215 8473 25249
rect 8507 25215 8565 25249
rect 8599 25215 8657 25249
rect 8691 25215 8749 25249
rect 8783 25215 8841 25249
rect 8875 25215 8933 25249
rect 8967 25215 9025 25249
rect 9059 25215 9117 25249
rect 9151 25215 9209 25249
rect 9243 25215 9301 25249
rect 9335 25215 9393 25249
rect 9427 25215 9485 25249
rect 9519 25215 9577 25249
rect 9611 25215 9669 25249
rect 9703 25215 9761 25249
rect 9795 25215 9853 25249
rect 9887 25215 9945 25249
rect 9979 25215 10037 25249
rect 10071 25215 10129 25249
rect 10163 25215 10221 25249
rect 10255 25215 10313 25249
rect 10347 25215 10405 25249
rect 10439 25215 10497 25249
rect 10531 25215 10589 25249
rect 10623 25215 10681 25249
rect 10715 25215 10773 25249
rect 10807 25215 10865 25249
rect 10899 25215 10957 25249
rect 10991 25215 11049 25249
rect 11083 25215 11141 25249
rect 11175 25215 11233 25249
rect 11267 25215 11325 25249
rect 11359 25215 11417 25249
rect 11451 25215 11509 25249
rect 11543 25215 11601 25249
rect 11635 25215 11693 25249
rect 11727 25215 11785 25249
rect 11819 25215 11877 25249
rect 11911 25215 11969 25249
rect 12003 25215 12061 25249
rect 12095 25215 12153 25249
rect 12187 25215 12245 25249
rect 12279 25215 12337 25249
rect 12371 25215 12429 25249
rect 12463 25215 12521 25249
rect 12555 25215 12613 25249
rect 12647 25215 12705 25249
rect 12739 25215 12797 25249
rect 12831 25215 12889 25249
rect 12923 25215 12981 25249
rect 13015 25215 13073 25249
rect 13107 25215 13165 25249
rect 13199 25215 13257 25249
rect 13291 25215 13349 25249
rect 13383 25215 13441 25249
rect 13475 25215 13533 25249
rect 13567 25215 13625 25249
rect 13659 25215 13717 25249
rect 13751 25215 13809 25249
rect 13843 25215 13901 25249
rect 13935 25215 13993 25249
rect 14027 25215 14085 25249
rect 14119 25215 14177 25249
rect 14211 25215 14269 25249
rect 14303 25215 14361 25249
rect 14395 25215 14453 25249
rect 14487 25215 14545 25249
rect 14579 25215 14637 25249
rect 14671 25215 14729 25249
rect 14763 25215 14821 25249
rect 14855 25215 14913 25249
rect 14947 25215 15005 25249
rect 15039 25215 15097 25249
rect 15131 25215 15189 25249
rect 15223 25215 15281 25249
rect 15315 25215 15373 25249
rect 15407 25215 15465 25249
rect 15499 25215 15557 25249
rect 15591 25215 15649 25249
rect 15683 25215 15741 25249
rect 15775 25215 15833 25249
rect 15867 25215 15925 25249
rect 15959 25215 16017 25249
rect 16051 25215 16109 25249
rect 16143 25215 16201 25249
rect 16235 25215 16293 25249
rect 16327 25215 16385 25249
rect 16419 25215 16477 25249
rect 16511 25215 16569 25249
rect 16603 25215 16661 25249
rect 16695 25215 16753 25249
rect 16787 25215 16845 25249
rect 16879 25215 16937 25249
rect 16971 25215 17029 25249
rect 17063 25215 17121 25249
rect 17155 25215 17213 25249
rect 17247 25215 17305 25249
rect 17339 25215 17397 25249
rect 17431 25215 17489 25249
rect 17523 25215 17581 25249
rect 17615 25215 17673 25249
rect 17707 25215 17765 25249
rect 17799 25215 17857 25249
rect 17891 25215 17949 25249
rect 17983 25215 18041 25249
rect 18075 25215 18133 25249
rect 18167 25215 18225 25249
rect 18259 25215 18317 25249
rect 18351 25215 18409 25249
rect 18443 25215 18501 25249
rect 18535 25215 18593 25249
rect 18627 25215 18685 25249
rect 18719 25215 18777 25249
rect 18811 25215 18869 25249
rect 18903 25215 18961 25249
rect 18995 25215 19053 25249
rect 19087 25215 19145 25249
rect 19179 25215 19237 25249
rect 19271 25215 19329 25249
rect 19363 25215 19421 25249
rect 19455 25215 19513 25249
rect 19547 25215 19605 25249
rect 19639 25215 19697 25249
rect 19731 25215 19789 25249
rect 19823 25215 19881 25249
rect 19915 25215 19973 25249
rect 20007 25215 20065 25249
rect 20099 25215 20157 25249
rect 20191 25215 20220 25249
rect 4965 25152 5207 25215
rect 4965 25118 4983 25152
rect 5017 25118 5155 25152
rect 5189 25118 5207 25152
rect 4965 25065 5207 25118
rect 5426 25154 6495 25215
rect 5426 25120 5443 25154
rect 5477 25120 6443 25154
rect 6477 25120 6495 25154
rect 5426 25106 6495 25120
rect 6530 25154 7599 25215
rect 6530 25120 6547 25154
rect 6581 25120 7547 25154
rect 7581 25120 7599 25154
rect 6530 25106 7599 25120
rect 7634 25154 8703 25215
rect 7634 25120 7651 25154
rect 7685 25120 8651 25154
rect 8685 25120 8703 25154
rect 7634 25106 8703 25120
rect 8738 25154 9807 25215
rect 8738 25120 8755 25154
rect 8789 25120 9755 25154
rect 9789 25120 9807 25154
rect 8738 25106 9807 25120
rect 9841 25121 9899 25215
rect 4965 24991 5069 25065
rect 4965 24957 5015 24991
rect 5049 24957 5069 24991
rect 5103 24997 5123 25031
rect 5157 24997 5207 25031
rect 5103 24923 5207 24997
rect 4965 24876 5207 24923
rect 4965 24842 4983 24876
rect 5017 24842 5155 24876
rect 5189 24842 5207 24876
rect 4965 24781 5207 24842
rect 5744 25027 5814 25042
rect 5744 24993 5763 25027
rect 5797 24993 5814 25027
rect 5744 24792 5814 24993
rect 6110 24991 6178 25106
rect 6110 24957 6127 24991
rect 6161 24957 6178 24991
rect 6110 24940 6178 24957
rect 6848 25027 6918 25042
rect 6848 24993 6867 25027
rect 6901 24993 6918 25027
rect 6848 24792 6918 24993
rect 7214 24991 7282 25106
rect 7214 24957 7231 24991
rect 7265 24957 7282 24991
rect 7214 24940 7282 24957
rect 7952 25027 8022 25042
rect 7952 24993 7971 25027
rect 8005 24993 8022 25027
rect 7952 24792 8022 24993
rect 8318 24991 8386 25106
rect 8318 24957 8335 24991
rect 8369 24957 8386 24991
rect 8318 24940 8386 24957
rect 9056 25027 9126 25042
rect 9056 24993 9075 25027
rect 9109 24993 9126 25027
rect 9056 24792 9126 24993
rect 9422 24991 9490 25106
rect 9841 25087 9853 25121
rect 9887 25087 9899 25121
rect 9841 25070 9899 25087
rect 10025 25154 10543 25215
rect 10025 25120 10043 25154
rect 10077 25120 10491 25154
rect 10525 25120 10543 25154
rect 10025 25061 10543 25120
rect 10578 25154 11647 25215
rect 10578 25120 10595 25154
rect 10629 25120 11595 25154
rect 11629 25120 11647 25154
rect 10578 25106 11647 25120
rect 11682 25154 12751 25215
rect 11682 25120 11699 25154
rect 11733 25120 12699 25154
rect 12733 25120 12751 25154
rect 11682 25106 12751 25120
rect 12786 25154 13855 25215
rect 12786 25120 12803 25154
rect 12837 25120 13803 25154
rect 13837 25120 13855 25154
rect 12786 25106 13855 25120
rect 13890 25154 14959 25215
rect 13890 25120 13907 25154
rect 13941 25120 14907 25154
rect 14941 25120 14959 25154
rect 13890 25106 14959 25120
rect 14993 25121 15051 25215
rect 9422 24957 9439 24991
rect 9473 24957 9490 24991
rect 9422 24940 9490 24957
rect 10025 24993 10103 25027
rect 10137 24993 10213 25027
rect 10247 24993 10267 25027
rect 9841 24903 9899 24938
rect 9841 24869 9853 24903
rect 9887 24869 9899 24903
rect 9841 24810 9899 24869
rect 4965 24747 4983 24781
rect 5017 24747 5155 24781
rect 5189 24747 5207 24781
rect 4965 24705 5207 24747
rect 5426 24781 6495 24792
rect 5426 24747 5443 24781
rect 5477 24747 6443 24781
rect 6477 24747 6495 24781
rect 5426 24705 6495 24747
rect 6530 24781 7599 24792
rect 6530 24747 6547 24781
rect 6581 24747 7547 24781
rect 7581 24747 7599 24781
rect 6530 24705 7599 24747
rect 7634 24781 8703 24792
rect 7634 24747 7651 24781
rect 7685 24747 8651 24781
rect 8685 24747 8703 24781
rect 7634 24705 8703 24747
rect 8738 24781 9807 24792
rect 8738 24747 8755 24781
rect 8789 24747 9755 24781
rect 9789 24747 9807 24781
rect 8738 24705 9807 24747
rect 9841 24776 9853 24810
rect 9887 24776 9899 24810
rect 9841 24705 9899 24776
rect 10025 24923 10267 24993
rect 10301 24991 10543 25061
rect 10301 24957 10321 24991
rect 10355 24957 10431 24991
rect 10465 24957 10543 24991
rect 10896 25027 10966 25042
rect 10896 24993 10915 25027
rect 10949 24993 10966 25027
rect 10025 24883 10543 24923
rect 10025 24849 10043 24883
rect 10077 24849 10491 24883
rect 10525 24849 10543 24883
rect 10025 24781 10543 24849
rect 10896 24792 10966 24993
rect 11262 24991 11330 25106
rect 11262 24957 11279 24991
rect 11313 24957 11330 24991
rect 11262 24940 11330 24957
rect 12000 25027 12070 25042
rect 12000 24993 12019 25027
rect 12053 24993 12070 25027
rect 12000 24792 12070 24993
rect 12366 24991 12434 25106
rect 12366 24957 12383 24991
rect 12417 24957 12434 24991
rect 12366 24940 12434 24957
rect 13104 25027 13174 25042
rect 13104 24993 13123 25027
rect 13157 24993 13174 25027
rect 13104 24792 13174 24993
rect 13470 24991 13538 25106
rect 13470 24957 13487 24991
rect 13521 24957 13538 24991
rect 13470 24940 13538 24957
rect 14208 25027 14278 25042
rect 14208 24993 14227 25027
rect 14261 24993 14278 25027
rect 14208 24792 14278 24993
rect 14574 24991 14642 25106
rect 14993 25087 15005 25121
rect 15039 25087 15051 25121
rect 14993 25070 15051 25087
rect 15177 25147 15511 25215
rect 15177 25113 15195 25147
rect 15229 25113 15459 25147
rect 15493 25113 15511 25147
rect 15177 25061 15511 25113
rect 15546 25154 16615 25215
rect 15546 25120 15563 25154
rect 15597 25120 16563 25154
rect 16597 25120 16615 25154
rect 15546 25106 16615 25120
rect 16650 25154 17719 25215
rect 16650 25120 16667 25154
rect 16701 25120 17667 25154
rect 17701 25120 17719 25154
rect 16650 25106 17719 25120
rect 17754 25154 18823 25215
rect 17754 25120 17771 25154
rect 17805 25120 18771 25154
rect 18805 25120 18823 25154
rect 17754 25106 18823 25120
rect 18858 25154 19927 25215
rect 18858 25120 18875 25154
rect 18909 25120 19875 25154
rect 19909 25120 19927 25154
rect 18858 25106 19927 25120
rect 19961 25152 20203 25215
rect 19961 25118 19979 25152
rect 20013 25118 20151 25152
rect 20185 25118 20203 25152
rect 14574 24957 14591 24991
rect 14625 24957 14642 24991
rect 14574 24940 14642 24957
rect 15177 24993 15197 25027
rect 15231 24993 15327 25027
rect 14993 24903 15051 24938
rect 14993 24869 15005 24903
rect 15039 24869 15051 24903
rect 14993 24810 15051 24869
rect 10025 24747 10043 24781
rect 10077 24747 10491 24781
rect 10525 24747 10543 24781
rect 10025 24705 10543 24747
rect 10578 24781 11647 24792
rect 10578 24747 10595 24781
rect 10629 24747 11595 24781
rect 11629 24747 11647 24781
rect 10578 24705 11647 24747
rect 11682 24781 12751 24792
rect 11682 24747 11699 24781
rect 11733 24747 12699 24781
rect 12733 24747 12751 24781
rect 11682 24705 12751 24747
rect 12786 24781 13855 24792
rect 12786 24747 12803 24781
rect 12837 24747 13803 24781
rect 13837 24747 13855 24781
rect 12786 24705 13855 24747
rect 13890 24781 14959 24792
rect 13890 24747 13907 24781
rect 13941 24747 14907 24781
rect 14941 24747 14959 24781
rect 13890 24705 14959 24747
rect 14993 24776 15005 24810
rect 15039 24776 15051 24810
rect 14993 24705 15051 24776
rect 15177 24923 15327 24993
rect 15361 24991 15511 25061
rect 15361 24957 15457 24991
rect 15491 24957 15511 24991
rect 15864 25027 15934 25042
rect 15864 24993 15883 25027
rect 15917 24993 15934 25027
rect 15177 24883 15511 24923
rect 15177 24849 15195 24883
rect 15229 24849 15459 24883
rect 15493 24849 15511 24883
rect 15177 24781 15511 24849
rect 15864 24792 15934 24993
rect 16230 24991 16298 25106
rect 16230 24957 16247 24991
rect 16281 24957 16298 24991
rect 16230 24940 16298 24957
rect 16968 25027 17038 25042
rect 16968 24993 16987 25027
rect 17021 24993 17038 25027
rect 16968 24792 17038 24993
rect 17334 24991 17402 25106
rect 17334 24957 17351 24991
rect 17385 24957 17402 24991
rect 17334 24940 17402 24957
rect 18072 25027 18142 25042
rect 18072 24993 18091 25027
rect 18125 24993 18142 25027
rect 18072 24792 18142 24993
rect 18438 24991 18506 25106
rect 18438 24957 18455 24991
rect 18489 24957 18506 24991
rect 18438 24940 18506 24957
rect 19176 25027 19246 25042
rect 19176 24993 19195 25027
rect 19229 24993 19246 25027
rect 19176 24792 19246 24993
rect 19542 24991 19610 25106
rect 19961 25065 20203 25118
rect 19542 24957 19559 24991
rect 19593 24957 19610 24991
rect 19542 24940 19610 24957
rect 19961 24997 20011 25031
rect 20045 24997 20065 25031
rect 19961 24923 20065 24997
rect 20099 24991 20203 25065
rect 20099 24957 20119 24991
rect 20153 24957 20203 24991
rect 19961 24876 20203 24923
rect 19961 24842 19979 24876
rect 20013 24842 20151 24876
rect 20185 24842 20203 24876
rect 15177 24747 15195 24781
rect 15229 24747 15459 24781
rect 15493 24747 15511 24781
rect 15177 24705 15511 24747
rect 15546 24781 16615 24792
rect 15546 24747 15563 24781
rect 15597 24747 16563 24781
rect 16597 24747 16615 24781
rect 15546 24705 16615 24747
rect 16650 24781 17719 24792
rect 16650 24747 16667 24781
rect 16701 24747 17667 24781
rect 17701 24747 17719 24781
rect 16650 24705 17719 24747
rect 17754 24781 18823 24792
rect 17754 24747 17771 24781
rect 17805 24747 18771 24781
rect 18805 24747 18823 24781
rect 17754 24705 18823 24747
rect 18858 24781 19927 24792
rect 18858 24747 18875 24781
rect 18909 24747 19875 24781
rect 19909 24747 19927 24781
rect 18858 24705 19927 24747
rect 19961 24781 20203 24842
rect 19961 24747 19979 24781
rect 20013 24747 20151 24781
rect 20185 24747 20203 24781
rect 19961 24705 20203 24747
rect 4948 24671 4977 24705
rect 5011 24671 5069 24705
rect 5103 24671 5161 24705
rect 5195 24671 5253 24705
rect 5287 24671 5345 24705
rect 5379 24671 5437 24705
rect 5471 24671 5529 24705
rect 5563 24671 5621 24705
rect 5655 24671 5713 24705
rect 5747 24671 5805 24705
rect 5839 24671 5897 24705
rect 5931 24671 5989 24705
rect 6023 24671 6081 24705
rect 6115 24671 6173 24705
rect 6207 24671 6265 24705
rect 6299 24671 6357 24705
rect 6391 24671 6449 24705
rect 6483 24671 6541 24705
rect 6575 24671 6633 24705
rect 6667 24671 6725 24705
rect 6759 24671 6817 24705
rect 6851 24671 6909 24705
rect 6943 24671 7001 24705
rect 7035 24671 7093 24705
rect 7127 24671 7185 24705
rect 7219 24671 7277 24705
rect 7311 24671 7369 24705
rect 7403 24671 7461 24705
rect 7495 24671 7553 24705
rect 7587 24671 7645 24705
rect 7679 24671 7737 24705
rect 7771 24671 7829 24705
rect 7863 24671 7921 24705
rect 7955 24671 8013 24705
rect 8047 24671 8105 24705
rect 8139 24671 8197 24705
rect 8231 24671 8289 24705
rect 8323 24671 8381 24705
rect 8415 24671 8473 24705
rect 8507 24671 8565 24705
rect 8599 24671 8657 24705
rect 8691 24671 8749 24705
rect 8783 24671 8841 24705
rect 8875 24671 8933 24705
rect 8967 24671 9025 24705
rect 9059 24671 9117 24705
rect 9151 24671 9209 24705
rect 9243 24671 9301 24705
rect 9335 24671 9393 24705
rect 9427 24671 9485 24705
rect 9519 24671 9577 24705
rect 9611 24671 9669 24705
rect 9703 24671 9761 24705
rect 9795 24671 9853 24705
rect 9887 24671 9945 24705
rect 9979 24671 10037 24705
rect 10071 24671 10129 24705
rect 10163 24671 10221 24705
rect 10255 24671 10313 24705
rect 10347 24671 10405 24705
rect 10439 24671 10497 24705
rect 10531 24671 10589 24705
rect 10623 24671 10681 24705
rect 10715 24671 10773 24705
rect 10807 24671 10865 24705
rect 10899 24671 10957 24705
rect 10991 24671 11049 24705
rect 11083 24671 11141 24705
rect 11175 24671 11233 24705
rect 11267 24671 11325 24705
rect 11359 24671 11417 24705
rect 11451 24671 11509 24705
rect 11543 24671 11601 24705
rect 11635 24671 11693 24705
rect 11727 24671 11785 24705
rect 11819 24671 11877 24705
rect 11911 24671 11969 24705
rect 12003 24671 12061 24705
rect 12095 24671 12153 24705
rect 12187 24671 12245 24705
rect 12279 24671 12337 24705
rect 12371 24671 12429 24705
rect 12463 24671 12521 24705
rect 12555 24671 12613 24705
rect 12647 24671 12705 24705
rect 12739 24671 12797 24705
rect 12831 24671 12889 24705
rect 12923 24671 12981 24705
rect 13015 24671 13073 24705
rect 13107 24671 13165 24705
rect 13199 24671 13257 24705
rect 13291 24671 13349 24705
rect 13383 24671 13441 24705
rect 13475 24671 13533 24705
rect 13567 24671 13625 24705
rect 13659 24671 13717 24705
rect 13751 24671 13809 24705
rect 13843 24671 13901 24705
rect 13935 24671 13993 24705
rect 14027 24671 14085 24705
rect 14119 24671 14177 24705
rect 14211 24671 14269 24705
rect 14303 24671 14361 24705
rect 14395 24671 14453 24705
rect 14487 24671 14545 24705
rect 14579 24671 14637 24705
rect 14671 24671 14729 24705
rect 14763 24671 14821 24705
rect 14855 24671 14913 24705
rect 14947 24671 15005 24705
rect 15039 24671 15097 24705
rect 15131 24671 15189 24705
rect 15223 24671 15281 24705
rect 15315 24671 15373 24705
rect 15407 24671 15465 24705
rect 15499 24671 15557 24705
rect 15591 24671 15649 24705
rect 15683 24671 15741 24705
rect 15775 24671 15833 24705
rect 15867 24671 15925 24705
rect 15959 24671 16017 24705
rect 16051 24671 16109 24705
rect 16143 24671 16201 24705
rect 16235 24671 16293 24705
rect 16327 24671 16385 24705
rect 16419 24671 16477 24705
rect 16511 24671 16569 24705
rect 16603 24671 16661 24705
rect 16695 24671 16753 24705
rect 16787 24671 16845 24705
rect 16879 24671 16937 24705
rect 16971 24671 17029 24705
rect 17063 24671 17121 24705
rect 17155 24671 17213 24705
rect 17247 24671 17305 24705
rect 17339 24671 17397 24705
rect 17431 24671 17489 24705
rect 17523 24671 17581 24705
rect 17615 24671 17673 24705
rect 17707 24671 17765 24705
rect 17799 24671 17857 24705
rect 17891 24671 17949 24705
rect 17983 24671 18041 24705
rect 18075 24671 18133 24705
rect 18167 24671 18225 24705
rect 18259 24671 18317 24705
rect 18351 24671 18409 24705
rect 18443 24671 18501 24705
rect 18535 24671 18593 24705
rect 18627 24671 18685 24705
rect 18719 24671 18777 24705
rect 18811 24671 18869 24705
rect 18903 24671 18961 24705
rect 18995 24671 19053 24705
rect 19087 24671 19145 24705
rect 19179 24671 19237 24705
rect 19271 24671 19329 24705
rect 19363 24671 19421 24705
rect 19455 24671 19513 24705
rect 19547 24671 19605 24705
rect 19639 24671 19697 24705
rect 19731 24671 19789 24705
rect 19823 24671 19881 24705
rect 19915 24671 19973 24705
rect 20007 24671 20065 24705
rect 20099 24671 20157 24705
rect 20191 24671 20220 24705
rect 4965 24629 5207 24671
rect 4965 24595 4983 24629
rect 5017 24595 5155 24629
rect 5189 24595 5207 24629
rect 4965 24534 5207 24595
rect 4965 24500 4983 24534
rect 5017 24500 5155 24534
rect 5189 24500 5207 24534
rect 4965 24453 5207 24500
rect 4965 24385 5015 24419
rect 5049 24385 5069 24419
rect 4965 24311 5069 24385
rect 5103 24379 5207 24453
rect 5103 24345 5123 24379
rect 5157 24345 5207 24379
rect 5425 24629 6127 24671
rect 5425 24595 5443 24629
rect 5477 24595 6075 24629
rect 6109 24595 6127 24629
rect 5425 24527 6127 24595
rect 6162 24629 7231 24671
rect 6162 24595 6179 24629
rect 6213 24595 7179 24629
rect 7213 24595 7231 24629
rect 6162 24584 7231 24595
rect 7265 24600 7323 24671
rect 5425 24493 5443 24527
rect 5477 24493 6075 24527
rect 6109 24493 6127 24527
rect 5425 24453 6127 24493
rect 5425 24383 5763 24453
rect 5425 24349 5503 24383
rect 5537 24349 5606 24383
rect 5640 24349 5709 24383
rect 5743 24349 5763 24383
rect 5797 24385 5817 24419
rect 5851 24385 5916 24419
rect 5950 24385 6015 24419
rect 6049 24385 6127 24419
rect 5797 24315 6127 24385
rect 6480 24383 6550 24584
rect 7265 24566 7277 24600
rect 7311 24566 7323 24600
rect 7265 24507 7323 24566
rect 7265 24473 7277 24507
rect 7311 24473 7323 24507
rect 7265 24438 7323 24473
rect 7449 24629 7967 24671
rect 7449 24595 7467 24629
rect 7501 24595 7915 24629
rect 7949 24595 7967 24629
rect 7449 24527 7967 24595
rect 8002 24629 9071 24671
rect 8002 24595 8019 24629
rect 8053 24595 9019 24629
rect 9053 24595 9071 24629
rect 8002 24584 9071 24595
rect 9106 24629 10175 24671
rect 9106 24595 9123 24629
rect 9157 24595 10123 24629
rect 10157 24595 10175 24629
rect 9106 24584 10175 24595
rect 10210 24629 11279 24671
rect 10210 24595 10227 24629
rect 10261 24595 11227 24629
rect 11261 24595 11279 24629
rect 10210 24584 11279 24595
rect 11314 24629 12383 24671
rect 11314 24595 11331 24629
rect 11365 24595 12331 24629
rect 12365 24595 12383 24629
rect 11314 24584 12383 24595
rect 12417 24600 12475 24671
rect 7449 24493 7467 24527
rect 7501 24493 7915 24527
rect 7949 24493 7967 24527
rect 7449 24453 7967 24493
rect 6480 24349 6499 24383
rect 6533 24349 6550 24383
rect 6480 24334 6550 24349
rect 6846 24419 6914 24436
rect 6846 24385 6863 24419
rect 6897 24385 6914 24419
rect 4965 24258 5207 24311
rect 4965 24224 4983 24258
rect 5017 24224 5155 24258
rect 5189 24224 5207 24258
rect 4965 24161 5207 24224
rect 5425 24256 6127 24315
rect 6846 24270 6914 24385
rect 7449 24383 7691 24453
rect 7449 24349 7527 24383
rect 7561 24349 7637 24383
rect 7671 24349 7691 24383
rect 7725 24385 7745 24419
rect 7779 24385 7855 24419
rect 7889 24385 7967 24419
rect 7725 24315 7967 24385
rect 8320 24383 8390 24584
rect 8320 24349 8339 24383
rect 8373 24349 8390 24383
rect 8320 24334 8390 24349
rect 8686 24419 8754 24436
rect 8686 24385 8703 24419
rect 8737 24385 8754 24419
rect 7265 24289 7323 24306
rect 5425 24222 5443 24256
rect 5477 24222 6075 24256
rect 6109 24222 6127 24256
rect 5425 24161 6127 24222
rect 6162 24256 7231 24270
rect 6162 24222 6179 24256
rect 6213 24222 7179 24256
rect 7213 24222 7231 24256
rect 6162 24161 7231 24222
rect 7265 24255 7277 24289
rect 7311 24255 7323 24289
rect 7265 24161 7323 24255
rect 7449 24256 7967 24315
rect 8686 24270 8754 24385
rect 9424 24383 9494 24584
rect 9424 24349 9443 24383
rect 9477 24349 9494 24383
rect 9424 24334 9494 24349
rect 9790 24419 9858 24436
rect 9790 24385 9807 24419
rect 9841 24385 9858 24419
rect 9790 24270 9858 24385
rect 10528 24383 10598 24584
rect 10528 24349 10547 24383
rect 10581 24349 10598 24383
rect 10528 24334 10598 24349
rect 10894 24419 10962 24436
rect 10894 24385 10911 24419
rect 10945 24385 10962 24419
rect 10894 24270 10962 24385
rect 11632 24383 11702 24584
rect 12417 24566 12429 24600
rect 12463 24566 12475 24600
rect 12417 24507 12475 24566
rect 12417 24473 12429 24507
rect 12463 24473 12475 24507
rect 12417 24438 12475 24473
rect 12601 24629 13119 24671
rect 12601 24595 12619 24629
rect 12653 24595 13067 24629
rect 13101 24595 13119 24629
rect 12601 24527 13119 24595
rect 13154 24629 14223 24671
rect 13154 24595 13171 24629
rect 13205 24595 14171 24629
rect 14205 24595 14223 24629
rect 13154 24584 14223 24595
rect 14258 24629 15327 24671
rect 14258 24595 14275 24629
rect 14309 24595 15275 24629
rect 15309 24595 15327 24629
rect 14258 24584 15327 24595
rect 15362 24629 16431 24671
rect 15362 24595 15379 24629
rect 15413 24595 16379 24629
rect 16413 24595 16431 24629
rect 15362 24584 16431 24595
rect 16466 24629 17535 24671
rect 16466 24595 16483 24629
rect 16517 24595 17483 24629
rect 17517 24595 17535 24629
rect 16466 24584 17535 24595
rect 17569 24600 17627 24671
rect 12601 24493 12619 24527
rect 12653 24493 13067 24527
rect 13101 24493 13119 24527
rect 12601 24453 13119 24493
rect 11632 24349 11651 24383
rect 11685 24349 11702 24383
rect 11632 24334 11702 24349
rect 11998 24419 12066 24436
rect 11998 24385 12015 24419
rect 12049 24385 12066 24419
rect 11998 24270 12066 24385
rect 12601 24383 12843 24453
rect 12601 24349 12679 24383
rect 12713 24349 12789 24383
rect 12823 24349 12843 24383
rect 12877 24385 12897 24419
rect 12931 24385 13007 24419
rect 13041 24385 13119 24419
rect 12877 24315 13119 24385
rect 13472 24383 13542 24584
rect 13472 24349 13491 24383
rect 13525 24349 13542 24383
rect 13472 24334 13542 24349
rect 13838 24419 13906 24436
rect 13838 24385 13855 24419
rect 13889 24385 13906 24419
rect 12417 24289 12475 24306
rect 7449 24222 7467 24256
rect 7501 24222 7915 24256
rect 7949 24222 7967 24256
rect 7449 24161 7967 24222
rect 8002 24256 9071 24270
rect 8002 24222 8019 24256
rect 8053 24222 9019 24256
rect 9053 24222 9071 24256
rect 8002 24161 9071 24222
rect 9106 24256 10175 24270
rect 9106 24222 9123 24256
rect 9157 24222 10123 24256
rect 10157 24222 10175 24256
rect 9106 24161 10175 24222
rect 10210 24256 11279 24270
rect 10210 24222 10227 24256
rect 10261 24222 11227 24256
rect 11261 24222 11279 24256
rect 10210 24161 11279 24222
rect 11314 24256 12383 24270
rect 11314 24222 11331 24256
rect 11365 24222 12331 24256
rect 12365 24222 12383 24256
rect 11314 24161 12383 24222
rect 12417 24255 12429 24289
rect 12463 24255 12475 24289
rect 12417 24161 12475 24255
rect 12601 24256 13119 24315
rect 13838 24270 13906 24385
rect 14576 24383 14646 24584
rect 14576 24349 14595 24383
rect 14629 24349 14646 24383
rect 14576 24334 14646 24349
rect 14942 24419 15010 24436
rect 14942 24385 14959 24419
rect 14993 24385 15010 24419
rect 14942 24270 15010 24385
rect 15680 24383 15750 24584
rect 15680 24349 15699 24383
rect 15733 24349 15750 24383
rect 15680 24334 15750 24349
rect 16046 24419 16114 24436
rect 16046 24385 16063 24419
rect 16097 24385 16114 24419
rect 16046 24270 16114 24385
rect 16784 24383 16854 24584
rect 17569 24566 17581 24600
rect 17615 24566 17627 24600
rect 17754 24629 18823 24671
rect 17754 24595 17771 24629
rect 17805 24595 18771 24629
rect 18805 24595 18823 24629
rect 17754 24584 18823 24595
rect 18858 24629 19927 24671
rect 18858 24595 18875 24629
rect 18909 24595 19875 24629
rect 19909 24595 19927 24629
rect 18858 24584 19927 24595
rect 19961 24629 20203 24671
rect 19961 24595 19979 24629
rect 20013 24595 20151 24629
rect 20185 24595 20203 24629
rect 17569 24507 17627 24566
rect 17569 24473 17581 24507
rect 17615 24473 17627 24507
rect 17569 24438 17627 24473
rect 16784 24349 16803 24383
rect 16837 24349 16854 24383
rect 16784 24334 16854 24349
rect 17150 24419 17218 24436
rect 17150 24385 17167 24419
rect 17201 24385 17218 24419
rect 17150 24270 17218 24385
rect 18072 24383 18142 24584
rect 18072 24349 18091 24383
rect 18125 24349 18142 24383
rect 18072 24334 18142 24349
rect 18438 24419 18506 24436
rect 18438 24385 18455 24419
rect 18489 24385 18506 24419
rect 17569 24289 17627 24306
rect 12601 24222 12619 24256
rect 12653 24222 13067 24256
rect 13101 24222 13119 24256
rect 12601 24161 13119 24222
rect 13154 24256 14223 24270
rect 13154 24222 13171 24256
rect 13205 24222 14171 24256
rect 14205 24222 14223 24256
rect 13154 24161 14223 24222
rect 14258 24256 15327 24270
rect 14258 24222 14275 24256
rect 14309 24222 15275 24256
rect 15309 24222 15327 24256
rect 14258 24161 15327 24222
rect 15362 24256 16431 24270
rect 15362 24222 15379 24256
rect 15413 24222 16379 24256
rect 16413 24222 16431 24256
rect 15362 24161 16431 24222
rect 16466 24256 17535 24270
rect 16466 24222 16483 24256
rect 16517 24222 17483 24256
rect 17517 24222 17535 24256
rect 16466 24161 17535 24222
rect 17569 24255 17581 24289
rect 17615 24255 17627 24289
rect 18438 24270 18506 24385
rect 19176 24383 19246 24584
rect 19961 24534 20203 24595
rect 19961 24500 19979 24534
rect 20013 24500 20151 24534
rect 20185 24500 20203 24534
rect 19961 24453 20203 24500
rect 19176 24349 19195 24383
rect 19229 24349 19246 24383
rect 19176 24334 19246 24349
rect 19542 24419 19610 24436
rect 19542 24385 19559 24419
rect 19593 24385 19610 24419
rect 19542 24270 19610 24385
rect 19961 24379 20065 24453
rect 19961 24345 20011 24379
rect 20045 24345 20065 24379
rect 20099 24385 20119 24419
rect 20153 24385 20203 24419
rect 20099 24311 20203 24385
rect 17569 24161 17627 24255
rect 17754 24256 18823 24270
rect 17754 24222 17771 24256
rect 17805 24222 18771 24256
rect 18805 24222 18823 24256
rect 17754 24161 18823 24222
rect 18858 24256 19927 24270
rect 18858 24222 18875 24256
rect 18909 24222 19875 24256
rect 19909 24222 19927 24256
rect 18858 24161 19927 24222
rect 19961 24258 20203 24311
rect 19961 24224 19979 24258
rect 20013 24224 20151 24258
rect 20185 24224 20203 24258
rect 19961 24161 20203 24224
rect 4948 24127 4977 24161
rect 5011 24127 5069 24161
rect 5103 24127 5161 24161
rect 5195 24127 5253 24161
rect 5287 24127 5345 24161
rect 5379 24127 5437 24161
rect 5471 24127 5529 24161
rect 5563 24127 5621 24161
rect 5655 24127 5713 24161
rect 5747 24127 5805 24161
rect 5839 24127 5897 24161
rect 5931 24127 5989 24161
rect 6023 24127 6081 24161
rect 6115 24127 6173 24161
rect 6207 24127 6265 24161
rect 6299 24127 6357 24161
rect 6391 24127 6449 24161
rect 6483 24127 6541 24161
rect 6575 24127 6633 24161
rect 6667 24127 6725 24161
rect 6759 24127 6817 24161
rect 6851 24127 6909 24161
rect 6943 24127 7001 24161
rect 7035 24127 7093 24161
rect 7127 24127 7185 24161
rect 7219 24127 7277 24161
rect 7311 24127 7369 24161
rect 7403 24127 7461 24161
rect 7495 24127 7553 24161
rect 7587 24127 7645 24161
rect 7679 24127 7737 24161
rect 7771 24127 7829 24161
rect 7863 24127 7921 24161
rect 7955 24127 8013 24161
rect 8047 24127 8105 24161
rect 8139 24127 8197 24161
rect 8231 24127 8289 24161
rect 8323 24127 8381 24161
rect 8415 24127 8473 24161
rect 8507 24127 8565 24161
rect 8599 24127 8657 24161
rect 8691 24127 8749 24161
rect 8783 24127 8841 24161
rect 8875 24127 8933 24161
rect 8967 24127 9025 24161
rect 9059 24127 9117 24161
rect 9151 24127 9209 24161
rect 9243 24127 9301 24161
rect 9335 24127 9393 24161
rect 9427 24127 9485 24161
rect 9519 24127 9577 24161
rect 9611 24127 9669 24161
rect 9703 24127 9761 24161
rect 9795 24127 9853 24161
rect 9887 24127 9945 24161
rect 9979 24127 10037 24161
rect 10071 24127 10129 24161
rect 10163 24127 10221 24161
rect 10255 24127 10313 24161
rect 10347 24127 10405 24161
rect 10439 24127 10497 24161
rect 10531 24127 10589 24161
rect 10623 24127 10681 24161
rect 10715 24127 10773 24161
rect 10807 24127 10865 24161
rect 10899 24127 10957 24161
rect 10991 24127 11049 24161
rect 11083 24127 11141 24161
rect 11175 24127 11233 24161
rect 11267 24127 11325 24161
rect 11359 24127 11417 24161
rect 11451 24127 11509 24161
rect 11543 24127 11601 24161
rect 11635 24127 11693 24161
rect 11727 24127 11785 24161
rect 11819 24127 11877 24161
rect 11911 24127 11969 24161
rect 12003 24127 12061 24161
rect 12095 24127 12153 24161
rect 12187 24127 12245 24161
rect 12279 24127 12337 24161
rect 12371 24127 12429 24161
rect 12463 24127 12521 24161
rect 12555 24127 12613 24161
rect 12647 24127 12705 24161
rect 12739 24127 12797 24161
rect 12831 24127 12889 24161
rect 12923 24127 12981 24161
rect 13015 24127 13073 24161
rect 13107 24127 13165 24161
rect 13199 24127 13257 24161
rect 13291 24127 13349 24161
rect 13383 24127 13441 24161
rect 13475 24127 13533 24161
rect 13567 24127 13625 24161
rect 13659 24127 13717 24161
rect 13751 24127 13809 24161
rect 13843 24127 13901 24161
rect 13935 24127 13993 24161
rect 14027 24127 14085 24161
rect 14119 24127 14177 24161
rect 14211 24127 14269 24161
rect 14303 24127 14361 24161
rect 14395 24127 14453 24161
rect 14487 24127 14545 24161
rect 14579 24127 14637 24161
rect 14671 24127 14729 24161
rect 14763 24127 14821 24161
rect 14855 24127 14913 24161
rect 14947 24127 15005 24161
rect 15039 24127 15097 24161
rect 15131 24127 15189 24161
rect 15223 24127 15281 24161
rect 15315 24127 15373 24161
rect 15407 24127 15465 24161
rect 15499 24127 15557 24161
rect 15591 24127 15649 24161
rect 15683 24127 15741 24161
rect 15775 24127 15833 24161
rect 15867 24127 15925 24161
rect 15959 24127 16017 24161
rect 16051 24127 16109 24161
rect 16143 24127 16201 24161
rect 16235 24127 16293 24161
rect 16327 24127 16385 24161
rect 16419 24127 16477 24161
rect 16511 24127 16569 24161
rect 16603 24127 16661 24161
rect 16695 24127 16753 24161
rect 16787 24127 16845 24161
rect 16879 24127 16937 24161
rect 16971 24127 17029 24161
rect 17063 24127 17121 24161
rect 17155 24127 17213 24161
rect 17247 24127 17305 24161
rect 17339 24127 17397 24161
rect 17431 24127 17489 24161
rect 17523 24127 17581 24161
rect 17615 24127 17673 24161
rect 17707 24127 17765 24161
rect 17799 24127 17857 24161
rect 17891 24127 17949 24161
rect 17983 24127 18041 24161
rect 18075 24127 18133 24161
rect 18167 24127 18225 24161
rect 18259 24127 18317 24161
rect 18351 24127 18409 24161
rect 18443 24127 18501 24161
rect 18535 24127 18593 24161
rect 18627 24127 18685 24161
rect 18719 24127 18777 24161
rect 18811 24127 18869 24161
rect 18903 24127 18961 24161
rect 18995 24127 19053 24161
rect 19087 24127 19145 24161
rect 19179 24127 19237 24161
rect 19271 24127 19329 24161
rect 19363 24127 19421 24161
rect 19455 24127 19513 24161
rect 19547 24127 19605 24161
rect 19639 24127 19697 24161
rect 19731 24127 19789 24161
rect 19823 24127 19881 24161
rect 19915 24127 19973 24161
rect 20007 24127 20065 24161
rect 20099 24127 20157 24161
rect 20191 24127 20220 24161
rect 4965 24064 5207 24127
rect 4965 24030 4983 24064
rect 5017 24030 5155 24064
rect 5189 24030 5207 24064
rect 4965 23977 5207 24030
rect 5426 24066 6495 24127
rect 5426 24032 5443 24066
rect 5477 24032 6443 24066
rect 6477 24032 6495 24066
rect 5426 24018 6495 24032
rect 6530 24066 7599 24127
rect 6530 24032 6547 24066
rect 6581 24032 7547 24066
rect 7581 24032 7599 24066
rect 6530 24018 7599 24032
rect 7634 24066 8703 24127
rect 7634 24032 7651 24066
rect 7685 24032 8651 24066
rect 8685 24032 8703 24066
rect 7634 24018 8703 24032
rect 8738 24066 9807 24127
rect 8738 24032 8755 24066
rect 8789 24032 9755 24066
rect 9789 24032 9807 24066
rect 8738 24018 9807 24032
rect 9841 24033 9899 24127
rect 4965 23903 5069 23977
rect 4965 23869 5015 23903
rect 5049 23869 5069 23903
rect 5103 23909 5123 23943
rect 5157 23909 5207 23943
rect 5103 23835 5207 23909
rect 4965 23788 5207 23835
rect 4965 23754 4983 23788
rect 5017 23754 5155 23788
rect 5189 23754 5207 23788
rect 4965 23693 5207 23754
rect 5744 23939 5814 23954
rect 5744 23905 5763 23939
rect 5797 23905 5814 23939
rect 5744 23704 5814 23905
rect 6110 23903 6178 24018
rect 6110 23869 6127 23903
rect 6161 23869 6178 23903
rect 6110 23852 6178 23869
rect 6848 23939 6918 23954
rect 6848 23905 6867 23939
rect 6901 23905 6918 23939
rect 6848 23704 6918 23905
rect 7214 23903 7282 24018
rect 7214 23869 7231 23903
rect 7265 23869 7282 23903
rect 7214 23852 7282 23869
rect 7952 23939 8022 23954
rect 7952 23905 7971 23939
rect 8005 23905 8022 23939
rect 7952 23704 8022 23905
rect 8318 23903 8386 24018
rect 8318 23869 8335 23903
rect 8369 23869 8386 23903
rect 8318 23852 8386 23869
rect 9056 23939 9126 23954
rect 9056 23905 9075 23939
rect 9109 23905 9126 23939
rect 9056 23704 9126 23905
rect 9422 23903 9490 24018
rect 9841 23999 9853 24033
rect 9887 23999 9899 24033
rect 9841 23982 9899 23999
rect 10025 24066 10543 24127
rect 10025 24032 10043 24066
rect 10077 24032 10491 24066
rect 10525 24032 10543 24066
rect 10025 23973 10543 24032
rect 10578 24066 11647 24127
rect 10578 24032 10595 24066
rect 10629 24032 11595 24066
rect 11629 24032 11647 24066
rect 10578 24018 11647 24032
rect 11682 24066 12751 24127
rect 11682 24032 11699 24066
rect 11733 24032 12699 24066
rect 12733 24032 12751 24066
rect 11682 24018 12751 24032
rect 12786 24066 13855 24127
rect 12786 24032 12803 24066
rect 12837 24032 13803 24066
rect 13837 24032 13855 24066
rect 12786 24018 13855 24032
rect 13890 24066 14959 24127
rect 13890 24032 13907 24066
rect 13941 24032 14907 24066
rect 14941 24032 14959 24066
rect 13890 24018 14959 24032
rect 14993 24033 15051 24127
rect 9422 23869 9439 23903
rect 9473 23869 9490 23903
rect 9422 23852 9490 23869
rect 10025 23905 10103 23939
rect 10137 23905 10213 23939
rect 10247 23905 10267 23939
rect 9841 23815 9899 23850
rect 9841 23781 9853 23815
rect 9887 23781 9899 23815
rect 9841 23722 9899 23781
rect 4965 23659 4983 23693
rect 5017 23659 5155 23693
rect 5189 23659 5207 23693
rect 4965 23617 5207 23659
rect 5426 23693 6495 23704
rect 5426 23659 5443 23693
rect 5477 23659 6443 23693
rect 6477 23659 6495 23693
rect 5426 23617 6495 23659
rect 6530 23693 7599 23704
rect 6530 23659 6547 23693
rect 6581 23659 7547 23693
rect 7581 23659 7599 23693
rect 6530 23617 7599 23659
rect 7634 23693 8703 23704
rect 7634 23659 7651 23693
rect 7685 23659 8651 23693
rect 8685 23659 8703 23693
rect 7634 23617 8703 23659
rect 8738 23693 9807 23704
rect 8738 23659 8755 23693
rect 8789 23659 9755 23693
rect 9789 23659 9807 23693
rect 8738 23617 9807 23659
rect 9841 23688 9853 23722
rect 9887 23688 9899 23722
rect 9841 23617 9899 23688
rect 10025 23835 10267 23905
rect 10301 23903 10543 23973
rect 10301 23869 10321 23903
rect 10355 23869 10431 23903
rect 10465 23869 10543 23903
rect 10896 23939 10966 23954
rect 10896 23905 10915 23939
rect 10949 23905 10966 23939
rect 10025 23795 10543 23835
rect 10025 23761 10043 23795
rect 10077 23761 10491 23795
rect 10525 23761 10543 23795
rect 10025 23693 10543 23761
rect 10896 23704 10966 23905
rect 11262 23903 11330 24018
rect 11262 23869 11279 23903
rect 11313 23869 11330 23903
rect 11262 23852 11330 23869
rect 12000 23939 12070 23954
rect 12000 23905 12019 23939
rect 12053 23905 12070 23939
rect 12000 23704 12070 23905
rect 12366 23903 12434 24018
rect 12366 23869 12383 23903
rect 12417 23869 12434 23903
rect 12366 23852 12434 23869
rect 13104 23939 13174 23954
rect 13104 23905 13123 23939
rect 13157 23905 13174 23939
rect 13104 23704 13174 23905
rect 13470 23903 13538 24018
rect 13470 23869 13487 23903
rect 13521 23869 13538 23903
rect 13470 23852 13538 23869
rect 14208 23939 14278 23954
rect 14208 23905 14227 23939
rect 14261 23905 14278 23939
rect 14208 23704 14278 23905
rect 14574 23903 14642 24018
rect 14993 23999 15005 24033
rect 15039 23999 15051 24033
rect 14993 23982 15051 23999
rect 15177 24059 15511 24127
rect 15177 24025 15195 24059
rect 15229 24025 15459 24059
rect 15493 24025 15511 24059
rect 15177 23973 15511 24025
rect 15546 24066 16615 24127
rect 15546 24032 15563 24066
rect 15597 24032 16563 24066
rect 16597 24032 16615 24066
rect 15546 24018 16615 24032
rect 16650 24066 17719 24127
rect 16650 24032 16667 24066
rect 16701 24032 17667 24066
rect 17701 24032 17719 24066
rect 16650 24018 17719 24032
rect 17754 24066 18823 24127
rect 17754 24032 17771 24066
rect 17805 24032 18771 24066
rect 18805 24032 18823 24066
rect 17754 24018 18823 24032
rect 18858 24066 19927 24127
rect 18858 24032 18875 24066
rect 18909 24032 19875 24066
rect 19909 24032 19927 24066
rect 18858 24018 19927 24032
rect 19961 24064 20203 24127
rect 19961 24030 19979 24064
rect 20013 24030 20151 24064
rect 20185 24030 20203 24064
rect 14574 23869 14591 23903
rect 14625 23869 14642 23903
rect 14574 23852 14642 23869
rect 15177 23905 15197 23939
rect 15231 23905 15327 23939
rect 14993 23815 15051 23850
rect 14993 23781 15005 23815
rect 15039 23781 15051 23815
rect 14993 23722 15051 23781
rect 10025 23659 10043 23693
rect 10077 23659 10491 23693
rect 10525 23659 10543 23693
rect 10025 23617 10543 23659
rect 10578 23693 11647 23704
rect 10578 23659 10595 23693
rect 10629 23659 11595 23693
rect 11629 23659 11647 23693
rect 10578 23617 11647 23659
rect 11682 23693 12751 23704
rect 11682 23659 11699 23693
rect 11733 23659 12699 23693
rect 12733 23659 12751 23693
rect 11682 23617 12751 23659
rect 12786 23693 13855 23704
rect 12786 23659 12803 23693
rect 12837 23659 13803 23693
rect 13837 23659 13855 23693
rect 12786 23617 13855 23659
rect 13890 23693 14959 23704
rect 13890 23659 13907 23693
rect 13941 23659 14907 23693
rect 14941 23659 14959 23693
rect 13890 23617 14959 23659
rect 14993 23688 15005 23722
rect 15039 23688 15051 23722
rect 14993 23617 15051 23688
rect 15177 23835 15327 23905
rect 15361 23903 15511 23973
rect 15361 23869 15457 23903
rect 15491 23869 15511 23903
rect 15864 23939 15934 23954
rect 15864 23905 15883 23939
rect 15917 23905 15934 23939
rect 15177 23795 15511 23835
rect 15177 23761 15195 23795
rect 15229 23761 15459 23795
rect 15493 23761 15511 23795
rect 15177 23693 15511 23761
rect 15864 23704 15934 23905
rect 16230 23903 16298 24018
rect 16230 23869 16247 23903
rect 16281 23869 16298 23903
rect 16230 23852 16298 23869
rect 16968 23939 17038 23954
rect 16968 23905 16987 23939
rect 17021 23905 17038 23939
rect 16968 23704 17038 23905
rect 17334 23903 17402 24018
rect 17334 23869 17351 23903
rect 17385 23869 17402 23903
rect 17334 23852 17402 23869
rect 18072 23939 18142 23954
rect 18072 23905 18091 23939
rect 18125 23905 18142 23939
rect 18072 23704 18142 23905
rect 18438 23903 18506 24018
rect 18438 23869 18455 23903
rect 18489 23869 18506 23903
rect 18438 23852 18506 23869
rect 19176 23939 19246 23954
rect 19176 23905 19195 23939
rect 19229 23905 19246 23939
rect 19176 23704 19246 23905
rect 19542 23903 19610 24018
rect 19961 23977 20203 24030
rect 19542 23869 19559 23903
rect 19593 23869 19610 23903
rect 19542 23852 19610 23869
rect 19961 23909 20011 23943
rect 20045 23909 20065 23943
rect 19961 23835 20065 23909
rect 20099 23903 20203 23977
rect 20099 23869 20119 23903
rect 20153 23869 20203 23903
rect 19961 23788 20203 23835
rect 19961 23754 19979 23788
rect 20013 23754 20151 23788
rect 20185 23754 20203 23788
rect 15177 23659 15195 23693
rect 15229 23659 15459 23693
rect 15493 23659 15511 23693
rect 15177 23617 15511 23659
rect 15546 23693 16615 23704
rect 15546 23659 15563 23693
rect 15597 23659 16563 23693
rect 16597 23659 16615 23693
rect 15546 23617 16615 23659
rect 16650 23693 17719 23704
rect 16650 23659 16667 23693
rect 16701 23659 17667 23693
rect 17701 23659 17719 23693
rect 16650 23617 17719 23659
rect 17754 23693 18823 23704
rect 17754 23659 17771 23693
rect 17805 23659 18771 23693
rect 18805 23659 18823 23693
rect 17754 23617 18823 23659
rect 18858 23693 19927 23704
rect 18858 23659 18875 23693
rect 18909 23659 19875 23693
rect 19909 23659 19927 23693
rect 18858 23617 19927 23659
rect 19961 23693 20203 23754
rect 19961 23659 19979 23693
rect 20013 23659 20151 23693
rect 20185 23659 20203 23693
rect 19961 23617 20203 23659
rect 4948 23583 4977 23617
rect 5011 23583 5069 23617
rect 5103 23583 5161 23617
rect 5195 23583 5253 23617
rect 5287 23583 5345 23617
rect 5379 23583 5437 23617
rect 5471 23583 5529 23617
rect 5563 23583 5621 23617
rect 5655 23583 5713 23617
rect 5747 23583 5805 23617
rect 5839 23583 5897 23617
rect 5931 23583 5989 23617
rect 6023 23583 6081 23617
rect 6115 23583 6173 23617
rect 6207 23583 6265 23617
rect 6299 23583 6357 23617
rect 6391 23583 6449 23617
rect 6483 23583 6541 23617
rect 6575 23583 6633 23617
rect 6667 23583 6725 23617
rect 6759 23583 6817 23617
rect 6851 23583 6909 23617
rect 6943 23583 7001 23617
rect 7035 23583 7093 23617
rect 7127 23583 7185 23617
rect 7219 23583 7277 23617
rect 7311 23583 7369 23617
rect 7403 23583 7461 23617
rect 7495 23583 7553 23617
rect 7587 23583 7645 23617
rect 7679 23583 7737 23617
rect 7771 23583 7829 23617
rect 7863 23583 7921 23617
rect 7955 23583 8013 23617
rect 8047 23583 8105 23617
rect 8139 23583 8197 23617
rect 8231 23583 8289 23617
rect 8323 23583 8381 23617
rect 8415 23583 8473 23617
rect 8507 23583 8565 23617
rect 8599 23583 8657 23617
rect 8691 23583 8749 23617
rect 8783 23583 8841 23617
rect 8875 23583 8933 23617
rect 8967 23583 9025 23617
rect 9059 23583 9117 23617
rect 9151 23583 9209 23617
rect 9243 23583 9301 23617
rect 9335 23583 9393 23617
rect 9427 23583 9485 23617
rect 9519 23583 9577 23617
rect 9611 23583 9669 23617
rect 9703 23583 9761 23617
rect 9795 23583 9853 23617
rect 9887 23583 9945 23617
rect 9979 23583 10037 23617
rect 10071 23583 10129 23617
rect 10163 23583 10221 23617
rect 10255 23583 10313 23617
rect 10347 23583 10405 23617
rect 10439 23583 10497 23617
rect 10531 23583 10589 23617
rect 10623 23583 10681 23617
rect 10715 23583 10773 23617
rect 10807 23583 10865 23617
rect 10899 23583 10957 23617
rect 10991 23583 11049 23617
rect 11083 23583 11141 23617
rect 11175 23583 11233 23617
rect 11267 23583 11325 23617
rect 11359 23583 11417 23617
rect 11451 23583 11509 23617
rect 11543 23583 11601 23617
rect 11635 23583 11693 23617
rect 11727 23583 11785 23617
rect 11819 23583 11877 23617
rect 11911 23583 11969 23617
rect 12003 23583 12061 23617
rect 12095 23583 12153 23617
rect 12187 23583 12245 23617
rect 12279 23583 12337 23617
rect 12371 23583 12429 23617
rect 12463 23583 12521 23617
rect 12555 23583 12613 23617
rect 12647 23583 12705 23617
rect 12739 23583 12797 23617
rect 12831 23583 12889 23617
rect 12923 23583 12981 23617
rect 13015 23583 13073 23617
rect 13107 23583 13165 23617
rect 13199 23583 13257 23617
rect 13291 23583 13349 23617
rect 13383 23583 13441 23617
rect 13475 23583 13533 23617
rect 13567 23583 13625 23617
rect 13659 23583 13717 23617
rect 13751 23583 13809 23617
rect 13843 23583 13901 23617
rect 13935 23583 13993 23617
rect 14027 23583 14085 23617
rect 14119 23583 14177 23617
rect 14211 23583 14269 23617
rect 14303 23583 14361 23617
rect 14395 23583 14453 23617
rect 14487 23583 14545 23617
rect 14579 23583 14637 23617
rect 14671 23583 14729 23617
rect 14763 23583 14821 23617
rect 14855 23583 14913 23617
rect 14947 23583 15005 23617
rect 15039 23583 15097 23617
rect 15131 23583 15189 23617
rect 15223 23583 15281 23617
rect 15315 23583 15373 23617
rect 15407 23583 15465 23617
rect 15499 23583 15557 23617
rect 15591 23583 15649 23617
rect 15683 23583 15741 23617
rect 15775 23583 15833 23617
rect 15867 23583 15925 23617
rect 15959 23583 16017 23617
rect 16051 23583 16109 23617
rect 16143 23583 16201 23617
rect 16235 23583 16293 23617
rect 16327 23583 16385 23617
rect 16419 23583 16477 23617
rect 16511 23583 16569 23617
rect 16603 23583 16661 23617
rect 16695 23583 16753 23617
rect 16787 23583 16845 23617
rect 16879 23583 16937 23617
rect 16971 23583 17029 23617
rect 17063 23583 17121 23617
rect 17155 23583 17213 23617
rect 17247 23583 17305 23617
rect 17339 23583 17397 23617
rect 17431 23583 17489 23617
rect 17523 23583 17581 23617
rect 17615 23583 17673 23617
rect 17707 23583 17765 23617
rect 17799 23583 17857 23617
rect 17891 23583 17949 23617
rect 17983 23583 18041 23617
rect 18075 23583 18133 23617
rect 18167 23583 18225 23617
rect 18259 23583 18317 23617
rect 18351 23583 18409 23617
rect 18443 23583 18501 23617
rect 18535 23583 18593 23617
rect 18627 23583 18685 23617
rect 18719 23583 18777 23617
rect 18811 23583 18869 23617
rect 18903 23583 18961 23617
rect 18995 23583 19053 23617
rect 19087 23583 19145 23617
rect 19179 23583 19237 23617
rect 19271 23583 19329 23617
rect 19363 23583 19421 23617
rect 19455 23583 19513 23617
rect 19547 23583 19605 23617
rect 19639 23583 19697 23617
rect 19731 23583 19789 23617
rect 19823 23583 19881 23617
rect 19915 23583 19973 23617
rect 20007 23583 20065 23617
rect 20099 23583 20157 23617
rect 20191 23583 20220 23617
rect 4965 23541 5207 23583
rect 4965 23507 4983 23541
rect 5017 23507 5155 23541
rect 5189 23507 5207 23541
rect 4965 23446 5207 23507
rect 4965 23412 4983 23446
rect 5017 23412 5155 23446
rect 5189 23412 5207 23446
rect 4965 23365 5207 23412
rect 4965 23297 5015 23331
rect 5049 23297 5069 23331
rect 4965 23223 5069 23297
rect 5103 23291 5207 23365
rect 5103 23257 5123 23291
rect 5157 23257 5207 23291
rect 5425 23541 6127 23583
rect 5425 23507 5443 23541
rect 5477 23507 6075 23541
rect 6109 23507 6127 23541
rect 5425 23439 6127 23507
rect 6162 23541 7231 23583
rect 6162 23507 6179 23541
rect 6213 23507 7179 23541
rect 7213 23507 7231 23541
rect 6162 23496 7231 23507
rect 7265 23512 7323 23583
rect 5425 23405 5443 23439
rect 5477 23405 6075 23439
rect 6109 23405 6127 23439
rect 5425 23365 6127 23405
rect 5425 23295 5763 23365
rect 5425 23261 5503 23295
rect 5537 23261 5606 23295
rect 5640 23261 5709 23295
rect 5743 23261 5763 23295
rect 5797 23297 5817 23331
rect 5851 23297 5916 23331
rect 5950 23297 6015 23331
rect 6049 23297 6127 23331
rect 5797 23227 6127 23297
rect 6480 23295 6550 23496
rect 7265 23478 7277 23512
rect 7311 23478 7323 23512
rect 7265 23419 7323 23478
rect 7265 23385 7277 23419
rect 7311 23385 7323 23419
rect 7265 23350 7323 23385
rect 7449 23541 7967 23583
rect 7449 23507 7467 23541
rect 7501 23507 7915 23541
rect 7949 23507 7967 23541
rect 7449 23439 7967 23507
rect 8002 23541 9071 23583
rect 8002 23507 8019 23541
rect 8053 23507 9019 23541
rect 9053 23507 9071 23541
rect 8002 23496 9071 23507
rect 9106 23541 10175 23583
rect 9106 23507 9123 23541
rect 9157 23507 10123 23541
rect 10157 23507 10175 23541
rect 9106 23496 10175 23507
rect 10210 23541 11279 23583
rect 10210 23507 10227 23541
rect 10261 23507 11227 23541
rect 11261 23507 11279 23541
rect 10210 23496 11279 23507
rect 11314 23541 12383 23583
rect 11314 23507 11331 23541
rect 11365 23507 12331 23541
rect 12365 23507 12383 23541
rect 11314 23496 12383 23507
rect 12417 23512 12475 23583
rect 7449 23405 7467 23439
rect 7501 23405 7915 23439
rect 7949 23405 7967 23439
rect 7449 23365 7967 23405
rect 6480 23261 6499 23295
rect 6533 23261 6550 23295
rect 6480 23246 6550 23261
rect 6846 23331 6914 23348
rect 6846 23297 6863 23331
rect 6897 23297 6914 23331
rect 4965 23170 5207 23223
rect 4965 23136 4983 23170
rect 5017 23136 5155 23170
rect 5189 23136 5207 23170
rect 4965 23073 5207 23136
rect 5425 23168 6127 23227
rect 6846 23182 6914 23297
rect 7449 23295 7691 23365
rect 7449 23261 7527 23295
rect 7561 23261 7637 23295
rect 7671 23261 7691 23295
rect 7725 23297 7745 23331
rect 7779 23297 7855 23331
rect 7889 23297 7967 23331
rect 7725 23227 7967 23297
rect 8320 23295 8390 23496
rect 8320 23261 8339 23295
rect 8373 23261 8390 23295
rect 8320 23246 8390 23261
rect 8686 23331 8754 23348
rect 8686 23297 8703 23331
rect 8737 23297 8754 23331
rect 7265 23201 7323 23218
rect 5425 23134 5443 23168
rect 5477 23134 6075 23168
rect 6109 23134 6127 23168
rect 5425 23073 6127 23134
rect 6162 23168 7231 23182
rect 6162 23134 6179 23168
rect 6213 23134 7179 23168
rect 7213 23134 7231 23168
rect 6162 23073 7231 23134
rect 7265 23167 7277 23201
rect 7311 23167 7323 23201
rect 7265 23073 7323 23167
rect 7449 23168 7967 23227
rect 8686 23182 8754 23297
rect 9424 23295 9494 23496
rect 9424 23261 9443 23295
rect 9477 23261 9494 23295
rect 9424 23246 9494 23261
rect 9790 23331 9858 23348
rect 9790 23297 9807 23331
rect 9841 23297 9858 23331
rect 9790 23182 9858 23297
rect 10528 23295 10598 23496
rect 10528 23261 10547 23295
rect 10581 23261 10598 23295
rect 10528 23246 10598 23261
rect 10894 23331 10962 23348
rect 10894 23297 10911 23331
rect 10945 23297 10962 23331
rect 10894 23182 10962 23297
rect 11632 23295 11702 23496
rect 12417 23478 12429 23512
rect 12463 23478 12475 23512
rect 12417 23419 12475 23478
rect 12417 23385 12429 23419
rect 12463 23385 12475 23419
rect 12417 23350 12475 23385
rect 12601 23541 13119 23583
rect 12601 23507 12619 23541
rect 12653 23507 13067 23541
rect 13101 23507 13119 23541
rect 12601 23439 13119 23507
rect 13154 23541 14223 23583
rect 13154 23507 13171 23541
rect 13205 23507 14171 23541
rect 14205 23507 14223 23541
rect 13154 23496 14223 23507
rect 14258 23541 15327 23583
rect 14258 23507 14275 23541
rect 14309 23507 15275 23541
rect 15309 23507 15327 23541
rect 14258 23496 15327 23507
rect 15362 23541 16431 23583
rect 15362 23507 15379 23541
rect 15413 23507 16379 23541
rect 16413 23507 16431 23541
rect 15362 23496 16431 23507
rect 16466 23541 17535 23583
rect 16466 23507 16483 23541
rect 16517 23507 17483 23541
rect 17517 23507 17535 23541
rect 16466 23496 17535 23507
rect 17569 23512 17627 23583
rect 12601 23405 12619 23439
rect 12653 23405 13067 23439
rect 13101 23405 13119 23439
rect 12601 23365 13119 23405
rect 11632 23261 11651 23295
rect 11685 23261 11702 23295
rect 11632 23246 11702 23261
rect 11998 23331 12066 23348
rect 11998 23297 12015 23331
rect 12049 23297 12066 23331
rect 11998 23182 12066 23297
rect 12601 23295 12843 23365
rect 12601 23261 12679 23295
rect 12713 23261 12789 23295
rect 12823 23261 12843 23295
rect 12877 23297 12897 23331
rect 12931 23297 13007 23331
rect 13041 23297 13119 23331
rect 12877 23227 13119 23297
rect 13472 23295 13542 23496
rect 13472 23261 13491 23295
rect 13525 23261 13542 23295
rect 13472 23246 13542 23261
rect 13838 23331 13906 23348
rect 13838 23297 13855 23331
rect 13889 23297 13906 23331
rect 12417 23201 12475 23218
rect 7449 23134 7467 23168
rect 7501 23134 7915 23168
rect 7949 23134 7967 23168
rect 7449 23073 7967 23134
rect 8002 23168 9071 23182
rect 8002 23134 8019 23168
rect 8053 23134 9019 23168
rect 9053 23134 9071 23168
rect 8002 23073 9071 23134
rect 9106 23168 10175 23182
rect 9106 23134 9123 23168
rect 9157 23134 10123 23168
rect 10157 23134 10175 23168
rect 9106 23073 10175 23134
rect 10210 23168 11279 23182
rect 10210 23134 10227 23168
rect 10261 23134 11227 23168
rect 11261 23134 11279 23168
rect 10210 23073 11279 23134
rect 11314 23168 12383 23182
rect 11314 23134 11331 23168
rect 11365 23134 12331 23168
rect 12365 23134 12383 23168
rect 11314 23073 12383 23134
rect 12417 23167 12429 23201
rect 12463 23167 12475 23201
rect 12417 23073 12475 23167
rect 12601 23168 13119 23227
rect 13838 23182 13906 23297
rect 14576 23295 14646 23496
rect 14576 23261 14595 23295
rect 14629 23261 14646 23295
rect 14576 23246 14646 23261
rect 14942 23331 15010 23348
rect 14942 23297 14959 23331
rect 14993 23297 15010 23331
rect 14942 23182 15010 23297
rect 15680 23295 15750 23496
rect 15680 23261 15699 23295
rect 15733 23261 15750 23295
rect 15680 23246 15750 23261
rect 16046 23331 16114 23348
rect 16046 23297 16063 23331
rect 16097 23297 16114 23331
rect 16046 23182 16114 23297
rect 16784 23295 16854 23496
rect 17569 23478 17581 23512
rect 17615 23478 17627 23512
rect 17754 23541 18823 23583
rect 17754 23507 17771 23541
rect 17805 23507 18771 23541
rect 18805 23507 18823 23541
rect 17754 23496 18823 23507
rect 18858 23541 19927 23583
rect 18858 23507 18875 23541
rect 18909 23507 19875 23541
rect 19909 23507 19927 23541
rect 18858 23496 19927 23507
rect 19961 23541 20203 23583
rect 19961 23507 19979 23541
rect 20013 23507 20151 23541
rect 20185 23507 20203 23541
rect 17569 23419 17627 23478
rect 17569 23385 17581 23419
rect 17615 23385 17627 23419
rect 17569 23350 17627 23385
rect 16784 23261 16803 23295
rect 16837 23261 16854 23295
rect 16784 23246 16854 23261
rect 17150 23331 17218 23348
rect 17150 23297 17167 23331
rect 17201 23297 17218 23331
rect 17150 23182 17218 23297
rect 18072 23295 18142 23496
rect 18072 23261 18091 23295
rect 18125 23261 18142 23295
rect 18072 23246 18142 23261
rect 18438 23331 18506 23348
rect 18438 23297 18455 23331
rect 18489 23297 18506 23331
rect 17569 23201 17627 23218
rect 12601 23134 12619 23168
rect 12653 23134 13067 23168
rect 13101 23134 13119 23168
rect 12601 23073 13119 23134
rect 13154 23168 14223 23182
rect 13154 23134 13171 23168
rect 13205 23134 14171 23168
rect 14205 23134 14223 23168
rect 13154 23073 14223 23134
rect 14258 23168 15327 23182
rect 14258 23134 14275 23168
rect 14309 23134 15275 23168
rect 15309 23134 15327 23168
rect 14258 23073 15327 23134
rect 15362 23168 16431 23182
rect 15362 23134 15379 23168
rect 15413 23134 16379 23168
rect 16413 23134 16431 23168
rect 15362 23073 16431 23134
rect 16466 23168 17535 23182
rect 16466 23134 16483 23168
rect 16517 23134 17483 23168
rect 17517 23134 17535 23168
rect 16466 23073 17535 23134
rect 17569 23167 17581 23201
rect 17615 23167 17627 23201
rect 18438 23182 18506 23297
rect 19176 23295 19246 23496
rect 19961 23446 20203 23507
rect 19961 23412 19979 23446
rect 20013 23412 20151 23446
rect 20185 23412 20203 23446
rect 19961 23365 20203 23412
rect 19176 23261 19195 23295
rect 19229 23261 19246 23295
rect 19176 23246 19246 23261
rect 19542 23331 19610 23348
rect 19542 23297 19559 23331
rect 19593 23297 19610 23331
rect 19542 23182 19610 23297
rect 19961 23291 20065 23365
rect 19961 23257 20011 23291
rect 20045 23257 20065 23291
rect 20099 23297 20119 23331
rect 20153 23297 20203 23331
rect 20099 23223 20203 23297
rect 17569 23073 17627 23167
rect 17754 23168 18823 23182
rect 17754 23134 17771 23168
rect 17805 23134 18771 23168
rect 18805 23134 18823 23168
rect 17754 23073 18823 23134
rect 18858 23168 19927 23182
rect 18858 23134 18875 23168
rect 18909 23134 19875 23168
rect 19909 23134 19927 23168
rect 18858 23073 19927 23134
rect 19961 23170 20203 23223
rect 19961 23136 19979 23170
rect 20013 23136 20151 23170
rect 20185 23136 20203 23170
rect 19961 23073 20203 23136
rect 4948 23039 4977 23073
rect 5011 23039 5069 23073
rect 5103 23039 5161 23073
rect 5195 23039 5253 23073
rect 5287 23039 5345 23073
rect 5379 23039 5437 23073
rect 5471 23039 5529 23073
rect 5563 23039 5621 23073
rect 5655 23039 5713 23073
rect 5747 23039 5805 23073
rect 5839 23039 5897 23073
rect 5931 23039 5989 23073
rect 6023 23039 6081 23073
rect 6115 23039 6173 23073
rect 6207 23039 6265 23073
rect 6299 23039 6357 23073
rect 6391 23039 6449 23073
rect 6483 23039 6541 23073
rect 6575 23039 6633 23073
rect 6667 23039 6725 23073
rect 6759 23039 6817 23073
rect 6851 23039 6909 23073
rect 6943 23039 7001 23073
rect 7035 23039 7093 23073
rect 7127 23039 7185 23073
rect 7219 23039 7277 23073
rect 7311 23039 7369 23073
rect 7403 23039 7461 23073
rect 7495 23039 7553 23073
rect 7587 23039 7645 23073
rect 7679 23039 7737 23073
rect 7771 23039 7829 23073
rect 7863 23039 7921 23073
rect 7955 23039 8013 23073
rect 8047 23039 8105 23073
rect 8139 23039 8197 23073
rect 8231 23039 8289 23073
rect 8323 23039 8381 23073
rect 8415 23039 8473 23073
rect 8507 23039 8565 23073
rect 8599 23039 8657 23073
rect 8691 23039 8749 23073
rect 8783 23039 8841 23073
rect 8875 23039 8933 23073
rect 8967 23039 9025 23073
rect 9059 23039 9117 23073
rect 9151 23039 9209 23073
rect 9243 23039 9301 23073
rect 9335 23039 9393 23073
rect 9427 23039 9485 23073
rect 9519 23039 9577 23073
rect 9611 23039 9669 23073
rect 9703 23039 9761 23073
rect 9795 23039 9853 23073
rect 9887 23039 9945 23073
rect 9979 23039 10037 23073
rect 10071 23039 10129 23073
rect 10163 23039 10221 23073
rect 10255 23039 10313 23073
rect 10347 23039 10405 23073
rect 10439 23039 10497 23073
rect 10531 23039 10589 23073
rect 10623 23039 10681 23073
rect 10715 23039 10773 23073
rect 10807 23039 10865 23073
rect 10899 23039 10957 23073
rect 10991 23039 11049 23073
rect 11083 23039 11141 23073
rect 11175 23039 11233 23073
rect 11267 23039 11325 23073
rect 11359 23039 11417 23073
rect 11451 23039 11509 23073
rect 11543 23039 11601 23073
rect 11635 23039 11693 23073
rect 11727 23039 11785 23073
rect 11819 23039 11877 23073
rect 11911 23039 11969 23073
rect 12003 23039 12061 23073
rect 12095 23039 12153 23073
rect 12187 23039 12245 23073
rect 12279 23039 12337 23073
rect 12371 23039 12429 23073
rect 12463 23039 12521 23073
rect 12555 23039 12613 23073
rect 12647 23039 12705 23073
rect 12739 23039 12797 23073
rect 12831 23039 12889 23073
rect 12923 23039 12981 23073
rect 13015 23039 13073 23073
rect 13107 23039 13165 23073
rect 13199 23039 13257 23073
rect 13291 23039 13349 23073
rect 13383 23039 13441 23073
rect 13475 23039 13533 23073
rect 13567 23039 13625 23073
rect 13659 23039 13717 23073
rect 13751 23039 13809 23073
rect 13843 23039 13901 23073
rect 13935 23039 13993 23073
rect 14027 23039 14085 23073
rect 14119 23039 14177 23073
rect 14211 23039 14269 23073
rect 14303 23039 14361 23073
rect 14395 23039 14453 23073
rect 14487 23039 14545 23073
rect 14579 23039 14637 23073
rect 14671 23039 14729 23073
rect 14763 23039 14821 23073
rect 14855 23039 14913 23073
rect 14947 23039 15005 23073
rect 15039 23039 15097 23073
rect 15131 23039 15189 23073
rect 15223 23039 15281 23073
rect 15315 23039 15373 23073
rect 15407 23039 15465 23073
rect 15499 23039 15557 23073
rect 15591 23039 15649 23073
rect 15683 23039 15741 23073
rect 15775 23039 15833 23073
rect 15867 23039 15925 23073
rect 15959 23039 16017 23073
rect 16051 23039 16109 23073
rect 16143 23039 16201 23073
rect 16235 23039 16293 23073
rect 16327 23039 16385 23073
rect 16419 23039 16477 23073
rect 16511 23039 16569 23073
rect 16603 23039 16661 23073
rect 16695 23039 16753 23073
rect 16787 23039 16845 23073
rect 16879 23039 16937 23073
rect 16971 23039 17029 23073
rect 17063 23039 17121 23073
rect 17155 23039 17213 23073
rect 17247 23039 17305 23073
rect 17339 23039 17397 23073
rect 17431 23039 17489 23073
rect 17523 23039 17581 23073
rect 17615 23039 17673 23073
rect 17707 23039 17765 23073
rect 17799 23039 17857 23073
rect 17891 23039 17949 23073
rect 17983 23039 18041 23073
rect 18075 23039 18133 23073
rect 18167 23039 18225 23073
rect 18259 23039 18317 23073
rect 18351 23039 18409 23073
rect 18443 23039 18501 23073
rect 18535 23039 18593 23073
rect 18627 23039 18685 23073
rect 18719 23039 18777 23073
rect 18811 23039 18869 23073
rect 18903 23039 18961 23073
rect 18995 23039 19053 23073
rect 19087 23039 19145 23073
rect 19179 23039 19237 23073
rect 19271 23039 19329 23073
rect 19363 23039 19421 23073
rect 19455 23039 19513 23073
rect 19547 23039 19605 23073
rect 19639 23039 19697 23073
rect 19731 23039 19789 23073
rect 19823 23039 19881 23073
rect 19915 23039 19973 23073
rect 20007 23039 20065 23073
rect 20099 23039 20157 23073
rect 20191 23039 20220 23073
rect 4965 22976 5207 23039
rect 4965 22942 4983 22976
rect 5017 22942 5155 22976
rect 5189 22942 5207 22976
rect 4965 22889 5207 22942
rect 5426 22978 6495 23039
rect 5426 22944 5443 22978
rect 5477 22944 6443 22978
rect 6477 22944 6495 22978
rect 5426 22930 6495 22944
rect 6530 22978 7599 23039
rect 6530 22944 6547 22978
rect 6581 22944 7547 22978
rect 7581 22944 7599 22978
rect 6530 22930 7599 22944
rect 7634 22978 8703 23039
rect 7634 22944 7651 22978
rect 7685 22944 8651 22978
rect 8685 22944 8703 22978
rect 7634 22930 8703 22944
rect 8738 22978 9807 23039
rect 8738 22944 8755 22978
rect 8789 22944 9755 22978
rect 9789 22944 9807 22978
rect 8738 22930 9807 22944
rect 9841 22945 9899 23039
rect 4965 22815 5069 22889
rect 4965 22781 5015 22815
rect 5049 22781 5069 22815
rect 5103 22821 5123 22855
rect 5157 22821 5207 22855
rect 5103 22747 5207 22821
rect 4965 22700 5207 22747
rect 4965 22666 4983 22700
rect 5017 22666 5155 22700
rect 5189 22666 5207 22700
rect 4965 22605 5207 22666
rect 5744 22851 5814 22866
rect 5744 22817 5763 22851
rect 5797 22817 5814 22851
rect 5744 22616 5814 22817
rect 6110 22815 6178 22930
rect 6110 22781 6127 22815
rect 6161 22781 6178 22815
rect 6110 22764 6178 22781
rect 6848 22851 6918 22866
rect 6848 22817 6867 22851
rect 6901 22817 6918 22851
rect 6848 22616 6918 22817
rect 7214 22815 7282 22930
rect 7214 22781 7231 22815
rect 7265 22781 7282 22815
rect 7214 22764 7282 22781
rect 7952 22851 8022 22866
rect 7952 22817 7971 22851
rect 8005 22817 8022 22851
rect 7952 22616 8022 22817
rect 8318 22815 8386 22930
rect 8318 22781 8335 22815
rect 8369 22781 8386 22815
rect 8318 22764 8386 22781
rect 9056 22851 9126 22866
rect 9056 22817 9075 22851
rect 9109 22817 9126 22851
rect 9056 22616 9126 22817
rect 9422 22815 9490 22930
rect 9841 22911 9853 22945
rect 9887 22911 9899 22945
rect 9841 22894 9899 22911
rect 10025 22978 10543 23039
rect 10025 22944 10043 22978
rect 10077 22944 10491 22978
rect 10525 22944 10543 22978
rect 10025 22885 10543 22944
rect 10578 22978 11647 23039
rect 10578 22944 10595 22978
rect 10629 22944 11595 22978
rect 11629 22944 11647 22978
rect 10578 22930 11647 22944
rect 11682 22978 12751 23039
rect 11682 22944 11699 22978
rect 11733 22944 12699 22978
rect 12733 22944 12751 22978
rect 11682 22930 12751 22944
rect 12786 22978 13855 23039
rect 12786 22944 12803 22978
rect 12837 22944 13803 22978
rect 13837 22944 13855 22978
rect 12786 22930 13855 22944
rect 13890 22978 14959 23039
rect 13890 22944 13907 22978
rect 13941 22944 14907 22978
rect 14941 22944 14959 22978
rect 13890 22930 14959 22944
rect 14993 22945 15051 23039
rect 9422 22781 9439 22815
rect 9473 22781 9490 22815
rect 9422 22764 9490 22781
rect 10025 22817 10103 22851
rect 10137 22817 10213 22851
rect 10247 22817 10267 22851
rect 9841 22727 9899 22762
rect 9841 22693 9853 22727
rect 9887 22693 9899 22727
rect 9841 22634 9899 22693
rect 4965 22571 4983 22605
rect 5017 22571 5155 22605
rect 5189 22571 5207 22605
rect 4965 22529 5207 22571
rect 5426 22605 6495 22616
rect 5426 22571 5443 22605
rect 5477 22571 6443 22605
rect 6477 22571 6495 22605
rect 5426 22529 6495 22571
rect 6530 22605 7599 22616
rect 6530 22571 6547 22605
rect 6581 22571 7547 22605
rect 7581 22571 7599 22605
rect 6530 22529 7599 22571
rect 7634 22605 8703 22616
rect 7634 22571 7651 22605
rect 7685 22571 8651 22605
rect 8685 22571 8703 22605
rect 7634 22529 8703 22571
rect 8738 22605 9807 22616
rect 8738 22571 8755 22605
rect 8789 22571 9755 22605
rect 9789 22571 9807 22605
rect 8738 22529 9807 22571
rect 9841 22600 9853 22634
rect 9887 22600 9899 22634
rect 9841 22529 9899 22600
rect 10025 22747 10267 22817
rect 10301 22815 10543 22885
rect 10301 22781 10321 22815
rect 10355 22781 10431 22815
rect 10465 22781 10543 22815
rect 10896 22851 10966 22866
rect 10896 22817 10915 22851
rect 10949 22817 10966 22851
rect 10025 22707 10543 22747
rect 10025 22673 10043 22707
rect 10077 22673 10491 22707
rect 10525 22673 10543 22707
rect 10025 22605 10543 22673
rect 10896 22616 10966 22817
rect 11262 22815 11330 22930
rect 11262 22781 11279 22815
rect 11313 22781 11330 22815
rect 11262 22764 11330 22781
rect 12000 22851 12070 22866
rect 12000 22817 12019 22851
rect 12053 22817 12070 22851
rect 12000 22616 12070 22817
rect 12366 22815 12434 22930
rect 12366 22781 12383 22815
rect 12417 22781 12434 22815
rect 12366 22764 12434 22781
rect 13104 22851 13174 22866
rect 13104 22817 13123 22851
rect 13157 22817 13174 22851
rect 13104 22616 13174 22817
rect 13470 22815 13538 22930
rect 13470 22781 13487 22815
rect 13521 22781 13538 22815
rect 13470 22764 13538 22781
rect 14208 22851 14278 22866
rect 14208 22817 14227 22851
rect 14261 22817 14278 22851
rect 14208 22616 14278 22817
rect 14574 22815 14642 22930
rect 14993 22911 15005 22945
rect 15039 22911 15051 22945
rect 14993 22894 15051 22911
rect 15177 22971 15511 23039
rect 15177 22937 15195 22971
rect 15229 22937 15459 22971
rect 15493 22937 15511 22971
rect 15177 22885 15511 22937
rect 15546 22978 16615 23039
rect 15546 22944 15563 22978
rect 15597 22944 16563 22978
rect 16597 22944 16615 22978
rect 15546 22930 16615 22944
rect 16650 22978 17719 23039
rect 16650 22944 16667 22978
rect 16701 22944 17667 22978
rect 17701 22944 17719 22978
rect 16650 22930 17719 22944
rect 17754 22978 18823 23039
rect 17754 22944 17771 22978
rect 17805 22944 18771 22978
rect 18805 22944 18823 22978
rect 17754 22930 18823 22944
rect 18858 22978 19927 23039
rect 18858 22944 18875 22978
rect 18909 22944 19875 22978
rect 19909 22944 19927 22978
rect 18858 22930 19927 22944
rect 19961 22976 20203 23039
rect 19961 22942 19979 22976
rect 20013 22942 20151 22976
rect 20185 22942 20203 22976
rect 14574 22781 14591 22815
rect 14625 22781 14642 22815
rect 14574 22764 14642 22781
rect 15177 22817 15197 22851
rect 15231 22817 15327 22851
rect 14993 22727 15051 22762
rect 14993 22693 15005 22727
rect 15039 22693 15051 22727
rect 14993 22634 15051 22693
rect 10025 22571 10043 22605
rect 10077 22571 10491 22605
rect 10525 22571 10543 22605
rect 10025 22529 10543 22571
rect 10578 22605 11647 22616
rect 10578 22571 10595 22605
rect 10629 22571 11595 22605
rect 11629 22571 11647 22605
rect 10578 22529 11647 22571
rect 11682 22605 12751 22616
rect 11682 22571 11699 22605
rect 11733 22571 12699 22605
rect 12733 22571 12751 22605
rect 11682 22529 12751 22571
rect 12786 22605 13855 22616
rect 12786 22571 12803 22605
rect 12837 22571 13803 22605
rect 13837 22571 13855 22605
rect 12786 22529 13855 22571
rect 13890 22605 14959 22616
rect 13890 22571 13907 22605
rect 13941 22571 14907 22605
rect 14941 22571 14959 22605
rect 13890 22529 14959 22571
rect 14993 22600 15005 22634
rect 15039 22600 15051 22634
rect 14993 22529 15051 22600
rect 15177 22747 15327 22817
rect 15361 22815 15511 22885
rect 15361 22781 15457 22815
rect 15491 22781 15511 22815
rect 15864 22851 15934 22866
rect 15864 22817 15883 22851
rect 15917 22817 15934 22851
rect 15177 22707 15511 22747
rect 15177 22673 15195 22707
rect 15229 22673 15459 22707
rect 15493 22673 15511 22707
rect 15177 22605 15511 22673
rect 15864 22616 15934 22817
rect 16230 22815 16298 22930
rect 16230 22781 16247 22815
rect 16281 22781 16298 22815
rect 16230 22764 16298 22781
rect 16968 22851 17038 22866
rect 16968 22817 16987 22851
rect 17021 22817 17038 22851
rect 16968 22616 17038 22817
rect 17334 22815 17402 22930
rect 17334 22781 17351 22815
rect 17385 22781 17402 22815
rect 17334 22764 17402 22781
rect 18072 22851 18142 22866
rect 18072 22817 18091 22851
rect 18125 22817 18142 22851
rect 18072 22616 18142 22817
rect 18438 22815 18506 22930
rect 18438 22781 18455 22815
rect 18489 22781 18506 22815
rect 18438 22764 18506 22781
rect 19176 22851 19246 22866
rect 19176 22817 19195 22851
rect 19229 22817 19246 22851
rect 19176 22616 19246 22817
rect 19542 22815 19610 22930
rect 19961 22889 20203 22942
rect 19542 22781 19559 22815
rect 19593 22781 19610 22815
rect 19542 22764 19610 22781
rect 19961 22821 20011 22855
rect 20045 22821 20065 22855
rect 19961 22747 20065 22821
rect 20099 22815 20203 22889
rect 20099 22781 20119 22815
rect 20153 22781 20203 22815
rect 19961 22700 20203 22747
rect 19961 22666 19979 22700
rect 20013 22666 20151 22700
rect 20185 22666 20203 22700
rect 15177 22571 15195 22605
rect 15229 22571 15459 22605
rect 15493 22571 15511 22605
rect 15177 22529 15511 22571
rect 15546 22605 16615 22616
rect 15546 22571 15563 22605
rect 15597 22571 16563 22605
rect 16597 22571 16615 22605
rect 15546 22529 16615 22571
rect 16650 22605 17719 22616
rect 16650 22571 16667 22605
rect 16701 22571 17667 22605
rect 17701 22571 17719 22605
rect 16650 22529 17719 22571
rect 17754 22605 18823 22616
rect 17754 22571 17771 22605
rect 17805 22571 18771 22605
rect 18805 22571 18823 22605
rect 17754 22529 18823 22571
rect 18858 22605 19927 22616
rect 18858 22571 18875 22605
rect 18909 22571 19875 22605
rect 19909 22571 19927 22605
rect 18858 22529 19927 22571
rect 19961 22605 20203 22666
rect 19961 22571 19979 22605
rect 20013 22571 20151 22605
rect 20185 22571 20203 22605
rect 19961 22529 20203 22571
rect 4948 22495 4977 22529
rect 5011 22495 5069 22529
rect 5103 22495 5161 22529
rect 5195 22495 5253 22529
rect 5287 22495 5345 22529
rect 5379 22495 5437 22529
rect 5471 22495 5529 22529
rect 5563 22495 5621 22529
rect 5655 22495 5713 22529
rect 5747 22495 5805 22529
rect 5839 22495 5897 22529
rect 5931 22495 5989 22529
rect 6023 22495 6081 22529
rect 6115 22495 6173 22529
rect 6207 22495 6265 22529
rect 6299 22495 6357 22529
rect 6391 22495 6449 22529
rect 6483 22495 6541 22529
rect 6575 22495 6633 22529
rect 6667 22495 6725 22529
rect 6759 22495 6817 22529
rect 6851 22495 6909 22529
rect 6943 22495 7001 22529
rect 7035 22495 7093 22529
rect 7127 22495 7185 22529
rect 7219 22495 7277 22529
rect 7311 22495 7369 22529
rect 7403 22495 7461 22529
rect 7495 22495 7553 22529
rect 7587 22495 7645 22529
rect 7679 22495 7737 22529
rect 7771 22495 7829 22529
rect 7863 22495 7921 22529
rect 7955 22495 8013 22529
rect 8047 22495 8105 22529
rect 8139 22495 8197 22529
rect 8231 22495 8289 22529
rect 8323 22495 8381 22529
rect 8415 22495 8473 22529
rect 8507 22495 8565 22529
rect 8599 22495 8657 22529
rect 8691 22495 8749 22529
rect 8783 22495 8841 22529
rect 8875 22495 8933 22529
rect 8967 22495 9025 22529
rect 9059 22495 9117 22529
rect 9151 22495 9209 22529
rect 9243 22495 9301 22529
rect 9335 22495 9393 22529
rect 9427 22495 9485 22529
rect 9519 22495 9577 22529
rect 9611 22495 9669 22529
rect 9703 22495 9761 22529
rect 9795 22495 9853 22529
rect 9887 22495 9945 22529
rect 9979 22495 10037 22529
rect 10071 22495 10129 22529
rect 10163 22495 10221 22529
rect 10255 22495 10313 22529
rect 10347 22495 10405 22529
rect 10439 22495 10497 22529
rect 10531 22495 10589 22529
rect 10623 22495 10681 22529
rect 10715 22495 10773 22529
rect 10807 22495 10865 22529
rect 10899 22495 10957 22529
rect 10991 22495 11049 22529
rect 11083 22495 11141 22529
rect 11175 22495 11233 22529
rect 11267 22495 11325 22529
rect 11359 22495 11417 22529
rect 11451 22495 11509 22529
rect 11543 22495 11601 22529
rect 11635 22495 11693 22529
rect 11727 22495 11785 22529
rect 11819 22495 11877 22529
rect 11911 22495 11969 22529
rect 12003 22495 12061 22529
rect 12095 22495 12153 22529
rect 12187 22495 12245 22529
rect 12279 22495 12337 22529
rect 12371 22495 12429 22529
rect 12463 22495 12521 22529
rect 12555 22495 12613 22529
rect 12647 22495 12705 22529
rect 12739 22495 12797 22529
rect 12831 22495 12889 22529
rect 12923 22495 12981 22529
rect 13015 22495 13073 22529
rect 13107 22495 13165 22529
rect 13199 22495 13257 22529
rect 13291 22495 13349 22529
rect 13383 22495 13441 22529
rect 13475 22495 13533 22529
rect 13567 22495 13625 22529
rect 13659 22495 13717 22529
rect 13751 22495 13809 22529
rect 13843 22495 13901 22529
rect 13935 22495 13993 22529
rect 14027 22495 14085 22529
rect 14119 22495 14177 22529
rect 14211 22495 14269 22529
rect 14303 22495 14361 22529
rect 14395 22495 14453 22529
rect 14487 22495 14545 22529
rect 14579 22495 14637 22529
rect 14671 22495 14729 22529
rect 14763 22495 14821 22529
rect 14855 22495 14913 22529
rect 14947 22495 15005 22529
rect 15039 22495 15097 22529
rect 15131 22495 15189 22529
rect 15223 22495 15281 22529
rect 15315 22495 15373 22529
rect 15407 22495 15465 22529
rect 15499 22495 15557 22529
rect 15591 22495 15649 22529
rect 15683 22495 15741 22529
rect 15775 22495 15833 22529
rect 15867 22495 15925 22529
rect 15959 22495 16017 22529
rect 16051 22495 16109 22529
rect 16143 22495 16201 22529
rect 16235 22495 16293 22529
rect 16327 22495 16385 22529
rect 16419 22495 16477 22529
rect 16511 22495 16569 22529
rect 16603 22495 16661 22529
rect 16695 22495 16753 22529
rect 16787 22495 16845 22529
rect 16879 22495 16937 22529
rect 16971 22495 17029 22529
rect 17063 22495 17121 22529
rect 17155 22495 17213 22529
rect 17247 22495 17305 22529
rect 17339 22495 17397 22529
rect 17431 22495 17489 22529
rect 17523 22495 17581 22529
rect 17615 22495 17673 22529
rect 17707 22495 17765 22529
rect 17799 22495 17857 22529
rect 17891 22495 17949 22529
rect 17983 22495 18041 22529
rect 18075 22495 18133 22529
rect 18167 22495 18225 22529
rect 18259 22495 18317 22529
rect 18351 22495 18409 22529
rect 18443 22495 18501 22529
rect 18535 22495 18593 22529
rect 18627 22495 18685 22529
rect 18719 22495 18777 22529
rect 18811 22495 18869 22529
rect 18903 22495 18961 22529
rect 18995 22495 19053 22529
rect 19087 22495 19145 22529
rect 19179 22495 19237 22529
rect 19271 22495 19329 22529
rect 19363 22495 19421 22529
rect 19455 22495 19513 22529
rect 19547 22495 19605 22529
rect 19639 22495 19697 22529
rect 19731 22495 19789 22529
rect 19823 22495 19881 22529
rect 19915 22495 19973 22529
rect 20007 22495 20065 22529
rect 20099 22495 20157 22529
rect 20191 22495 20220 22529
rect 4965 22453 5207 22495
rect 4965 22419 4983 22453
rect 5017 22419 5155 22453
rect 5189 22419 5207 22453
rect 4965 22358 5207 22419
rect 4965 22324 4983 22358
rect 5017 22324 5155 22358
rect 5189 22324 5207 22358
rect 4965 22277 5207 22324
rect 4965 22209 5015 22243
rect 5049 22209 5069 22243
rect 4965 22135 5069 22209
rect 5103 22203 5207 22277
rect 5103 22169 5123 22203
rect 5157 22169 5207 22203
rect 5425 22453 6127 22495
rect 5425 22419 5443 22453
rect 5477 22419 6075 22453
rect 6109 22419 6127 22453
rect 5425 22351 6127 22419
rect 6162 22453 7231 22495
rect 6162 22419 6179 22453
rect 6213 22419 7179 22453
rect 7213 22419 7231 22453
rect 6162 22408 7231 22419
rect 7265 22424 7323 22495
rect 5425 22317 5443 22351
rect 5477 22317 6075 22351
rect 6109 22317 6127 22351
rect 5425 22277 6127 22317
rect 5425 22207 5763 22277
rect 5425 22173 5503 22207
rect 5537 22173 5606 22207
rect 5640 22173 5709 22207
rect 5743 22173 5763 22207
rect 5797 22209 5817 22243
rect 5851 22209 5916 22243
rect 5950 22209 6015 22243
rect 6049 22209 6127 22243
rect 5797 22139 6127 22209
rect 6480 22207 6550 22408
rect 7265 22390 7277 22424
rect 7311 22390 7323 22424
rect 7265 22331 7323 22390
rect 7265 22297 7277 22331
rect 7311 22297 7323 22331
rect 7265 22262 7323 22297
rect 7449 22453 7967 22495
rect 7449 22419 7467 22453
rect 7501 22419 7915 22453
rect 7949 22419 7967 22453
rect 7449 22351 7967 22419
rect 8002 22453 9071 22495
rect 8002 22419 8019 22453
rect 8053 22419 9019 22453
rect 9053 22419 9071 22453
rect 8002 22408 9071 22419
rect 9106 22453 10175 22495
rect 9106 22419 9123 22453
rect 9157 22419 10123 22453
rect 10157 22419 10175 22453
rect 9106 22408 10175 22419
rect 10210 22453 11279 22495
rect 10210 22419 10227 22453
rect 10261 22419 11227 22453
rect 11261 22419 11279 22453
rect 10210 22408 11279 22419
rect 11314 22453 12383 22495
rect 11314 22419 11331 22453
rect 11365 22419 12331 22453
rect 12365 22419 12383 22453
rect 11314 22408 12383 22419
rect 12417 22424 12475 22495
rect 7449 22317 7467 22351
rect 7501 22317 7915 22351
rect 7949 22317 7967 22351
rect 7449 22277 7967 22317
rect 6480 22173 6499 22207
rect 6533 22173 6550 22207
rect 6480 22158 6550 22173
rect 6846 22243 6914 22260
rect 6846 22209 6863 22243
rect 6897 22209 6914 22243
rect 4965 22082 5207 22135
rect 4965 22048 4983 22082
rect 5017 22048 5155 22082
rect 5189 22048 5207 22082
rect 4965 21985 5207 22048
rect 5425 22080 6127 22139
rect 6846 22094 6914 22209
rect 7449 22207 7691 22277
rect 7449 22173 7527 22207
rect 7561 22173 7637 22207
rect 7671 22173 7691 22207
rect 7725 22209 7745 22243
rect 7779 22209 7855 22243
rect 7889 22209 7967 22243
rect 7725 22139 7967 22209
rect 8320 22207 8390 22408
rect 8320 22173 8339 22207
rect 8373 22173 8390 22207
rect 8320 22158 8390 22173
rect 8686 22243 8754 22260
rect 8686 22209 8703 22243
rect 8737 22209 8754 22243
rect 7265 22113 7323 22130
rect 5425 22046 5443 22080
rect 5477 22046 6075 22080
rect 6109 22046 6127 22080
rect 5425 21985 6127 22046
rect 6162 22080 7231 22094
rect 6162 22046 6179 22080
rect 6213 22046 7179 22080
rect 7213 22046 7231 22080
rect 6162 21985 7231 22046
rect 7265 22079 7277 22113
rect 7311 22079 7323 22113
rect 7265 21985 7323 22079
rect 7449 22080 7967 22139
rect 8686 22094 8754 22209
rect 9424 22207 9494 22408
rect 9424 22173 9443 22207
rect 9477 22173 9494 22207
rect 9424 22158 9494 22173
rect 9790 22243 9858 22260
rect 9790 22209 9807 22243
rect 9841 22209 9858 22243
rect 9790 22094 9858 22209
rect 10528 22207 10598 22408
rect 10528 22173 10547 22207
rect 10581 22173 10598 22207
rect 10528 22158 10598 22173
rect 10894 22243 10962 22260
rect 10894 22209 10911 22243
rect 10945 22209 10962 22243
rect 10894 22094 10962 22209
rect 11632 22207 11702 22408
rect 12417 22390 12429 22424
rect 12463 22390 12475 22424
rect 12417 22331 12475 22390
rect 12417 22297 12429 22331
rect 12463 22297 12475 22331
rect 12417 22262 12475 22297
rect 12601 22453 13119 22495
rect 12601 22419 12619 22453
rect 12653 22419 13067 22453
rect 13101 22419 13119 22453
rect 12601 22351 13119 22419
rect 13154 22453 14223 22495
rect 13154 22419 13171 22453
rect 13205 22419 14171 22453
rect 14205 22419 14223 22453
rect 13154 22408 14223 22419
rect 14258 22453 15327 22495
rect 14258 22419 14275 22453
rect 14309 22419 15275 22453
rect 15309 22419 15327 22453
rect 14258 22408 15327 22419
rect 15362 22453 16431 22495
rect 15362 22419 15379 22453
rect 15413 22419 16379 22453
rect 16413 22419 16431 22453
rect 15362 22408 16431 22419
rect 16466 22453 17535 22495
rect 16466 22419 16483 22453
rect 16517 22419 17483 22453
rect 17517 22419 17535 22453
rect 16466 22408 17535 22419
rect 17569 22424 17627 22495
rect 12601 22317 12619 22351
rect 12653 22317 13067 22351
rect 13101 22317 13119 22351
rect 12601 22277 13119 22317
rect 11632 22173 11651 22207
rect 11685 22173 11702 22207
rect 11632 22158 11702 22173
rect 11998 22243 12066 22260
rect 11998 22209 12015 22243
rect 12049 22209 12066 22243
rect 11998 22094 12066 22209
rect 12601 22207 12843 22277
rect 12601 22173 12679 22207
rect 12713 22173 12789 22207
rect 12823 22173 12843 22207
rect 12877 22209 12897 22243
rect 12931 22209 13007 22243
rect 13041 22209 13119 22243
rect 12877 22139 13119 22209
rect 13472 22207 13542 22408
rect 13472 22173 13491 22207
rect 13525 22173 13542 22207
rect 13472 22158 13542 22173
rect 13838 22243 13906 22260
rect 13838 22209 13855 22243
rect 13889 22209 13906 22243
rect 12417 22113 12475 22130
rect 7449 22046 7467 22080
rect 7501 22046 7915 22080
rect 7949 22046 7967 22080
rect 7449 21985 7967 22046
rect 8002 22080 9071 22094
rect 8002 22046 8019 22080
rect 8053 22046 9019 22080
rect 9053 22046 9071 22080
rect 8002 21985 9071 22046
rect 9106 22080 10175 22094
rect 9106 22046 9123 22080
rect 9157 22046 10123 22080
rect 10157 22046 10175 22080
rect 9106 21985 10175 22046
rect 10210 22080 11279 22094
rect 10210 22046 10227 22080
rect 10261 22046 11227 22080
rect 11261 22046 11279 22080
rect 10210 21985 11279 22046
rect 11314 22080 12383 22094
rect 11314 22046 11331 22080
rect 11365 22046 12331 22080
rect 12365 22046 12383 22080
rect 11314 21985 12383 22046
rect 12417 22079 12429 22113
rect 12463 22079 12475 22113
rect 12417 21985 12475 22079
rect 12601 22080 13119 22139
rect 13838 22094 13906 22209
rect 14576 22207 14646 22408
rect 14576 22173 14595 22207
rect 14629 22173 14646 22207
rect 14576 22158 14646 22173
rect 14942 22243 15010 22260
rect 14942 22209 14959 22243
rect 14993 22209 15010 22243
rect 14942 22094 15010 22209
rect 15680 22207 15750 22408
rect 15680 22173 15699 22207
rect 15733 22173 15750 22207
rect 15680 22158 15750 22173
rect 16046 22243 16114 22260
rect 16046 22209 16063 22243
rect 16097 22209 16114 22243
rect 16046 22094 16114 22209
rect 16784 22207 16854 22408
rect 17569 22390 17581 22424
rect 17615 22390 17627 22424
rect 17754 22453 18823 22495
rect 17754 22419 17771 22453
rect 17805 22419 18771 22453
rect 18805 22419 18823 22453
rect 17754 22408 18823 22419
rect 18858 22453 19927 22495
rect 18858 22419 18875 22453
rect 18909 22419 19875 22453
rect 19909 22419 19927 22453
rect 18858 22408 19927 22419
rect 19961 22453 20203 22495
rect 19961 22419 19979 22453
rect 20013 22419 20151 22453
rect 20185 22419 20203 22453
rect 17569 22331 17627 22390
rect 17569 22297 17581 22331
rect 17615 22297 17627 22331
rect 17569 22262 17627 22297
rect 16784 22173 16803 22207
rect 16837 22173 16854 22207
rect 16784 22158 16854 22173
rect 17150 22243 17218 22260
rect 17150 22209 17167 22243
rect 17201 22209 17218 22243
rect 17150 22094 17218 22209
rect 18072 22207 18142 22408
rect 18072 22173 18091 22207
rect 18125 22173 18142 22207
rect 18072 22158 18142 22173
rect 18438 22243 18506 22260
rect 18438 22209 18455 22243
rect 18489 22209 18506 22243
rect 17569 22113 17627 22130
rect 12601 22046 12619 22080
rect 12653 22046 13067 22080
rect 13101 22046 13119 22080
rect 12601 21985 13119 22046
rect 13154 22080 14223 22094
rect 13154 22046 13171 22080
rect 13205 22046 14171 22080
rect 14205 22046 14223 22080
rect 13154 21985 14223 22046
rect 14258 22080 15327 22094
rect 14258 22046 14275 22080
rect 14309 22046 15275 22080
rect 15309 22046 15327 22080
rect 14258 21985 15327 22046
rect 15362 22080 16431 22094
rect 15362 22046 15379 22080
rect 15413 22046 16379 22080
rect 16413 22046 16431 22080
rect 15362 21985 16431 22046
rect 16466 22080 17535 22094
rect 16466 22046 16483 22080
rect 16517 22046 17483 22080
rect 17517 22046 17535 22080
rect 16466 21985 17535 22046
rect 17569 22079 17581 22113
rect 17615 22079 17627 22113
rect 18438 22094 18506 22209
rect 19176 22207 19246 22408
rect 19961 22358 20203 22419
rect 19961 22324 19979 22358
rect 20013 22324 20151 22358
rect 20185 22324 20203 22358
rect 19961 22277 20203 22324
rect 19176 22173 19195 22207
rect 19229 22173 19246 22207
rect 19176 22158 19246 22173
rect 19542 22243 19610 22260
rect 19542 22209 19559 22243
rect 19593 22209 19610 22243
rect 19542 22094 19610 22209
rect 19961 22203 20065 22277
rect 19961 22169 20011 22203
rect 20045 22169 20065 22203
rect 20099 22209 20119 22243
rect 20153 22209 20203 22243
rect 20099 22135 20203 22209
rect 17569 21985 17627 22079
rect 17754 22080 18823 22094
rect 17754 22046 17771 22080
rect 17805 22046 18771 22080
rect 18805 22046 18823 22080
rect 17754 21985 18823 22046
rect 18858 22080 19927 22094
rect 18858 22046 18875 22080
rect 18909 22046 19875 22080
rect 19909 22046 19927 22080
rect 18858 21985 19927 22046
rect 19961 22082 20203 22135
rect 19961 22048 19979 22082
rect 20013 22048 20151 22082
rect 20185 22048 20203 22082
rect 19961 21985 20203 22048
rect 4948 21951 4977 21985
rect 5011 21951 5069 21985
rect 5103 21951 5161 21985
rect 5195 21951 5253 21985
rect 5287 21951 5345 21985
rect 5379 21951 5437 21985
rect 5471 21951 5529 21985
rect 5563 21951 5621 21985
rect 5655 21951 5713 21985
rect 5747 21951 5805 21985
rect 5839 21951 5897 21985
rect 5931 21951 5989 21985
rect 6023 21951 6081 21985
rect 6115 21951 6173 21985
rect 6207 21951 6265 21985
rect 6299 21951 6357 21985
rect 6391 21951 6449 21985
rect 6483 21951 6541 21985
rect 6575 21951 6633 21985
rect 6667 21951 6725 21985
rect 6759 21951 6817 21985
rect 6851 21951 6909 21985
rect 6943 21951 7001 21985
rect 7035 21951 7093 21985
rect 7127 21951 7185 21985
rect 7219 21951 7277 21985
rect 7311 21951 7369 21985
rect 7403 21951 7461 21985
rect 7495 21951 7553 21985
rect 7587 21951 7645 21985
rect 7679 21951 7737 21985
rect 7771 21951 7829 21985
rect 7863 21951 7921 21985
rect 7955 21951 8013 21985
rect 8047 21951 8105 21985
rect 8139 21951 8197 21985
rect 8231 21951 8289 21985
rect 8323 21951 8381 21985
rect 8415 21951 8473 21985
rect 8507 21951 8565 21985
rect 8599 21951 8657 21985
rect 8691 21951 8749 21985
rect 8783 21951 8841 21985
rect 8875 21951 8933 21985
rect 8967 21951 9025 21985
rect 9059 21951 9117 21985
rect 9151 21951 9209 21985
rect 9243 21951 9301 21985
rect 9335 21951 9393 21985
rect 9427 21951 9485 21985
rect 9519 21951 9577 21985
rect 9611 21951 9669 21985
rect 9703 21951 9761 21985
rect 9795 21951 9853 21985
rect 9887 21951 9945 21985
rect 9979 21951 10037 21985
rect 10071 21951 10129 21985
rect 10163 21951 10221 21985
rect 10255 21951 10313 21985
rect 10347 21951 10405 21985
rect 10439 21951 10497 21985
rect 10531 21951 10589 21985
rect 10623 21951 10681 21985
rect 10715 21951 10773 21985
rect 10807 21951 10865 21985
rect 10899 21951 10957 21985
rect 10991 21951 11049 21985
rect 11083 21951 11141 21985
rect 11175 21951 11233 21985
rect 11267 21951 11325 21985
rect 11359 21951 11417 21985
rect 11451 21951 11509 21985
rect 11543 21951 11601 21985
rect 11635 21951 11693 21985
rect 11727 21951 11785 21985
rect 11819 21951 11877 21985
rect 11911 21951 11969 21985
rect 12003 21951 12061 21985
rect 12095 21951 12153 21985
rect 12187 21951 12245 21985
rect 12279 21951 12337 21985
rect 12371 21951 12429 21985
rect 12463 21951 12521 21985
rect 12555 21951 12613 21985
rect 12647 21951 12705 21985
rect 12739 21951 12797 21985
rect 12831 21951 12889 21985
rect 12923 21951 12981 21985
rect 13015 21951 13073 21985
rect 13107 21951 13165 21985
rect 13199 21951 13257 21985
rect 13291 21951 13349 21985
rect 13383 21951 13441 21985
rect 13475 21951 13533 21985
rect 13567 21951 13625 21985
rect 13659 21951 13717 21985
rect 13751 21951 13809 21985
rect 13843 21951 13901 21985
rect 13935 21951 13993 21985
rect 14027 21951 14085 21985
rect 14119 21951 14177 21985
rect 14211 21951 14269 21985
rect 14303 21951 14361 21985
rect 14395 21951 14453 21985
rect 14487 21951 14545 21985
rect 14579 21951 14637 21985
rect 14671 21951 14729 21985
rect 14763 21951 14821 21985
rect 14855 21951 14913 21985
rect 14947 21951 15005 21985
rect 15039 21951 15097 21985
rect 15131 21951 15189 21985
rect 15223 21951 15281 21985
rect 15315 21951 15373 21985
rect 15407 21951 15465 21985
rect 15499 21951 15557 21985
rect 15591 21951 15649 21985
rect 15683 21951 15741 21985
rect 15775 21951 15833 21985
rect 15867 21951 15925 21985
rect 15959 21951 16017 21985
rect 16051 21951 16109 21985
rect 16143 21951 16201 21985
rect 16235 21951 16293 21985
rect 16327 21951 16385 21985
rect 16419 21951 16477 21985
rect 16511 21951 16569 21985
rect 16603 21951 16661 21985
rect 16695 21951 16753 21985
rect 16787 21951 16845 21985
rect 16879 21951 16937 21985
rect 16971 21951 17029 21985
rect 17063 21951 17121 21985
rect 17155 21951 17213 21985
rect 17247 21951 17305 21985
rect 17339 21951 17397 21985
rect 17431 21951 17489 21985
rect 17523 21951 17581 21985
rect 17615 21951 17673 21985
rect 17707 21951 17765 21985
rect 17799 21951 17857 21985
rect 17891 21951 17949 21985
rect 17983 21951 18041 21985
rect 18075 21951 18133 21985
rect 18167 21951 18225 21985
rect 18259 21951 18317 21985
rect 18351 21951 18409 21985
rect 18443 21951 18501 21985
rect 18535 21951 18593 21985
rect 18627 21951 18685 21985
rect 18719 21951 18777 21985
rect 18811 21951 18869 21985
rect 18903 21951 18961 21985
rect 18995 21951 19053 21985
rect 19087 21951 19145 21985
rect 19179 21951 19237 21985
rect 19271 21951 19329 21985
rect 19363 21951 19421 21985
rect 19455 21951 19513 21985
rect 19547 21951 19605 21985
rect 19639 21951 19697 21985
rect 19731 21951 19789 21985
rect 19823 21951 19881 21985
rect 19915 21951 19973 21985
rect 20007 21951 20065 21985
rect 20099 21951 20157 21985
rect 20191 21951 20220 21985
rect 4965 21888 5207 21951
rect 4965 21854 4983 21888
rect 5017 21854 5155 21888
rect 5189 21854 5207 21888
rect 4965 21801 5207 21854
rect 5426 21890 6495 21951
rect 5426 21856 5443 21890
rect 5477 21856 6443 21890
rect 6477 21856 6495 21890
rect 5426 21842 6495 21856
rect 6530 21890 7599 21951
rect 6530 21856 6547 21890
rect 6581 21856 7547 21890
rect 7581 21856 7599 21890
rect 6530 21842 7599 21856
rect 7634 21890 8703 21951
rect 7634 21856 7651 21890
rect 7685 21856 8651 21890
rect 8685 21856 8703 21890
rect 7634 21842 8703 21856
rect 8738 21890 9807 21951
rect 8738 21856 8755 21890
rect 8789 21856 9755 21890
rect 9789 21856 9807 21890
rect 8738 21842 9807 21856
rect 9841 21857 9899 21951
rect 4965 21727 5069 21801
rect 4965 21693 5015 21727
rect 5049 21693 5069 21727
rect 5103 21733 5123 21767
rect 5157 21733 5207 21767
rect 5103 21659 5207 21733
rect 4965 21612 5207 21659
rect 4965 21578 4983 21612
rect 5017 21578 5155 21612
rect 5189 21578 5207 21612
rect 4965 21517 5207 21578
rect 5744 21763 5814 21778
rect 5744 21729 5763 21763
rect 5797 21729 5814 21763
rect 5744 21528 5814 21729
rect 6110 21727 6178 21842
rect 6110 21693 6127 21727
rect 6161 21693 6178 21727
rect 6110 21676 6178 21693
rect 6848 21763 6918 21778
rect 6848 21729 6867 21763
rect 6901 21729 6918 21763
rect 6848 21528 6918 21729
rect 7214 21727 7282 21842
rect 7214 21693 7231 21727
rect 7265 21693 7282 21727
rect 7214 21676 7282 21693
rect 7952 21763 8022 21778
rect 7952 21729 7971 21763
rect 8005 21729 8022 21763
rect 7952 21528 8022 21729
rect 8318 21727 8386 21842
rect 8318 21693 8335 21727
rect 8369 21693 8386 21727
rect 8318 21676 8386 21693
rect 9056 21763 9126 21778
rect 9056 21729 9075 21763
rect 9109 21729 9126 21763
rect 9056 21528 9126 21729
rect 9422 21727 9490 21842
rect 9841 21823 9853 21857
rect 9887 21823 9899 21857
rect 9841 21806 9899 21823
rect 10025 21890 10543 21951
rect 10025 21856 10043 21890
rect 10077 21856 10491 21890
rect 10525 21856 10543 21890
rect 10025 21797 10543 21856
rect 10578 21890 11647 21951
rect 10578 21856 10595 21890
rect 10629 21856 11595 21890
rect 11629 21856 11647 21890
rect 10578 21842 11647 21856
rect 11682 21890 12751 21951
rect 11682 21856 11699 21890
rect 11733 21856 12699 21890
rect 12733 21856 12751 21890
rect 11682 21842 12751 21856
rect 12786 21890 13855 21951
rect 12786 21856 12803 21890
rect 12837 21856 13803 21890
rect 13837 21856 13855 21890
rect 12786 21842 13855 21856
rect 13890 21890 14959 21951
rect 13890 21856 13907 21890
rect 13941 21856 14907 21890
rect 14941 21856 14959 21890
rect 13890 21842 14959 21856
rect 14993 21857 15051 21951
rect 9422 21693 9439 21727
rect 9473 21693 9490 21727
rect 9422 21676 9490 21693
rect 10025 21729 10103 21763
rect 10137 21729 10213 21763
rect 10247 21729 10267 21763
rect 9841 21639 9899 21674
rect 9841 21605 9853 21639
rect 9887 21605 9899 21639
rect 9841 21546 9899 21605
rect 4965 21483 4983 21517
rect 5017 21483 5155 21517
rect 5189 21483 5207 21517
rect 4965 21441 5207 21483
rect 5426 21517 6495 21528
rect 5426 21483 5443 21517
rect 5477 21483 6443 21517
rect 6477 21483 6495 21517
rect 5426 21441 6495 21483
rect 6530 21517 7599 21528
rect 6530 21483 6547 21517
rect 6581 21483 7547 21517
rect 7581 21483 7599 21517
rect 6530 21441 7599 21483
rect 7634 21517 8703 21528
rect 7634 21483 7651 21517
rect 7685 21483 8651 21517
rect 8685 21483 8703 21517
rect 7634 21441 8703 21483
rect 8738 21517 9807 21528
rect 8738 21483 8755 21517
rect 8789 21483 9755 21517
rect 9789 21483 9807 21517
rect 8738 21441 9807 21483
rect 9841 21512 9853 21546
rect 9887 21512 9899 21546
rect 9841 21441 9899 21512
rect 10025 21659 10267 21729
rect 10301 21727 10543 21797
rect 10301 21693 10321 21727
rect 10355 21693 10431 21727
rect 10465 21693 10543 21727
rect 10896 21763 10966 21778
rect 10896 21729 10915 21763
rect 10949 21729 10966 21763
rect 10025 21619 10543 21659
rect 10025 21585 10043 21619
rect 10077 21585 10491 21619
rect 10525 21585 10543 21619
rect 10025 21517 10543 21585
rect 10896 21528 10966 21729
rect 11262 21727 11330 21842
rect 11262 21693 11279 21727
rect 11313 21693 11330 21727
rect 11262 21676 11330 21693
rect 12000 21763 12070 21778
rect 12000 21729 12019 21763
rect 12053 21729 12070 21763
rect 12000 21528 12070 21729
rect 12366 21727 12434 21842
rect 12366 21693 12383 21727
rect 12417 21693 12434 21727
rect 12366 21676 12434 21693
rect 13104 21763 13174 21778
rect 13104 21729 13123 21763
rect 13157 21729 13174 21763
rect 13104 21528 13174 21729
rect 13470 21727 13538 21842
rect 13470 21693 13487 21727
rect 13521 21693 13538 21727
rect 13470 21676 13538 21693
rect 14208 21763 14278 21778
rect 14208 21729 14227 21763
rect 14261 21729 14278 21763
rect 14208 21528 14278 21729
rect 14574 21727 14642 21842
rect 14993 21823 15005 21857
rect 15039 21823 15051 21857
rect 14993 21806 15051 21823
rect 15177 21883 15511 21951
rect 15177 21849 15195 21883
rect 15229 21849 15459 21883
rect 15493 21849 15511 21883
rect 15177 21797 15511 21849
rect 15546 21890 16615 21951
rect 15546 21856 15563 21890
rect 15597 21856 16563 21890
rect 16597 21856 16615 21890
rect 15546 21842 16615 21856
rect 16650 21890 17719 21951
rect 16650 21856 16667 21890
rect 16701 21856 17667 21890
rect 17701 21856 17719 21890
rect 16650 21842 17719 21856
rect 17754 21890 18823 21951
rect 17754 21856 17771 21890
rect 17805 21856 18771 21890
rect 18805 21856 18823 21890
rect 17754 21842 18823 21856
rect 18858 21890 19927 21951
rect 18858 21856 18875 21890
rect 18909 21856 19875 21890
rect 19909 21856 19927 21890
rect 18858 21842 19927 21856
rect 19961 21888 20203 21951
rect 19961 21854 19979 21888
rect 20013 21854 20151 21888
rect 20185 21854 20203 21888
rect 14574 21693 14591 21727
rect 14625 21693 14642 21727
rect 14574 21676 14642 21693
rect 15177 21729 15197 21763
rect 15231 21729 15327 21763
rect 14993 21639 15051 21674
rect 14993 21605 15005 21639
rect 15039 21605 15051 21639
rect 14993 21546 15051 21605
rect 10025 21483 10043 21517
rect 10077 21483 10491 21517
rect 10525 21483 10543 21517
rect 10025 21441 10543 21483
rect 10578 21517 11647 21528
rect 10578 21483 10595 21517
rect 10629 21483 11595 21517
rect 11629 21483 11647 21517
rect 10578 21441 11647 21483
rect 11682 21517 12751 21528
rect 11682 21483 11699 21517
rect 11733 21483 12699 21517
rect 12733 21483 12751 21517
rect 11682 21441 12751 21483
rect 12786 21517 13855 21528
rect 12786 21483 12803 21517
rect 12837 21483 13803 21517
rect 13837 21483 13855 21517
rect 12786 21441 13855 21483
rect 13890 21517 14959 21528
rect 13890 21483 13907 21517
rect 13941 21483 14907 21517
rect 14941 21483 14959 21517
rect 13890 21441 14959 21483
rect 14993 21512 15005 21546
rect 15039 21512 15051 21546
rect 14993 21441 15051 21512
rect 15177 21659 15327 21729
rect 15361 21727 15511 21797
rect 15361 21693 15457 21727
rect 15491 21693 15511 21727
rect 15864 21763 15934 21778
rect 15864 21729 15883 21763
rect 15917 21729 15934 21763
rect 15177 21619 15511 21659
rect 15177 21585 15195 21619
rect 15229 21585 15459 21619
rect 15493 21585 15511 21619
rect 15177 21517 15511 21585
rect 15864 21528 15934 21729
rect 16230 21727 16298 21842
rect 16230 21693 16247 21727
rect 16281 21693 16298 21727
rect 16230 21676 16298 21693
rect 16968 21763 17038 21778
rect 16968 21729 16987 21763
rect 17021 21729 17038 21763
rect 16968 21528 17038 21729
rect 17334 21727 17402 21842
rect 17334 21693 17351 21727
rect 17385 21693 17402 21727
rect 17334 21676 17402 21693
rect 18072 21763 18142 21778
rect 18072 21729 18091 21763
rect 18125 21729 18142 21763
rect 18072 21528 18142 21729
rect 18438 21727 18506 21842
rect 18438 21693 18455 21727
rect 18489 21693 18506 21727
rect 18438 21676 18506 21693
rect 19176 21763 19246 21778
rect 19176 21729 19195 21763
rect 19229 21729 19246 21763
rect 19176 21528 19246 21729
rect 19542 21727 19610 21842
rect 19961 21801 20203 21854
rect 19542 21693 19559 21727
rect 19593 21693 19610 21727
rect 19542 21676 19610 21693
rect 19961 21733 20011 21767
rect 20045 21733 20065 21767
rect 19961 21659 20065 21733
rect 20099 21727 20203 21801
rect 20099 21693 20119 21727
rect 20153 21693 20203 21727
rect 19961 21612 20203 21659
rect 19961 21578 19979 21612
rect 20013 21578 20151 21612
rect 20185 21578 20203 21612
rect 15177 21483 15195 21517
rect 15229 21483 15459 21517
rect 15493 21483 15511 21517
rect 15177 21441 15511 21483
rect 15546 21517 16615 21528
rect 15546 21483 15563 21517
rect 15597 21483 16563 21517
rect 16597 21483 16615 21517
rect 15546 21441 16615 21483
rect 16650 21517 17719 21528
rect 16650 21483 16667 21517
rect 16701 21483 17667 21517
rect 17701 21483 17719 21517
rect 16650 21441 17719 21483
rect 17754 21517 18823 21528
rect 17754 21483 17771 21517
rect 17805 21483 18771 21517
rect 18805 21483 18823 21517
rect 17754 21441 18823 21483
rect 18858 21517 19927 21528
rect 18858 21483 18875 21517
rect 18909 21483 19875 21517
rect 19909 21483 19927 21517
rect 18858 21441 19927 21483
rect 19961 21517 20203 21578
rect 19961 21483 19979 21517
rect 20013 21483 20151 21517
rect 20185 21483 20203 21517
rect 19961 21441 20203 21483
rect 4948 21407 4977 21441
rect 5011 21407 5069 21441
rect 5103 21407 5161 21441
rect 5195 21407 5253 21441
rect 5287 21407 5345 21441
rect 5379 21407 5437 21441
rect 5471 21407 5529 21441
rect 5563 21407 5621 21441
rect 5655 21407 5713 21441
rect 5747 21407 5805 21441
rect 5839 21407 5897 21441
rect 5931 21407 5989 21441
rect 6023 21407 6081 21441
rect 6115 21407 6173 21441
rect 6207 21407 6265 21441
rect 6299 21407 6357 21441
rect 6391 21407 6449 21441
rect 6483 21407 6541 21441
rect 6575 21407 6633 21441
rect 6667 21407 6725 21441
rect 6759 21407 6817 21441
rect 6851 21407 6909 21441
rect 6943 21407 7001 21441
rect 7035 21407 7093 21441
rect 7127 21407 7185 21441
rect 7219 21407 7277 21441
rect 7311 21407 7369 21441
rect 7403 21407 7461 21441
rect 7495 21407 7553 21441
rect 7587 21407 7645 21441
rect 7679 21407 7737 21441
rect 7771 21407 7829 21441
rect 7863 21407 7921 21441
rect 7955 21407 8013 21441
rect 8047 21407 8105 21441
rect 8139 21407 8197 21441
rect 8231 21407 8289 21441
rect 8323 21407 8381 21441
rect 8415 21407 8473 21441
rect 8507 21407 8565 21441
rect 8599 21407 8657 21441
rect 8691 21407 8749 21441
rect 8783 21407 8841 21441
rect 8875 21407 8933 21441
rect 8967 21407 9025 21441
rect 9059 21407 9117 21441
rect 9151 21407 9209 21441
rect 9243 21407 9301 21441
rect 9335 21407 9393 21441
rect 9427 21407 9485 21441
rect 9519 21407 9577 21441
rect 9611 21407 9669 21441
rect 9703 21407 9761 21441
rect 9795 21407 9853 21441
rect 9887 21407 9945 21441
rect 9979 21407 10037 21441
rect 10071 21407 10129 21441
rect 10163 21407 10221 21441
rect 10255 21407 10313 21441
rect 10347 21407 10405 21441
rect 10439 21407 10497 21441
rect 10531 21407 10589 21441
rect 10623 21407 10681 21441
rect 10715 21407 10773 21441
rect 10807 21407 10865 21441
rect 10899 21407 10957 21441
rect 10991 21407 11049 21441
rect 11083 21407 11141 21441
rect 11175 21407 11233 21441
rect 11267 21407 11325 21441
rect 11359 21407 11417 21441
rect 11451 21407 11509 21441
rect 11543 21407 11601 21441
rect 11635 21407 11693 21441
rect 11727 21407 11785 21441
rect 11819 21407 11877 21441
rect 11911 21407 11969 21441
rect 12003 21407 12061 21441
rect 12095 21407 12153 21441
rect 12187 21407 12245 21441
rect 12279 21407 12337 21441
rect 12371 21407 12429 21441
rect 12463 21407 12521 21441
rect 12555 21407 12613 21441
rect 12647 21407 12705 21441
rect 12739 21407 12797 21441
rect 12831 21407 12889 21441
rect 12923 21407 12981 21441
rect 13015 21407 13073 21441
rect 13107 21407 13165 21441
rect 13199 21407 13257 21441
rect 13291 21407 13349 21441
rect 13383 21407 13441 21441
rect 13475 21407 13533 21441
rect 13567 21407 13625 21441
rect 13659 21407 13717 21441
rect 13751 21407 13809 21441
rect 13843 21407 13901 21441
rect 13935 21407 13993 21441
rect 14027 21407 14085 21441
rect 14119 21407 14177 21441
rect 14211 21407 14269 21441
rect 14303 21407 14361 21441
rect 14395 21407 14453 21441
rect 14487 21407 14545 21441
rect 14579 21407 14637 21441
rect 14671 21407 14729 21441
rect 14763 21407 14821 21441
rect 14855 21407 14913 21441
rect 14947 21407 15005 21441
rect 15039 21407 15097 21441
rect 15131 21407 15189 21441
rect 15223 21407 15281 21441
rect 15315 21407 15373 21441
rect 15407 21407 15465 21441
rect 15499 21407 15557 21441
rect 15591 21407 15649 21441
rect 15683 21407 15741 21441
rect 15775 21407 15833 21441
rect 15867 21407 15925 21441
rect 15959 21407 16017 21441
rect 16051 21407 16109 21441
rect 16143 21407 16201 21441
rect 16235 21407 16293 21441
rect 16327 21407 16385 21441
rect 16419 21407 16477 21441
rect 16511 21407 16569 21441
rect 16603 21407 16661 21441
rect 16695 21407 16753 21441
rect 16787 21407 16845 21441
rect 16879 21407 16937 21441
rect 16971 21407 17029 21441
rect 17063 21407 17121 21441
rect 17155 21407 17213 21441
rect 17247 21407 17305 21441
rect 17339 21407 17397 21441
rect 17431 21407 17489 21441
rect 17523 21407 17581 21441
rect 17615 21407 17673 21441
rect 17707 21407 17765 21441
rect 17799 21407 17857 21441
rect 17891 21407 17949 21441
rect 17983 21407 18041 21441
rect 18075 21407 18133 21441
rect 18167 21407 18225 21441
rect 18259 21407 18317 21441
rect 18351 21407 18409 21441
rect 18443 21407 18501 21441
rect 18535 21407 18593 21441
rect 18627 21407 18685 21441
rect 18719 21407 18777 21441
rect 18811 21407 18869 21441
rect 18903 21407 18961 21441
rect 18995 21407 19053 21441
rect 19087 21407 19145 21441
rect 19179 21407 19237 21441
rect 19271 21407 19329 21441
rect 19363 21407 19421 21441
rect 19455 21407 19513 21441
rect 19547 21407 19605 21441
rect 19639 21407 19697 21441
rect 19731 21407 19789 21441
rect 19823 21407 19881 21441
rect 19915 21407 19973 21441
rect 20007 21407 20065 21441
rect 20099 21407 20157 21441
rect 20191 21407 20220 21441
rect 4965 21365 5207 21407
rect 4965 21331 4983 21365
rect 5017 21331 5155 21365
rect 5189 21331 5207 21365
rect 4965 21270 5207 21331
rect 4965 21236 4983 21270
rect 5017 21236 5155 21270
rect 5189 21236 5207 21270
rect 4965 21189 5207 21236
rect 4965 21121 5015 21155
rect 5049 21121 5069 21155
rect 4965 21047 5069 21121
rect 5103 21115 5207 21189
rect 5103 21081 5123 21115
rect 5157 21081 5207 21115
rect 5425 21365 6127 21407
rect 5425 21331 5443 21365
rect 5477 21331 6075 21365
rect 6109 21331 6127 21365
rect 5425 21263 6127 21331
rect 6162 21365 7231 21407
rect 6162 21331 6179 21365
rect 6213 21331 7179 21365
rect 7213 21331 7231 21365
rect 6162 21320 7231 21331
rect 7265 21336 7323 21407
rect 5425 21229 5443 21263
rect 5477 21229 6075 21263
rect 6109 21229 6127 21263
rect 5425 21189 6127 21229
rect 5425 21119 5763 21189
rect 5425 21085 5503 21119
rect 5537 21085 5606 21119
rect 5640 21085 5709 21119
rect 5743 21085 5763 21119
rect 5797 21121 5817 21155
rect 5851 21121 5916 21155
rect 5950 21121 6015 21155
rect 6049 21121 6127 21155
rect 5797 21051 6127 21121
rect 6480 21119 6550 21320
rect 7265 21302 7277 21336
rect 7311 21302 7323 21336
rect 7265 21243 7323 21302
rect 7265 21209 7277 21243
rect 7311 21209 7323 21243
rect 7265 21174 7323 21209
rect 7449 21365 7967 21407
rect 7449 21331 7467 21365
rect 7501 21331 7915 21365
rect 7949 21331 7967 21365
rect 7449 21263 7967 21331
rect 8002 21365 9071 21407
rect 8002 21331 8019 21365
rect 8053 21331 9019 21365
rect 9053 21331 9071 21365
rect 8002 21320 9071 21331
rect 9106 21365 10175 21407
rect 9106 21331 9123 21365
rect 9157 21331 10123 21365
rect 10157 21331 10175 21365
rect 9106 21320 10175 21331
rect 10210 21365 11279 21407
rect 10210 21331 10227 21365
rect 10261 21331 11227 21365
rect 11261 21331 11279 21365
rect 10210 21320 11279 21331
rect 11314 21365 12383 21407
rect 11314 21331 11331 21365
rect 11365 21331 12331 21365
rect 12365 21331 12383 21365
rect 11314 21320 12383 21331
rect 12417 21336 12475 21407
rect 7449 21229 7467 21263
rect 7501 21229 7915 21263
rect 7949 21229 7967 21263
rect 7449 21189 7967 21229
rect 6480 21085 6499 21119
rect 6533 21085 6550 21119
rect 6480 21070 6550 21085
rect 6846 21155 6914 21172
rect 6846 21121 6863 21155
rect 6897 21121 6914 21155
rect 4965 20994 5207 21047
rect 4965 20960 4983 20994
rect 5017 20960 5155 20994
rect 5189 20960 5207 20994
rect 4965 20897 5207 20960
rect 5425 20992 6127 21051
rect 6846 21006 6914 21121
rect 7449 21119 7691 21189
rect 7449 21085 7527 21119
rect 7561 21085 7637 21119
rect 7671 21085 7691 21119
rect 7725 21121 7745 21155
rect 7779 21121 7855 21155
rect 7889 21121 7967 21155
rect 7725 21051 7967 21121
rect 8320 21119 8390 21320
rect 8320 21085 8339 21119
rect 8373 21085 8390 21119
rect 8320 21070 8390 21085
rect 8686 21155 8754 21172
rect 8686 21121 8703 21155
rect 8737 21121 8754 21155
rect 7265 21025 7323 21042
rect 5425 20958 5443 20992
rect 5477 20958 6075 20992
rect 6109 20958 6127 20992
rect 5425 20897 6127 20958
rect 6162 20992 7231 21006
rect 6162 20958 6179 20992
rect 6213 20958 7179 20992
rect 7213 20958 7231 20992
rect 6162 20897 7231 20958
rect 7265 20991 7277 21025
rect 7311 20991 7323 21025
rect 7265 20897 7323 20991
rect 7449 20992 7967 21051
rect 8686 21006 8754 21121
rect 9424 21119 9494 21320
rect 9424 21085 9443 21119
rect 9477 21085 9494 21119
rect 9424 21070 9494 21085
rect 9790 21155 9858 21172
rect 9790 21121 9807 21155
rect 9841 21121 9858 21155
rect 9790 21006 9858 21121
rect 10528 21119 10598 21320
rect 10528 21085 10547 21119
rect 10581 21085 10598 21119
rect 10528 21070 10598 21085
rect 10894 21155 10962 21172
rect 10894 21121 10911 21155
rect 10945 21121 10962 21155
rect 10894 21006 10962 21121
rect 11632 21119 11702 21320
rect 12417 21302 12429 21336
rect 12463 21302 12475 21336
rect 12417 21243 12475 21302
rect 12417 21209 12429 21243
rect 12463 21209 12475 21243
rect 12417 21174 12475 21209
rect 12601 21365 13119 21407
rect 12601 21331 12619 21365
rect 12653 21331 13067 21365
rect 13101 21331 13119 21365
rect 12601 21263 13119 21331
rect 13154 21365 14223 21407
rect 13154 21331 13171 21365
rect 13205 21331 14171 21365
rect 14205 21331 14223 21365
rect 13154 21320 14223 21331
rect 14258 21365 15327 21407
rect 14258 21331 14275 21365
rect 14309 21331 15275 21365
rect 15309 21331 15327 21365
rect 14258 21320 15327 21331
rect 15362 21365 16431 21407
rect 15362 21331 15379 21365
rect 15413 21331 16379 21365
rect 16413 21331 16431 21365
rect 15362 21320 16431 21331
rect 16466 21365 17535 21407
rect 16466 21331 16483 21365
rect 16517 21331 17483 21365
rect 17517 21331 17535 21365
rect 16466 21320 17535 21331
rect 17569 21336 17627 21407
rect 12601 21229 12619 21263
rect 12653 21229 13067 21263
rect 13101 21229 13119 21263
rect 12601 21189 13119 21229
rect 11632 21085 11651 21119
rect 11685 21085 11702 21119
rect 11632 21070 11702 21085
rect 11998 21155 12066 21172
rect 11998 21121 12015 21155
rect 12049 21121 12066 21155
rect 11998 21006 12066 21121
rect 12601 21119 12843 21189
rect 12601 21085 12679 21119
rect 12713 21085 12789 21119
rect 12823 21085 12843 21119
rect 12877 21121 12897 21155
rect 12931 21121 13007 21155
rect 13041 21121 13119 21155
rect 12877 21051 13119 21121
rect 13472 21119 13542 21320
rect 13472 21085 13491 21119
rect 13525 21085 13542 21119
rect 13472 21070 13542 21085
rect 13838 21155 13906 21172
rect 13838 21121 13855 21155
rect 13889 21121 13906 21155
rect 12417 21025 12475 21042
rect 7449 20958 7467 20992
rect 7501 20958 7915 20992
rect 7949 20958 7967 20992
rect 7449 20897 7967 20958
rect 8002 20992 9071 21006
rect 8002 20958 8019 20992
rect 8053 20958 9019 20992
rect 9053 20958 9071 20992
rect 8002 20897 9071 20958
rect 9106 20992 10175 21006
rect 9106 20958 9123 20992
rect 9157 20958 10123 20992
rect 10157 20958 10175 20992
rect 9106 20897 10175 20958
rect 10210 20992 11279 21006
rect 10210 20958 10227 20992
rect 10261 20958 11227 20992
rect 11261 20958 11279 20992
rect 10210 20897 11279 20958
rect 11314 20992 12383 21006
rect 11314 20958 11331 20992
rect 11365 20958 12331 20992
rect 12365 20958 12383 20992
rect 11314 20897 12383 20958
rect 12417 20991 12429 21025
rect 12463 20991 12475 21025
rect 12417 20897 12475 20991
rect 12601 20992 13119 21051
rect 13838 21006 13906 21121
rect 14576 21119 14646 21320
rect 14576 21085 14595 21119
rect 14629 21085 14646 21119
rect 14576 21070 14646 21085
rect 14942 21155 15010 21172
rect 14942 21121 14959 21155
rect 14993 21121 15010 21155
rect 14942 21006 15010 21121
rect 15680 21119 15750 21320
rect 15680 21085 15699 21119
rect 15733 21085 15750 21119
rect 15680 21070 15750 21085
rect 16046 21155 16114 21172
rect 16046 21121 16063 21155
rect 16097 21121 16114 21155
rect 16046 21006 16114 21121
rect 16784 21119 16854 21320
rect 17569 21302 17581 21336
rect 17615 21302 17627 21336
rect 17754 21365 18823 21407
rect 17754 21331 17771 21365
rect 17805 21331 18771 21365
rect 18805 21331 18823 21365
rect 17754 21320 18823 21331
rect 18858 21365 19927 21407
rect 18858 21331 18875 21365
rect 18909 21331 19875 21365
rect 19909 21331 19927 21365
rect 18858 21320 19927 21331
rect 19961 21365 20203 21407
rect 19961 21331 19979 21365
rect 20013 21331 20151 21365
rect 20185 21331 20203 21365
rect 17569 21243 17627 21302
rect 17569 21209 17581 21243
rect 17615 21209 17627 21243
rect 17569 21174 17627 21209
rect 16784 21085 16803 21119
rect 16837 21085 16854 21119
rect 16784 21070 16854 21085
rect 17150 21155 17218 21172
rect 17150 21121 17167 21155
rect 17201 21121 17218 21155
rect 17150 21006 17218 21121
rect 18072 21119 18142 21320
rect 18072 21085 18091 21119
rect 18125 21085 18142 21119
rect 18072 21070 18142 21085
rect 18438 21155 18506 21172
rect 18438 21121 18455 21155
rect 18489 21121 18506 21155
rect 17569 21025 17627 21042
rect 12601 20958 12619 20992
rect 12653 20958 13067 20992
rect 13101 20958 13119 20992
rect 12601 20897 13119 20958
rect 13154 20992 14223 21006
rect 13154 20958 13171 20992
rect 13205 20958 14171 20992
rect 14205 20958 14223 20992
rect 13154 20897 14223 20958
rect 14258 20992 15327 21006
rect 14258 20958 14275 20992
rect 14309 20958 15275 20992
rect 15309 20958 15327 20992
rect 14258 20897 15327 20958
rect 15362 20992 16431 21006
rect 15362 20958 15379 20992
rect 15413 20958 16379 20992
rect 16413 20958 16431 20992
rect 15362 20897 16431 20958
rect 16466 20992 17535 21006
rect 16466 20958 16483 20992
rect 16517 20958 17483 20992
rect 17517 20958 17535 20992
rect 16466 20897 17535 20958
rect 17569 20991 17581 21025
rect 17615 20991 17627 21025
rect 18438 21006 18506 21121
rect 19176 21119 19246 21320
rect 19961 21270 20203 21331
rect 19961 21236 19979 21270
rect 20013 21236 20151 21270
rect 20185 21236 20203 21270
rect 19961 21189 20203 21236
rect 19176 21085 19195 21119
rect 19229 21085 19246 21119
rect 19176 21070 19246 21085
rect 19542 21155 19610 21172
rect 19542 21121 19559 21155
rect 19593 21121 19610 21155
rect 19542 21006 19610 21121
rect 19961 21115 20065 21189
rect 19961 21081 20011 21115
rect 20045 21081 20065 21115
rect 20099 21121 20119 21155
rect 20153 21121 20203 21155
rect 20099 21047 20203 21121
rect 17569 20897 17627 20991
rect 17754 20992 18823 21006
rect 17754 20958 17771 20992
rect 17805 20958 18771 20992
rect 18805 20958 18823 20992
rect 17754 20897 18823 20958
rect 18858 20992 19927 21006
rect 18858 20958 18875 20992
rect 18909 20958 19875 20992
rect 19909 20958 19927 20992
rect 18858 20897 19927 20958
rect 19961 20994 20203 21047
rect 19961 20960 19979 20994
rect 20013 20960 20151 20994
rect 20185 20960 20203 20994
rect 19961 20897 20203 20960
rect 4948 20863 4977 20897
rect 5011 20863 5069 20897
rect 5103 20863 5161 20897
rect 5195 20863 5253 20897
rect 5287 20863 5345 20897
rect 5379 20863 5437 20897
rect 5471 20863 5529 20897
rect 5563 20863 5621 20897
rect 5655 20863 5713 20897
rect 5747 20863 5805 20897
rect 5839 20863 5897 20897
rect 5931 20863 5989 20897
rect 6023 20863 6081 20897
rect 6115 20863 6173 20897
rect 6207 20863 6265 20897
rect 6299 20863 6357 20897
rect 6391 20863 6449 20897
rect 6483 20863 6541 20897
rect 6575 20863 6633 20897
rect 6667 20863 6725 20897
rect 6759 20863 6817 20897
rect 6851 20863 6909 20897
rect 6943 20863 7001 20897
rect 7035 20863 7093 20897
rect 7127 20863 7185 20897
rect 7219 20863 7277 20897
rect 7311 20863 7369 20897
rect 7403 20863 7461 20897
rect 7495 20863 7553 20897
rect 7587 20863 7645 20897
rect 7679 20863 7737 20897
rect 7771 20863 7829 20897
rect 7863 20863 7921 20897
rect 7955 20863 8013 20897
rect 8047 20863 8105 20897
rect 8139 20863 8197 20897
rect 8231 20863 8289 20897
rect 8323 20863 8381 20897
rect 8415 20863 8473 20897
rect 8507 20863 8565 20897
rect 8599 20863 8657 20897
rect 8691 20863 8749 20897
rect 8783 20863 8841 20897
rect 8875 20863 8933 20897
rect 8967 20863 9025 20897
rect 9059 20863 9117 20897
rect 9151 20863 9209 20897
rect 9243 20863 9301 20897
rect 9335 20863 9393 20897
rect 9427 20863 9485 20897
rect 9519 20863 9577 20897
rect 9611 20863 9669 20897
rect 9703 20863 9761 20897
rect 9795 20863 9853 20897
rect 9887 20863 9945 20897
rect 9979 20863 10037 20897
rect 10071 20863 10129 20897
rect 10163 20863 10221 20897
rect 10255 20863 10313 20897
rect 10347 20863 10405 20897
rect 10439 20863 10497 20897
rect 10531 20863 10589 20897
rect 10623 20863 10681 20897
rect 10715 20863 10773 20897
rect 10807 20863 10865 20897
rect 10899 20863 10957 20897
rect 10991 20863 11049 20897
rect 11083 20863 11141 20897
rect 11175 20863 11233 20897
rect 11267 20863 11325 20897
rect 11359 20863 11417 20897
rect 11451 20863 11509 20897
rect 11543 20863 11601 20897
rect 11635 20863 11693 20897
rect 11727 20863 11785 20897
rect 11819 20863 11877 20897
rect 11911 20863 11969 20897
rect 12003 20863 12061 20897
rect 12095 20863 12153 20897
rect 12187 20863 12245 20897
rect 12279 20863 12337 20897
rect 12371 20863 12429 20897
rect 12463 20863 12521 20897
rect 12555 20863 12613 20897
rect 12647 20863 12705 20897
rect 12739 20863 12797 20897
rect 12831 20863 12889 20897
rect 12923 20863 12981 20897
rect 13015 20863 13073 20897
rect 13107 20863 13165 20897
rect 13199 20863 13257 20897
rect 13291 20863 13349 20897
rect 13383 20863 13441 20897
rect 13475 20863 13533 20897
rect 13567 20863 13625 20897
rect 13659 20863 13717 20897
rect 13751 20863 13809 20897
rect 13843 20863 13901 20897
rect 13935 20863 13993 20897
rect 14027 20863 14085 20897
rect 14119 20863 14177 20897
rect 14211 20863 14269 20897
rect 14303 20863 14361 20897
rect 14395 20863 14453 20897
rect 14487 20863 14545 20897
rect 14579 20863 14637 20897
rect 14671 20863 14729 20897
rect 14763 20863 14821 20897
rect 14855 20863 14913 20897
rect 14947 20863 15005 20897
rect 15039 20863 15097 20897
rect 15131 20863 15189 20897
rect 15223 20863 15281 20897
rect 15315 20863 15373 20897
rect 15407 20863 15465 20897
rect 15499 20863 15557 20897
rect 15591 20863 15649 20897
rect 15683 20863 15741 20897
rect 15775 20863 15833 20897
rect 15867 20863 15925 20897
rect 15959 20863 16017 20897
rect 16051 20863 16109 20897
rect 16143 20863 16201 20897
rect 16235 20863 16293 20897
rect 16327 20863 16385 20897
rect 16419 20863 16477 20897
rect 16511 20863 16569 20897
rect 16603 20863 16661 20897
rect 16695 20863 16753 20897
rect 16787 20863 16845 20897
rect 16879 20863 16937 20897
rect 16971 20863 17029 20897
rect 17063 20863 17121 20897
rect 17155 20863 17213 20897
rect 17247 20863 17305 20897
rect 17339 20863 17397 20897
rect 17431 20863 17489 20897
rect 17523 20863 17581 20897
rect 17615 20863 17673 20897
rect 17707 20863 17765 20897
rect 17799 20863 17857 20897
rect 17891 20863 17949 20897
rect 17983 20863 18041 20897
rect 18075 20863 18133 20897
rect 18167 20863 18225 20897
rect 18259 20863 18317 20897
rect 18351 20863 18409 20897
rect 18443 20863 18501 20897
rect 18535 20863 18593 20897
rect 18627 20863 18685 20897
rect 18719 20863 18777 20897
rect 18811 20863 18869 20897
rect 18903 20863 18961 20897
rect 18995 20863 19053 20897
rect 19087 20863 19145 20897
rect 19179 20863 19237 20897
rect 19271 20863 19329 20897
rect 19363 20863 19421 20897
rect 19455 20863 19513 20897
rect 19547 20863 19605 20897
rect 19639 20863 19697 20897
rect 19731 20863 19789 20897
rect 19823 20863 19881 20897
rect 19915 20863 19973 20897
rect 20007 20863 20065 20897
rect 20099 20863 20157 20897
rect 20191 20863 20220 20897
rect 4965 20800 5207 20863
rect 4965 20766 4983 20800
rect 5017 20766 5155 20800
rect 5189 20766 5207 20800
rect 4965 20713 5207 20766
rect 5426 20802 6495 20863
rect 5426 20768 5443 20802
rect 5477 20768 6443 20802
rect 6477 20768 6495 20802
rect 5426 20754 6495 20768
rect 6530 20802 7599 20863
rect 6530 20768 6547 20802
rect 6581 20768 7547 20802
rect 7581 20768 7599 20802
rect 6530 20754 7599 20768
rect 7634 20802 8703 20863
rect 7634 20768 7651 20802
rect 7685 20768 8651 20802
rect 8685 20768 8703 20802
rect 7634 20754 8703 20768
rect 8738 20802 9807 20863
rect 8738 20768 8755 20802
rect 8789 20768 9755 20802
rect 9789 20768 9807 20802
rect 8738 20754 9807 20768
rect 9841 20769 9899 20863
rect 4965 20639 5069 20713
rect 4965 20605 5015 20639
rect 5049 20605 5069 20639
rect 5103 20645 5123 20679
rect 5157 20645 5207 20679
rect 5103 20571 5207 20645
rect 4965 20524 5207 20571
rect 4965 20490 4983 20524
rect 5017 20490 5155 20524
rect 5189 20490 5207 20524
rect 4965 20429 5207 20490
rect 5744 20675 5814 20690
rect 5744 20641 5763 20675
rect 5797 20641 5814 20675
rect 5744 20440 5814 20641
rect 6110 20639 6178 20754
rect 6110 20605 6127 20639
rect 6161 20605 6178 20639
rect 6110 20588 6178 20605
rect 6848 20675 6918 20690
rect 6848 20641 6867 20675
rect 6901 20641 6918 20675
rect 6848 20440 6918 20641
rect 7214 20639 7282 20754
rect 7214 20605 7231 20639
rect 7265 20605 7282 20639
rect 7214 20588 7282 20605
rect 7952 20675 8022 20690
rect 7952 20641 7971 20675
rect 8005 20641 8022 20675
rect 7952 20440 8022 20641
rect 8318 20639 8386 20754
rect 8318 20605 8335 20639
rect 8369 20605 8386 20639
rect 8318 20588 8386 20605
rect 9056 20675 9126 20690
rect 9056 20641 9075 20675
rect 9109 20641 9126 20675
rect 9056 20440 9126 20641
rect 9422 20639 9490 20754
rect 9841 20735 9853 20769
rect 9887 20735 9899 20769
rect 9841 20718 9899 20735
rect 10025 20802 10543 20863
rect 10025 20768 10043 20802
rect 10077 20768 10491 20802
rect 10525 20768 10543 20802
rect 10025 20709 10543 20768
rect 10578 20802 11647 20863
rect 10578 20768 10595 20802
rect 10629 20768 11595 20802
rect 11629 20768 11647 20802
rect 10578 20754 11647 20768
rect 11682 20802 12751 20863
rect 11682 20768 11699 20802
rect 11733 20768 12699 20802
rect 12733 20768 12751 20802
rect 11682 20754 12751 20768
rect 12786 20802 13855 20863
rect 12786 20768 12803 20802
rect 12837 20768 13803 20802
rect 13837 20768 13855 20802
rect 12786 20754 13855 20768
rect 13890 20802 14959 20863
rect 13890 20768 13907 20802
rect 13941 20768 14907 20802
rect 14941 20768 14959 20802
rect 13890 20754 14959 20768
rect 14993 20769 15051 20863
rect 9422 20605 9439 20639
rect 9473 20605 9490 20639
rect 9422 20588 9490 20605
rect 10025 20641 10103 20675
rect 10137 20641 10213 20675
rect 10247 20641 10267 20675
rect 9841 20551 9899 20586
rect 9841 20517 9853 20551
rect 9887 20517 9899 20551
rect 9841 20458 9899 20517
rect 4965 20395 4983 20429
rect 5017 20395 5155 20429
rect 5189 20395 5207 20429
rect 4965 20353 5207 20395
rect 5426 20429 6495 20440
rect 5426 20395 5443 20429
rect 5477 20395 6443 20429
rect 6477 20395 6495 20429
rect 5426 20353 6495 20395
rect 6530 20429 7599 20440
rect 6530 20395 6547 20429
rect 6581 20395 7547 20429
rect 7581 20395 7599 20429
rect 6530 20353 7599 20395
rect 7634 20429 8703 20440
rect 7634 20395 7651 20429
rect 7685 20395 8651 20429
rect 8685 20395 8703 20429
rect 7634 20353 8703 20395
rect 8738 20429 9807 20440
rect 8738 20395 8755 20429
rect 8789 20395 9755 20429
rect 9789 20395 9807 20429
rect 8738 20353 9807 20395
rect 9841 20424 9853 20458
rect 9887 20424 9899 20458
rect 9841 20353 9899 20424
rect 10025 20571 10267 20641
rect 10301 20639 10543 20709
rect 10301 20605 10321 20639
rect 10355 20605 10431 20639
rect 10465 20605 10543 20639
rect 10896 20675 10966 20690
rect 10896 20641 10915 20675
rect 10949 20641 10966 20675
rect 10025 20531 10543 20571
rect 10025 20497 10043 20531
rect 10077 20497 10491 20531
rect 10525 20497 10543 20531
rect 10025 20429 10543 20497
rect 10896 20440 10966 20641
rect 11262 20639 11330 20754
rect 11262 20605 11279 20639
rect 11313 20605 11330 20639
rect 11262 20588 11330 20605
rect 12000 20675 12070 20690
rect 12000 20641 12019 20675
rect 12053 20641 12070 20675
rect 12000 20440 12070 20641
rect 12366 20639 12434 20754
rect 12366 20605 12383 20639
rect 12417 20605 12434 20639
rect 12366 20588 12434 20605
rect 13104 20675 13174 20690
rect 13104 20641 13123 20675
rect 13157 20641 13174 20675
rect 13104 20440 13174 20641
rect 13470 20639 13538 20754
rect 13470 20605 13487 20639
rect 13521 20605 13538 20639
rect 13470 20588 13538 20605
rect 14208 20675 14278 20690
rect 14208 20641 14227 20675
rect 14261 20641 14278 20675
rect 14208 20440 14278 20641
rect 14574 20639 14642 20754
rect 14993 20735 15005 20769
rect 15039 20735 15051 20769
rect 14993 20718 15051 20735
rect 15177 20795 15511 20863
rect 15177 20761 15195 20795
rect 15229 20761 15459 20795
rect 15493 20761 15511 20795
rect 15177 20709 15511 20761
rect 15546 20802 16615 20863
rect 15546 20768 15563 20802
rect 15597 20768 16563 20802
rect 16597 20768 16615 20802
rect 15546 20754 16615 20768
rect 16650 20802 17719 20863
rect 16650 20768 16667 20802
rect 16701 20768 17667 20802
rect 17701 20768 17719 20802
rect 16650 20754 17719 20768
rect 17754 20802 18823 20863
rect 17754 20768 17771 20802
rect 17805 20768 18771 20802
rect 18805 20768 18823 20802
rect 17754 20754 18823 20768
rect 18858 20802 19927 20863
rect 18858 20768 18875 20802
rect 18909 20768 19875 20802
rect 19909 20768 19927 20802
rect 18858 20754 19927 20768
rect 19961 20800 20203 20863
rect 19961 20766 19979 20800
rect 20013 20766 20151 20800
rect 20185 20766 20203 20800
rect 14574 20605 14591 20639
rect 14625 20605 14642 20639
rect 14574 20588 14642 20605
rect 15177 20641 15197 20675
rect 15231 20641 15327 20675
rect 14993 20551 15051 20586
rect 14993 20517 15005 20551
rect 15039 20517 15051 20551
rect 14993 20458 15051 20517
rect 10025 20395 10043 20429
rect 10077 20395 10491 20429
rect 10525 20395 10543 20429
rect 10025 20353 10543 20395
rect 10578 20429 11647 20440
rect 10578 20395 10595 20429
rect 10629 20395 11595 20429
rect 11629 20395 11647 20429
rect 10578 20353 11647 20395
rect 11682 20429 12751 20440
rect 11682 20395 11699 20429
rect 11733 20395 12699 20429
rect 12733 20395 12751 20429
rect 11682 20353 12751 20395
rect 12786 20429 13855 20440
rect 12786 20395 12803 20429
rect 12837 20395 13803 20429
rect 13837 20395 13855 20429
rect 12786 20353 13855 20395
rect 13890 20429 14959 20440
rect 13890 20395 13907 20429
rect 13941 20395 14907 20429
rect 14941 20395 14959 20429
rect 13890 20353 14959 20395
rect 14993 20424 15005 20458
rect 15039 20424 15051 20458
rect 14993 20353 15051 20424
rect 15177 20571 15327 20641
rect 15361 20639 15511 20709
rect 15361 20605 15457 20639
rect 15491 20605 15511 20639
rect 15864 20675 15934 20690
rect 15864 20641 15883 20675
rect 15917 20641 15934 20675
rect 15177 20531 15511 20571
rect 15177 20497 15195 20531
rect 15229 20497 15459 20531
rect 15493 20497 15511 20531
rect 15177 20429 15511 20497
rect 15864 20440 15934 20641
rect 16230 20639 16298 20754
rect 16230 20605 16247 20639
rect 16281 20605 16298 20639
rect 16230 20588 16298 20605
rect 16968 20675 17038 20690
rect 16968 20641 16987 20675
rect 17021 20641 17038 20675
rect 16968 20440 17038 20641
rect 17334 20639 17402 20754
rect 17334 20605 17351 20639
rect 17385 20605 17402 20639
rect 17334 20588 17402 20605
rect 18072 20675 18142 20690
rect 18072 20641 18091 20675
rect 18125 20641 18142 20675
rect 18072 20440 18142 20641
rect 18438 20639 18506 20754
rect 18438 20605 18455 20639
rect 18489 20605 18506 20639
rect 18438 20588 18506 20605
rect 19176 20675 19246 20690
rect 19176 20641 19195 20675
rect 19229 20641 19246 20675
rect 19176 20440 19246 20641
rect 19542 20639 19610 20754
rect 19961 20713 20203 20766
rect 19542 20605 19559 20639
rect 19593 20605 19610 20639
rect 19542 20588 19610 20605
rect 19961 20645 20011 20679
rect 20045 20645 20065 20679
rect 19961 20571 20065 20645
rect 20099 20639 20203 20713
rect 20099 20605 20119 20639
rect 20153 20605 20203 20639
rect 19961 20524 20203 20571
rect 19961 20490 19979 20524
rect 20013 20490 20151 20524
rect 20185 20490 20203 20524
rect 15177 20395 15195 20429
rect 15229 20395 15459 20429
rect 15493 20395 15511 20429
rect 15177 20353 15511 20395
rect 15546 20429 16615 20440
rect 15546 20395 15563 20429
rect 15597 20395 16563 20429
rect 16597 20395 16615 20429
rect 15546 20353 16615 20395
rect 16650 20429 17719 20440
rect 16650 20395 16667 20429
rect 16701 20395 17667 20429
rect 17701 20395 17719 20429
rect 16650 20353 17719 20395
rect 17754 20429 18823 20440
rect 17754 20395 17771 20429
rect 17805 20395 18771 20429
rect 18805 20395 18823 20429
rect 17754 20353 18823 20395
rect 18858 20429 19927 20440
rect 18858 20395 18875 20429
rect 18909 20395 19875 20429
rect 19909 20395 19927 20429
rect 18858 20353 19927 20395
rect 19961 20429 20203 20490
rect 19961 20395 19979 20429
rect 20013 20395 20151 20429
rect 20185 20395 20203 20429
rect 19961 20353 20203 20395
rect 4948 20319 4977 20353
rect 5011 20319 5069 20353
rect 5103 20319 5161 20353
rect 5195 20319 5253 20353
rect 5287 20319 5345 20353
rect 5379 20319 5437 20353
rect 5471 20319 5529 20353
rect 5563 20319 5621 20353
rect 5655 20319 5713 20353
rect 5747 20319 5805 20353
rect 5839 20319 5897 20353
rect 5931 20319 5989 20353
rect 6023 20319 6081 20353
rect 6115 20319 6173 20353
rect 6207 20319 6265 20353
rect 6299 20319 6357 20353
rect 6391 20319 6449 20353
rect 6483 20319 6541 20353
rect 6575 20319 6633 20353
rect 6667 20319 6725 20353
rect 6759 20319 6817 20353
rect 6851 20319 6909 20353
rect 6943 20319 7001 20353
rect 7035 20319 7093 20353
rect 7127 20319 7185 20353
rect 7219 20319 7277 20353
rect 7311 20319 7369 20353
rect 7403 20319 7461 20353
rect 7495 20319 7553 20353
rect 7587 20319 7645 20353
rect 7679 20319 7737 20353
rect 7771 20319 7829 20353
rect 7863 20319 7921 20353
rect 7955 20319 8013 20353
rect 8047 20319 8105 20353
rect 8139 20319 8197 20353
rect 8231 20319 8289 20353
rect 8323 20319 8381 20353
rect 8415 20319 8473 20353
rect 8507 20319 8565 20353
rect 8599 20319 8657 20353
rect 8691 20319 8749 20353
rect 8783 20319 8841 20353
rect 8875 20319 8933 20353
rect 8967 20319 9025 20353
rect 9059 20319 9117 20353
rect 9151 20319 9209 20353
rect 9243 20319 9301 20353
rect 9335 20319 9393 20353
rect 9427 20319 9485 20353
rect 9519 20319 9577 20353
rect 9611 20319 9669 20353
rect 9703 20319 9761 20353
rect 9795 20319 9853 20353
rect 9887 20319 9945 20353
rect 9979 20319 10037 20353
rect 10071 20319 10129 20353
rect 10163 20319 10221 20353
rect 10255 20319 10313 20353
rect 10347 20319 10405 20353
rect 10439 20319 10497 20353
rect 10531 20319 10589 20353
rect 10623 20319 10681 20353
rect 10715 20319 10773 20353
rect 10807 20319 10865 20353
rect 10899 20319 10957 20353
rect 10991 20319 11049 20353
rect 11083 20319 11141 20353
rect 11175 20319 11233 20353
rect 11267 20319 11325 20353
rect 11359 20319 11417 20353
rect 11451 20319 11509 20353
rect 11543 20319 11601 20353
rect 11635 20319 11693 20353
rect 11727 20319 11785 20353
rect 11819 20319 11877 20353
rect 11911 20319 11969 20353
rect 12003 20319 12061 20353
rect 12095 20319 12153 20353
rect 12187 20319 12245 20353
rect 12279 20319 12337 20353
rect 12371 20319 12429 20353
rect 12463 20319 12521 20353
rect 12555 20319 12613 20353
rect 12647 20319 12705 20353
rect 12739 20319 12797 20353
rect 12831 20319 12889 20353
rect 12923 20319 12981 20353
rect 13015 20319 13073 20353
rect 13107 20319 13165 20353
rect 13199 20319 13257 20353
rect 13291 20319 13349 20353
rect 13383 20319 13441 20353
rect 13475 20319 13533 20353
rect 13567 20319 13625 20353
rect 13659 20319 13717 20353
rect 13751 20319 13809 20353
rect 13843 20319 13901 20353
rect 13935 20319 13993 20353
rect 14027 20319 14085 20353
rect 14119 20319 14177 20353
rect 14211 20319 14269 20353
rect 14303 20319 14361 20353
rect 14395 20319 14453 20353
rect 14487 20319 14545 20353
rect 14579 20319 14637 20353
rect 14671 20319 14729 20353
rect 14763 20319 14821 20353
rect 14855 20319 14913 20353
rect 14947 20319 15005 20353
rect 15039 20319 15097 20353
rect 15131 20319 15189 20353
rect 15223 20319 15281 20353
rect 15315 20319 15373 20353
rect 15407 20319 15465 20353
rect 15499 20319 15557 20353
rect 15591 20319 15649 20353
rect 15683 20319 15741 20353
rect 15775 20319 15833 20353
rect 15867 20319 15925 20353
rect 15959 20319 16017 20353
rect 16051 20319 16109 20353
rect 16143 20319 16201 20353
rect 16235 20319 16293 20353
rect 16327 20319 16385 20353
rect 16419 20319 16477 20353
rect 16511 20319 16569 20353
rect 16603 20319 16661 20353
rect 16695 20319 16753 20353
rect 16787 20319 16845 20353
rect 16879 20319 16937 20353
rect 16971 20319 17029 20353
rect 17063 20319 17121 20353
rect 17155 20319 17213 20353
rect 17247 20319 17305 20353
rect 17339 20319 17397 20353
rect 17431 20319 17489 20353
rect 17523 20319 17581 20353
rect 17615 20319 17673 20353
rect 17707 20319 17765 20353
rect 17799 20319 17857 20353
rect 17891 20319 17949 20353
rect 17983 20319 18041 20353
rect 18075 20319 18133 20353
rect 18167 20319 18225 20353
rect 18259 20319 18317 20353
rect 18351 20319 18409 20353
rect 18443 20319 18501 20353
rect 18535 20319 18593 20353
rect 18627 20319 18685 20353
rect 18719 20319 18777 20353
rect 18811 20319 18869 20353
rect 18903 20319 18961 20353
rect 18995 20319 19053 20353
rect 19087 20319 19145 20353
rect 19179 20319 19237 20353
rect 19271 20319 19329 20353
rect 19363 20319 19421 20353
rect 19455 20319 19513 20353
rect 19547 20319 19605 20353
rect 19639 20319 19697 20353
rect 19731 20319 19789 20353
rect 19823 20319 19881 20353
rect 19915 20319 19973 20353
rect 20007 20319 20065 20353
rect 20099 20319 20157 20353
rect 20191 20319 20220 20353
rect 4965 20277 5207 20319
rect 4965 20243 4983 20277
rect 5017 20243 5155 20277
rect 5189 20243 5207 20277
rect 4965 20182 5207 20243
rect 4965 20148 4983 20182
rect 5017 20148 5155 20182
rect 5189 20148 5207 20182
rect 4965 20101 5207 20148
rect 4965 20033 5015 20067
rect 5049 20033 5069 20067
rect 4965 19959 5069 20033
rect 5103 20027 5207 20101
rect 5103 19993 5123 20027
rect 5157 19993 5207 20027
rect 5425 20277 6127 20319
rect 5425 20243 5443 20277
rect 5477 20243 6075 20277
rect 6109 20243 6127 20277
rect 5425 20175 6127 20243
rect 6162 20277 7231 20319
rect 6162 20243 6179 20277
rect 6213 20243 7179 20277
rect 7213 20243 7231 20277
rect 6162 20232 7231 20243
rect 7265 20248 7323 20319
rect 5425 20141 5443 20175
rect 5477 20141 6075 20175
rect 6109 20141 6127 20175
rect 5425 20101 6127 20141
rect 5425 20031 5763 20101
rect 5425 19997 5503 20031
rect 5537 19997 5606 20031
rect 5640 19997 5709 20031
rect 5743 19997 5763 20031
rect 5797 20033 5817 20067
rect 5851 20033 5916 20067
rect 5950 20033 6015 20067
rect 6049 20033 6127 20067
rect 5797 19963 6127 20033
rect 6480 20031 6550 20232
rect 7265 20214 7277 20248
rect 7311 20214 7323 20248
rect 7265 20155 7323 20214
rect 7265 20121 7277 20155
rect 7311 20121 7323 20155
rect 7265 20086 7323 20121
rect 7449 20277 7967 20319
rect 7449 20243 7467 20277
rect 7501 20243 7915 20277
rect 7949 20243 7967 20277
rect 7449 20175 7967 20243
rect 8002 20277 9071 20319
rect 8002 20243 8019 20277
rect 8053 20243 9019 20277
rect 9053 20243 9071 20277
rect 8002 20232 9071 20243
rect 9106 20277 10175 20319
rect 9106 20243 9123 20277
rect 9157 20243 10123 20277
rect 10157 20243 10175 20277
rect 9106 20232 10175 20243
rect 10210 20277 11279 20319
rect 10210 20243 10227 20277
rect 10261 20243 11227 20277
rect 11261 20243 11279 20277
rect 10210 20232 11279 20243
rect 11314 20277 12383 20319
rect 11314 20243 11331 20277
rect 11365 20243 12331 20277
rect 12365 20243 12383 20277
rect 11314 20232 12383 20243
rect 12417 20248 12475 20319
rect 7449 20141 7467 20175
rect 7501 20141 7915 20175
rect 7949 20141 7967 20175
rect 7449 20101 7967 20141
rect 6480 19997 6499 20031
rect 6533 19997 6550 20031
rect 6480 19982 6550 19997
rect 6846 20067 6914 20084
rect 6846 20033 6863 20067
rect 6897 20033 6914 20067
rect 4965 19906 5207 19959
rect 4965 19872 4983 19906
rect 5017 19872 5155 19906
rect 5189 19872 5207 19906
rect 4965 19809 5207 19872
rect 5425 19904 6127 19963
rect 6846 19918 6914 20033
rect 7449 20031 7691 20101
rect 7449 19997 7527 20031
rect 7561 19997 7637 20031
rect 7671 19997 7691 20031
rect 7725 20033 7745 20067
rect 7779 20033 7855 20067
rect 7889 20033 7967 20067
rect 7725 19963 7967 20033
rect 8320 20031 8390 20232
rect 8320 19997 8339 20031
rect 8373 19997 8390 20031
rect 8320 19982 8390 19997
rect 8686 20067 8754 20084
rect 8686 20033 8703 20067
rect 8737 20033 8754 20067
rect 7265 19937 7323 19954
rect 5425 19870 5443 19904
rect 5477 19870 6075 19904
rect 6109 19870 6127 19904
rect 5425 19809 6127 19870
rect 6162 19904 7231 19918
rect 6162 19870 6179 19904
rect 6213 19870 7179 19904
rect 7213 19870 7231 19904
rect 6162 19809 7231 19870
rect 7265 19903 7277 19937
rect 7311 19903 7323 19937
rect 7265 19809 7323 19903
rect 7449 19904 7967 19963
rect 8686 19918 8754 20033
rect 9424 20031 9494 20232
rect 9424 19997 9443 20031
rect 9477 19997 9494 20031
rect 9424 19982 9494 19997
rect 9790 20067 9858 20084
rect 9790 20033 9807 20067
rect 9841 20033 9858 20067
rect 9790 19918 9858 20033
rect 10528 20031 10598 20232
rect 10528 19997 10547 20031
rect 10581 19997 10598 20031
rect 10528 19982 10598 19997
rect 10894 20067 10962 20084
rect 10894 20033 10911 20067
rect 10945 20033 10962 20067
rect 10894 19918 10962 20033
rect 11632 20031 11702 20232
rect 12417 20214 12429 20248
rect 12463 20214 12475 20248
rect 12417 20155 12475 20214
rect 12417 20121 12429 20155
rect 12463 20121 12475 20155
rect 12417 20086 12475 20121
rect 12601 20277 13119 20319
rect 12601 20243 12619 20277
rect 12653 20243 13067 20277
rect 13101 20243 13119 20277
rect 12601 20175 13119 20243
rect 13154 20277 14223 20319
rect 13154 20243 13171 20277
rect 13205 20243 14171 20277
rect 14205 20243 14223 20277
rect 13154 20232 14223 20243
rect 14258 20277 15327 20319
rect 14258 20243 14275 20277
rect 14309 20243 15275 20277
rect 15309 20243 15327 20277
rect 14258 20232 15327 20243
rect 15362 20277 16431 20319
rect 15362 20243 15379 20277
rect 15413 20243 16379 20277
rect 16413 20243 16431 20277
rect 15362 20232 16431 20243
rect 16466 20277 17535 20319
rect 16466 20243 16483 20277
rect 16517 20243 17483 20277
rect 17517 20243 17535 20277
rect 16466 20232 17535 20243
rect 17569 20248 17627 20319
rect 12601 20141 12619 20175
rect 12653 20141 13067 20175
rect 13101 20141 13119 20175
rect 12601 20101 13119 20141
rect 11632 19997 11651 20031
rect 11685 19997 11702 20031
rect 11632 19982 11702 19997
rect 11998 20067 12066 20084
rect 11998 20033 12015 20067
rect 12049 20033 12066 20067
rect 11998 19918 12066 20033
rect 12601 20031 12843 20101
rect 12601 19997 12679 20031
rect 12713 19997 12789 20031
rect 12823 19997 12843 20031
rect 12877 20033 12897 20067
rect 12931 20033 13007 20067
rect 13041 20033 13119 20067
rect 12877 19963 13119 20033
rect 13472 20031 13542 20232
rect 13472 19997 13491 20031
rect 13525 19997 13542 20031
rect 13472 19982 13542 19997
rect 13838 20067 13906 20084
rect 13838 20033 13855 20067
rect 13889 20033 13906 20067
rect 12417 19937 12475 19954
rect 7449 19870 7467 19904
rect 7501 19870 7915 19904
rect 7949 19870 7967 19904
rect 7449 19809 7967 19870
rect 8002 19904 9071 19918
rect 8002 19870 8019 19904
rect 8053 19870 9019 19904
rect 9053 19870 9071 19904
rect 8002 19809 9071 19870
rect 9106 19904 10175 19918
rect 9106 19870 9123 19904
rect 9157 19870 10123 19904
rect 10157 19870 10175 19904
rect 9106 19809 10175 19870
rect 10210 19904 11279 19918
rect 10210 19870 10227 19904
rect 10261 19870 11227 19904
rect 11261 19870 11279 19904
rect 10210 19809 11279 19870
rect 11314 19904 12383 19918
rect 11314 19870 11331 19904
rect 11365 19870 12331 19904
rect 12365 19870 12383 19904
rect 11314 19809 12383 19870
rect 12417 19903 12429 19937
rect 12463 19903 12475 19937
rect 12417 19809 12475 19903
rect 12601 19904 13119 19963
rect 13838 19918 13906 20033
rect 14576 20031 14646 20232
rect 14576 19997 14595 20031
rect 14629 19997 14646 20031
rect 14576 19982 14646 19997
rect 14942 20067 15010 20084
rect 14942 20033 14959 20067
rect 14993 20033 15010 20067
rect 14942 19918 15010 20033
rect 15680 20031 15750 20232
rect 15680 19997 15699 20031
rect 15733 19997 15750 20031
rect 15680 19982 15750 19997
rect 16046 20067 16114 20084
rect 16046 20033 16063 20067
rect 16097 20033 16114 20067
rect 16046 19918 16114 20033
rect 16784 20031 16854 20232
rect 17569 20214 17581 20248
rect 17615 20214 17627 20248
rect 17754 20277 18823 20319
rect 17754 20243 17771 20277
rect 17805 20243 18771 20277
rect 18805 20243 18823 20277
rect 17754 20232 18823 20243
rect 18858 20277 19927 20319
rect 18858 20243 18875 20277
rect 18909 20243 19875 20277
rect 19909 20243 19927 20277
rect 18858 20232 19927 20243
rect 19961 20277 20203 20319
rect 19961 20243 19979 20277
rect 20013 20243 20151 20277
rect 20185 20243 20203 20277
rect 17569 20155 17627 20214
rect 17569 20121 17581 20155
rect 17615 20121 17627 20155
rect 17569 20086 17627 20121
rect 16784 19997 16803 20031
rect 16837 19997 16854 20031
rect 16784 19982 16854 19997
rect 17150 20067 17218 20084
rect 17150 20033 17167 20067
rect 17201 20033 17218 20067
rect 17150 19918 17218 20033
rect 18072 20031 18142 20232
rect 18072 19997 18091 20031
rect 18125 19997 18142 20031
rect 18072 19982 18142 19997
rect 18438 20067 18506 20084
rect 18438 20033 18455 20067
rect 18489 20033 18506 20067
rect 17569 19937 17627 19954
rect 12601 19870 12619 19904
rect 12653 19870 13067 19904
rect 13101 19870 13119 19904
rect 12601 19809 13119 19870
rect 13154 19904 14223 19918
rect 13154 19870 13171 19904
rect 13205 19870 14171 19904
rect 14205 19870 14223 19904
rect 13154 19809 14223 19870
rect 14258 19904 15327 19918
rect 14258 19870 14275 19904
rect 14309 19870 15275 19904
rect 15309 19870 15327 19904
rect 14258 19809 15327 19870
rect 15362 19904 16431 19918
rect 15362 19870 15379 19904
rect 15413 19870 16379 19904
rect 16413 19870 16431 19904
rect 15362 19809 16431 19870
rect 16466 19904 17535 19918
rect 16466 19870 16483 19904
rect 16517 19870 17483 19904
rect 17517 19870 17535 19904
rect 16466 19809 17535 19870
rect 17569 19903 17581 19937
rect 17615 19903 17627 19937
rect 18438 19918 18506 20033
rect 19176 20031 19246 20232
rect 19961 20182 20203 20243
rect 19961 20148 19979 20182
rect 20013 20148 20151 20182
rect 20185 20148 20203 20182
rect 19961 20101 20203 20148
rect 19176 19997 19195 20031
rect 19229 19997 19246 20031
rect 19176 19982 19246 19997
rect 19542 20067 19610 20084
rect 19542 20033 19559 20067
rect 19593 20033 19610 20067
rect 19542 19918 19610 20033
rect 19961 20027 20065 20101
rect 19961 19993 20011 20027
rect 20045 19993 20065 20027
rect 20099 20033 20119 20067
rect 20153 20033 20203 20067
rect 20099 19959 20203 20033
rect 17569 19809 17627 19903
rect 17754 19904 18823 19918
rect 17754 19870 17771 19904
rect 17805 19870 18771 19904
rect 18805 19870 18823 19904
rect 17754 19809 18823 19870
rect 18858 19904 19927 19918
rect 18858 19870 18875 19904
rect 18909 19870 19875 19904
rect 19909 19870 19927 19904
rect 18858 19809 19927 19870
rect 19961 19906 20203 19959
rect 19961 19872 19979 19906
rect 20013 19872 20151 19906
rect 20185 19872 20203 19906
rect 19961 19809 20203 19872
rect 4948 19775 4977 19809
rect 5011 19775 5069 19809
rect 5103 19775 5161 19809
rect 5195 19775 5253 19809
rect 5287 19775 5345 19809
rect 5379 19775 5437 19809
rect 5471 19775 5529 19809
rect 5563 19775 5621 19809
rect 5655 19775 5713 19809
rect 5747 19775 5805 19809
rect 5839 19775 5897 19809
rect 5931 19775 5989 19809
rect 6023 19775 6081 19809
rect 6115 19775 6173 19809
rect 6207 19775 6265 19809
rect 6299 19775 6357 19809
rect 6391 19775 6449 19809
rect 6483 19775 6541 19809
rect 6575 19775 6633 19809
rect 6667 19775 6725 19809
rect 6759 19775 6817 19809
rect 6851 19775 6909 19809
rect 6943 19775 7001 19809
rect 7035 19775 7093 19809
rect 7127 19775 7185 19809
rect 7219 19775 7277 19809
rect 7311 19775 7369 19809
rect 7403 19775 7461 19809
rect 7495 19775 7553 19809
rect 7587 19775 7645 19809
rect 7679 19775 7737 19809
rect 7771 19775 7829 19809
rect 7863 19775 7921 19809
rect 7955 19775 8013 19809
rect 8047 19775 8105 19809
rect 8139 19775 8197 19809
rect 8231 19775 8289 19809
rect 8323 19775 8381 19809
rect 8415 19775 8473 19809
rect 8507 19775 8565 19809
rect 8599 19775 8657 19809
rect 8691 19775 8749 19809
rect 8783 19775 8841 19809
rect 8875 19775 8933 19809
rect 8967 19775 9025 19809
rect 9059 19775 9117 19809
rect 9151 19775 9209 19809
rect 9243 19775 9301 19809
rect 9335 19775 9393 19809
rect 9427 19775 9485 19809
rect 9519 19775 9577 19809
rect 9611 19775 9669 19809
rect 9703 19775 9761 19809
rect 9795 19775 9853 19809
rect 9887 19775 9945 19809
rect 9979 19775 10037 19809
rect 10071 19775 10129 19809
rect 10163 19775 10221 19809
rect 10255 19775 10313 19809
rect 10347 19775 10405 19809
rect 10439 19775 10497 19809
rect 10531 19775 10589 19809
rect 10623 19775 10681 19809
rect 10715 19775 10773 19809
rect 10807 19775 10865 19809
rect 10899 19775 10957 19809
rect 10991 19775 11049 19809
rect 11083 19775 11141 19809
rect 11175 19775 11233 19809
rect 11267 19775 11325 19809
rect 11359 19775 11417 19809
rect 11451 19775 11509 19809
rect 11543 19775 11601 19809
rect 11635 19775 11693 19809
rect 11727 19775 11785 19809
rect 11819 19775 11877 19809
rect 11911 19775 11969 19809
rect 12003 19775 12061 19809
rect 12095 19775 12153 19809
rect 12187 19775 12245 19809
rect 12279 19775 12337 19809
rect 12371 19775 12429 19809
rect 12463 19775 12521 19809
rect 12555 19775 12613 19809
rect 12647 19775 12705 19809
rect 12739 19775 12797 19809
rect 12831 19775 12889 19809
rect 12923 19775 12981 19809
rect 13015 19775 13073 19809
rect 13107 19775 13165 19809
rect 13199 19775 13257 19809
rect 13291 19775 13349 19809
rect 13383 19775 13441 19809
rect 13475 19775 13533 19809
rect 13567 19775 13625 19809
rect 13659 19775 13717 19809
rect 13751 19775 13809 19809
rect 13843 19775 13901 19809
rect 13935 19775 13993 19809
rect 14027 19775 14085 19809
rect 14119 19775 14177 19809
rect 14211 19775 14269 19809
rect 14303 19775 14361 19809
rect 14395 19775 14453 19809
rect 14487 19775 14545 19809
rect 14579 19775 14637 19809
rect 14671 19775 14729 19809
rect 14763 19775 14821 19809
rect 14855 19775 14913 19809
rect 14947 19775 15005 19809
rect 15039 19775 15097 19809
rect 15131 19775 15189 19809
rect 15223 19775 15281 19809
rect 15315 19775 15373 19809
rect 15407 19775 15465 19809
rect 15499 19775 15557 19809
rect 15591 19775 15649 19809
rect 15683 19775 15741 19809
rect 15775 19775 15833 19809
rect 15867 19775 15925 19809
rect 15959 19775 16017 19809
rect 16051 19775 16109 19809
rect 16143 19775 16201 19809
rect 16235 19775 16293 19809
rect 16327 19775 16385 19809
rect 16419 19775 16477 19809
rect 16511 19775 16569 19809
rect 16603 19775 16661 19809
rect 16695 19775 16753 19809
rect 16787 19775 16845 19809
rect 16879 19775 16937 19809
rect 16971 19775 17029 19809
rect 17063 19775 17121 19809
rect 17155 19775 17213 19809
rect 17247 19775 17305 19809
rect 17339 19775 17397 19809
rect 17431 19775 17489 19809
rect 17523 19775 17581 19809
rect 17615 19775 17673 19809
rect 17707 19775 17765 19809
rect 17799 19775 17857 19809
rect 17891 19775 17949 19809
rect 17983 19775 18041 19809
rect 18075 19775 18133 19809
rect 18167 19775 18225 19809
rect 18259 19775 18317 19809
rect 18351 19775 18409 19809
rect 18443 19775 18501 19809
rect 18535 19775 18593 19809
rect 18627 19775 18685 19809
rect 18719 19775 18777 19809
rect 18811 19775 18869 19809
rect 18903 19775 18961 19809
rect 18995 19775 19053 19809
rect 19087 19775 19145 19809
rect 19179 19775 19237 19809
rect 19271 19775 19329 19809
rect 19363 19775 19421 19809
rect 19455 19775 19513 19809
rect 19547 19775 19605 19809
rect 19639 19775 19697 19809
rect 19731 19775 19789 19809
rect 19823 19775 19881 19809
rect 19915 19775 19973 19809
rect 20007 19775 20065 19809
rect 20099 19775 20157 19809
rect 20191 19775 20220 19809
rect 4965 19712 5207 19775
rect 4965 19678 4983 19712
rect 5017 19678 5155 19712
rect 5189 19678 5207 19712
rect 4965 19625 5207 19678
rect 5426 19714 6495 19775
rect 5426 19680 5443 19714
rect 5477 19680 6443 19714
rect 6477 19680 6495 19714
rect 5426 19666 6495 19680
rect 6530 19714 7599 19775
rect 6530 19680 6547 19714
rect 6581 19680 7547 19714
rect 7581 19680 7599 19714
rect 6530 19666 7599 19680
rect 7634 19714 8703 19775
rect 7634 19680 7651 19714
rect 7685 19680 8651 19714
rect 8685 19680 8703 19714
rect 7634 19666 8703 19680
rect 8738 19714 9807 19775
rect 8738 19680 8755 19714
rect 8789 19680 9755 19714
rect 9789 19680 9807 19714
rect 8738 19666 9807 19680
rect 9841 19681 9899 19775
rect 4965 19551 5069 19625
rect 4965 19517 5015 19551
rect 5049 19517 5069 19551
rect 5103 19557 5123 19591
rect 5157 19557 5207 19591
rect 5103 19483 5207 19557
rect 4965 19436 5207 19483
rect 4965 19402 4983 19436
rect 5017 19402 5155 19436
rect 5189 19402 5207 19436
rect 4965 19341 5207 19402
rect 5744 19587 5814 19602
rect 5744 19553 5763 19587
rect 5797 19553 5814 19587
rect 5744 19352 5814 19553
rect 6110 19551 6178 19666
rect 6110 19517 6127 19551
rect 6161 19517 6178 19551
rect 6110 19500 6178 19517
rect 6848 19587 6918 19602
rect 6848 19553 6867 19587
rect 6901 19553 6918 19587
rect 6848 19352 6918 19553
rect 7214 19551 7282 19666
rect 7214 19517 7231 19551
rect 7265 19517 7282 19551
rect 7214 19500 7282 19517
rect 7952 19587 8022 19602
rect 7952 19553 7971 19587
rect 8005 19553 8022 19587
rect 7952 19352 8022 19553
rect 8318 19551 8386 19666
rect 8318 19517 8335 19551
rect 8369 19517 8386 19551
rect 8318 19500 8386 19517
rect 9056 19587 9126 19602
rect 9056 19553 9075 19587
rect 9109 19553 9126 19587
rect 9056 19352 9126 19553
rect 9422 19551 9490 19666
rect 9841 19647 9853 19681
rect 9887 19647 9899 19681
rect 9841 19630 9899 19647
rect 10025 19714 10543 19775
rect 10025 19680 10043 19714
rect 10077 19680 10491 19714
rect 10525 19680 10543 19714
rect 10025 19621 10543 19680
rect 10578 19714 11647 19775
rect 10578 19680 10595 19714
rect 10629 19680 11595 19714
rect 11629 19680 11647 19714
rect 10578 19666 11647 19680
rect 11682 19714 12751 19775
rect 11682 19680 11699 19714
rect 11733 19680 12699 19714
rect 12733 19680 12751 19714
rect 11682 19666 12751 19680
rect 12786 19714 13855 19775
rect 12786 19680 12803 19714
rect 12837 19680 13803 19714
rect 13837 19680 13855 19714
rect 12786 19666 13855 19680
rect 13890 19714 14959 19775
rect 13890 19680 13907 19714
rect 13941 19680 14907 19714
rect 14941 19680 14959 19714
rect 13890 19666 14959 19680
rect 14993 19681 15051 19775
rect 9422 19517 9439 19551
rect 9473 19517 9490 19551
rect 9422 19500 9490 19517
rect 10025 19553 10103 19587
rect 10137 19553 10213 19587
rect 10247 19553 10267 19587
rect 9841 19463 9899 19498
rect 9841 19429 9853 19463
rect 9887 19429 9899 19463
rect 9841 19370 9899 19429
rect 4965 19307 4983 19341
rect 5017 19307 5155 19341
rect 5189 19307 5207 19341
rect 4965 19265 5207 19307
rect 5426 19341 6495 19352
rect 5426 19307 5443 19341
rect 5477 19307 6443 19341
rect 6477 19307 6495 19341
rect 5426 19265 6495 19307
rect 6530 19341 7599 19352
rect 6530 19307 6547 19341
rect 6581 19307 7547 19341
rect 7581 19307 7599 19341
rect 6530 19265 7599 19307
rect 7634 19341 8703 19352
rect 7634 19307 7651 19341
rect 7685 19307 8651 19341
rect 8685 19307 8703 19341
rect 7634 19265 8703 19307
rect 8738 19341 9807 19352
rect 8738 19307 8755 19341
rect 8789 19307 9755 19341
rect 9789 19307 9807 19341
rect 8738 19265 9807 19307
rect 9841 19336 9853 19370
rect 9887 19336 9899 19370
rect 9841 19265 9899 19336
rect 10025 19483 10267 19553
rect 10301 19551 10543 19621
rect 10301 19517 10321 19551
rect 10355 19517 10431 19551
rect 10465 19517 10543 19551
rect 10896 19587 10966 19602
rect 10896 19553 10915 19587
rect 10949 19553 10966 19587
rect 10025 19443 10543 19483
rect 10025 19409 10043 19443
rect 10077 19409 10491 19443
rect 10525 19409 10543 19443
rect 10025 19341 10543 19409
rect 10896 19352 10966 19553
rect 11262 19551 11330 19666
rect 11262 19517 11279 19551
rect 11313 19517 11330 19551
rect 11262 19500 11330 19517
rect 12000 19587 12070 19602
rect 12000 19553 12019 19587
rect 12053 19553 12070 19587
rect 12000 19352 12070 19553
rect 12366 19551 12434 19666
rect 12366 19517 12383 19551
rect 12417 19517 12434 19551
rect 12366 19500 12434 19517
rect 13104 19587 13174 19602
rect 13104 19553 13123 19587
rect 13157 19553 13174 19587
rect 13104 19352 13174 19553
rect 13470 19551 13538 19666
rect 13470 19517 13487 19551
rect 13521 19517 13538 19551
rect 13470 19500 13538 19517
rect 14208 19587 14278 19602
rect 14208 19553 14227 19587
rect 14261 19553 14278 19587
rect 14208 19352 14278 19553
rect 14574 19551 14642 19666
rect 14993 19647 15005 19681
rect 15039 19647 15051 19681
rect 14993 19630 15051 19647
rect 15177 19707 15511 19775
rect 15177 19673 15195 19707
rect 15229 19673 15459 19707
rect 15493 19673 15511 19707
rect 15177 19621 15511 19673
rect 15546 19714 16615 19775
rect 15546 19680 15563 19714
rect 15597 19680 16563 19714
rect 16597 19680 16615 19714
rect 15546 19666 16615 19680
rect 16650 19714 17719 19775
rect 16650 19680 16667 19714
rect 16701 19680 17667 19714
rect 17701 19680 17719 19714
rect 16650 19666 17719 19680
rect 17754 19714 18823 19775
rect 17754 19680 17771 19714
rect 17805 19680 18771 19714
rect 18805 19680 18823 19714
rect 17754 19666 18823 19680
rect 18858 19714 19927 19775
rect 18858 19680 18875 19714
rect 18909 19680 19875 19714
rect 19909 19680 19927 19714
rect 18858 19666 19927 19680
rect 19961 19712 20203 19775
rect 19961 19678 19979 19712
rect 20013 19678 20151 19712
rect 20185 19678 20203 19712
rect 14574 19517 14591 19551
rect 14625 19517 14642 19551
rect 14574 19500 14642 19517
rect 15177 19553 15197 19587
rect 15231 19553 15327 19587
rect 14993 19463 15051 19498
rect 14993 19429 15005 19463
rect 15039 19429 15051 19463
rect 14993 19370 15051 19429
rect 10025 19307 10043 19341
rect 10077 19307 10491 19341
rect 10525 19307 10543 19341
rect 10025 19265 10543 19307
rect 10578 19341 11647 19352
rect 10578 19307 10595 19341
rect 10629 19307 11595 19341
rect 11629 19307 11647 19341
rect 10578 19265 11647 19307
rect 11682 19341 12751 19352
rect 11682 19307 11699 19341
rect 11733 19307 12699 19341
rect 12733 19307 12751 19341
rect 11682 19265 12751 19307
rect 12786 19341 13855 19352
rect 12786 19307 12803 19341
rect 12837 19307 13803 19341
rect 13837 19307 13855 19341
rect 12786 19265 13855 19307
rect 13890 19341 14959 19352
rect 13890 19307 13907 19341
rect 13941 19307 14907 19341
rect 14941 19307 14959 19341
rect 13890 19265 14959 19307
rect 14993 19336 15005 19370
rect 15039 19336 15051 19370
rect 14993 19265 15051 19336
rect 15177 19483 15327 19553
rect 15361 19551 15511 19621
rect 15361 19517 15457 19551
rect 15491 19517 15511 19551
rect 15864 19587 15934 19602
rect 15864 19553 15883 19587
rect 15917 19553 15934 19587
rect 15177 19443 15511 19483
rect 15177 19409 15195 19443
rect 15229 19409 15459 19443
rect 15493 19409 15511 19443
rect 15177 19341 15511 19409
rect 15864 19352 15934 19553
rect 16230 19551 16298 19666
rect 16230 19517 16247 19551
rect 16281 19517 16298 19551
rect 16230 19500 16298 19517
rect 16968 19587 17038 19602
rect 16968 19553 16987 19587
rect 17021 19553 17038 19587
rect 16968 19352 17038 19553
rect 17334 19551 17402 19666
rect 17334 19517 17351 19551
rect 17385 19517 17402 19551
rect 17334 19500 17402 19517
rect 18072 19587 18142 19602
rect 18072 19553 18091 19587
rect 18125 19553 18142 19587
rect 18072 19352 18142 19553
rect 18438 19551 18506 19666
rect 18438 19517 18455 19551
rect 18489 19517 18506 19551
rect 18438 19500 18506 19517
rect 19176 19587 19246 19602
rect 19176 19553 19195 19587
rect 19229 19553 19246 19587
rect 19176 19352 19246 19553
rect 19542 19551 19610 19666
rect 19961 19625 20203 19678
rect 19542 19517 19559 19551
rect 19593 19517 19610 19551
rect 19542 19500 19610 19517
rect 19961 19557 20011 19591
rect 20045 19557 20065 19591
rect 19961 19483 20065 19557
rect 20099 19551 20203 19625
rect 20099 19517 20119 19551
rect 20153 19517 20203 19551
rect 19961 19436 20203 19483
rect 19961 19402 19979 19436
rect 20013 19402 20151 19436
rect 20185 19402 20203 19436
rect 15177 19307 15195 19341
rect 15229 19307 15459 19341
rect 15493 19307 15511 19341
rect 15177 19265 15511 19307
rect 15546 19341 16615 19352
rect 15546 19307 15563 19341
rect 15597 19307 16563 19341
rect 16597 19307 16615 19341
rect 15546 19265 16615 19307
rect 16650 19341 17719 19352
rect 16650 19307 16667 19341
rect 16701 19307 17667 19341
rect 17701 19307 17719 19341
rect 16650 19265 17719 19307
rect 17754 19341 18823 19352
rect 17754 19307 17771 19341
rect 17805 19307 18771 19341
rect 18805 19307 18823 19341
rect 17754 19265 18823 19307
rect 18858 19341 19927 19352
rect 18858 19307 18875 19341
rect 18909 19307 19875 19341
rect 19909 19307 19927 19341
rect 18858 19265 19927 19307
rect 19961 19341 20203 19402
rect 19961 19307 19979 19341
rect 20013 19307 20151 19341
rect 20185 19307 20203 19341
rect 19961 19265 20203 19307
rect 4948 19231 4977 19265
rect 5011 19231 5069 19265
rect 5103 19231 5161 19265
rect 5195 19231 5253 19265
rect 5287 19231 5345 19265
rect 5379 19231 5437 19265
rect 5471 19231 5529 19265
rect 5563 19231 5621 19265
rect 5655 19231 5713 19265
rect 5747 19231 5805 19265
rect 5839 19231 5897 19265
rect 5931 19231 5989 19265
rect 6023 19231 6081 19265
rect 6115 19231 6173 19265
rect 6207 19231 6265 19265
rect 6299 19231 6357 19265
rect 6391 19231 6449 19265
rect 6483 19231 6541 19265
rect 6575 19231 6633 19265
rect 6667 19231 6725 19265
rect 6759 19231 6817 19265
rect 6851 19231 6909 19265
rect 6943 19231 7001 19265
rect 7035 19231 7093 19265
rect 7127 19231 7185 19265
rect 7219 19231 7277 19265
rect 7311 19231 7369 19265
rect 7403 19231 7461 19265
rect 7495 19231 7553 19265
rect 7587 19231 7645 19265
rect 7679 19231 7737 19265
rect 7771 19231 7829 19265
rect 7863 19231 7921 19265
rect 7955 19231 8013 19265
rect 8047 19231 8105 19265
rect 8139 19231 8197 19265
rect 8231 19231 8289 19265
rect 8323 19231 8381 19265
rect 8415 19231 8473 19265
rect 8507 19231 8565 19265
rect 8599 19231 8657 19265
rect 8691 19231 8749 19265
rect 8783 19231 8841 19265
rect 8875 19231 8933 19265
rect 8967 19231 9025 19265
rect 9059 19231 9117 19265
rect 9151 19231 9209 19265
rect 9243 19231 9301 19265
rect 9335 19231 9393 19265
rect 9427 19231 9485 19265
rect 9519 19231 9577 19265
rect 9611 19231 9669 19265
rect 9703 19231 9761 19265
rect 9795 19231 9853 19265
rect 9887 19231 9945 19265
rect 9979 19231 10037 19265
rect 10071 19231 10129 19265
rect 10163 19231 10221 19265
rect 10255 19231 10313 19265
rect 10347 19231 10405 19265
rect 10439 19231 10497 19265
rect 10531 19231 10589 19265
rect 10623 19231 10681 19265
rect 10715 19231 10773 19265
rect 10807 19231 10865 19265
rect 10899 19231 10957 19265
rect 10991 19231 11049 19265
rect 11083 19231 11141 19265
rect 11175 19231 11233 19265
rect 11267 19231 11325 19265
rect 11359 19231 11417 19265
rect 11451 19231 11509 19265
rect 11543 19231 11601 19265
rect 11635 19231 11693 19265
rect 11727 19231 11785 19265
rect 11819 19231 11877 19265
rect 11911 19231 11969 19265
rect 12003 19231 12061 19265
rect 12095 19231 12153 19265
rect 12187 19231 12245 19265
rect 12279 19231 12337 19265
rect 12371 19231 12429 19265
rect 12463 19231 12521 19265
rect 12555 19231 12613 19265
rect 12647 19231 12705 19265
rect 12739 19231 12797 19265
rect 12831 19231 12889 19265
rect 12923 19231 12981 19265
rect 13015 19231 13073 19265
rect 13107 19231 13165 19265
rect 13199 19231 13257 19265
rect 13291 19231 13349 19265
rect 13383 19231 13441 19265
rect 13475 19231 13533 19265
rect 13567 19231 13625 19265
rect 13659 19231 13717 19265
rect 13751 19231 13809 19265
rect 13843 19231 13901 19265
rect 13935 19231 13993 19265
rect 14027 19231 14085 19265
rect 14119 19231 14177 19265
rect 14211 19231 14269 19265
rect 14303 19231 14361 19265
rect 14395 19231 14453 19265
rect 14487 19231 14545 19265
rect 14579 19231 14637 19265
rect 14671 19231 14729 19265
rect 14763 19231 14821 19265
rect 14855 19231 14913 19265
rect 14947 19231 15005 19265
rect 15039 19231 15097 19265
rect 15131 19231 15189 19265
rect 15223 19231 15281 19265
rect 15315 19231 15373 19265
rect 15407 19231 15465 19265
rect 15499 19231 15557 19265
rect 15591 19231 15649 19265
rect 15683 19231 15741 19265
rect 15775 19231 15833 19265
rect 15867 19231 15925 19265
rect 15959 19231 16017 19265
rect 16051 19231 16109 19265
rect 16143 19231 16201 19265
rect 16235 19231 16293 19265
rect 16327 19231 16385 19265
rect 16419 19231 16477 19265
rect 16511 19231 16569 19265
rect 16603 19231 16661 19265
rect 16695 19231 16753 19265
rect 16787 19231 16845 19265
rect 16879 19231 16937 19265
rect 16971 19231 17029 19265
rect 17063 19231 17121 19265
rect 17155 19231 17213 19265
rect 17247 19231 17305 19265
rect 17339 19231 17397 19265
rect 17431 19231 17489 19265
rect 17523 19231 17581 19265
rect 17615 19231 17673 19265
rect 17707 19231 17765 19265
rect 17799 19231 17857 19265
rect 17891 19231 17949 19265
rect 17983 19231 18041 19265
rect 18075 19231 18133 19265
rect 18167 19231 18225 19265
rect 18259 19231 18317 19265
rect 18351 19231 18409 19265
rect 18443 19231 18501 19265
rect 18535 19231 18593 19265
rect 18627 19231 18685 19265
rect 18719 19231 18777 19265
rect 18811 19231 18869 19265
rect 18903 19231 18961 19265
rect 18995 19231 19053 19265
rect 19087 19231 19145 19265
rect 19179 19231 19237 19265
rect 19271 19231 19329 19265
rect 19363 19231 19421 19265
rect 19455 19231 19513 19265
rect 19547 19231 19605 19265
rect 19639 19231 19697 19265
rect 19731 19231 19789 19265
rect 19823 19231 19881 19265
rect 19915 19231 19973 19265
rect 20007 19231 20065 19265
rect 20099 19231 20157 19265
rect 20191 19231 20220 19265
rect 4965 19189 5207 19231
rect 4965 19155 4983 19189
rect 5017 19155 5155 19189
rect 5189 19155 5207 19189
rect 4965 19094 5207 19155
rect 4965 19060 4983 19094
rect 5017 19060 5155 19094
rect 5189 19060 5207 19094
rect 4965 19013 5207 19060
rect 4965 18945 5015 18979
rect 5049 18945 5069 18979
rect 4965 18871 5069 18945
rect 5103 18939 5207 19013
rect 5103 18905 5123 18939
rect 5157 18905 5207 18939
rect 5425 19189 6127 19231
rect 5425 19155 5443 19189
rect 5477 19155 6075 19189
rect 6109 19155 6127 19189
rect 5425 19087 6127 19155
rect 6162 19189 7231 19231
rect 6162 19155 6179 19189
rect 6213 19155 7179 19189
rect 7213 19155 7231 19189
rect 6162 19144 7231 19155
rect 7265 19160 7323 19231
rect 5425 19053 5443 19087
rect 5477 19053 6075 19087
rect 6109 19053 6127 19087
rect 5425 19013 6127 19053
rect 5425 18943 5763 19013
rect 5425 18909 5503 18943
rect 5537 18909 5606 18943
rect 5640 18909 5709 18943
rect 5743 18909 5763 18943
rect 5797 18945 5817 18979
rect 5851 18945 5916 18979
rect 5950 18945 6015 18979
rect 6049 18945 6127 18979
rect 5797 18875 6127 18945
rect 6480 18943 6550 19144
rect 7265 19126 7277 19160
rect 7311 19126 7323 19160
rect 7265 19067 7323 19126
rect 7265 19033 7277 19067
rect 7311 19033 7323 19067
rect 7265 18998 7323 19033
rect 7449 19189 7967 19231
rect 7449 19155 7467 19189
rect 7501 19155 7915 19189
rect 7949 19155 7967 19189
rect 7449 19087 7967 19155
rect 8002 19189 9071 19231
rect 8002 19155 8019 19189
rect 8053 19155 9019 19189
rect 9053 19155 9071 19189
rect 8002 19144 9071 19155
rect 9106 19189 10175 19231
rect 9106 19155 9123 19189
rect 9157 19155 10123 19189
rect 10157 19155 10175 19189
rect 9106 19144 10175 19155
rect 10210 19189 11279 19231
rect 10210 19155 10227 19189
rect 10261 19155 11227 19189
rect 11261 19155 11279 19189
rect 10210 19144 11279 19155
rect 11314 19189 12383 19231
rect 11314 19155 11331 19189
rect 11365 19155 12331 19189
rect 12365 19155 12383 19189
rect 11314 19144 12383 19155
rect 12417 19160 12475 19231
rect 7449 19053 7467 19087
rect 7501 19053 7915 19087
rect 7949 19053 7967 19087
rect 7449 19013 7967 19053
rect 6480 18909 6499 18943
rect 6533 18909 6550 18943
rect 6480 18894 6550 18909
rect 6846 18979 6914 18996
rect 6846 18945 6863 18979
rect 6897 18945 6914 18979
rect 4965 18818 5207 18871
rect 4965 18784 4983 18818
rect 5017 18784 5155 18818
rect 5189 18784 5207 18818
rect 4965 18721 5207 18784
rect 5425 18816 6127 18875
rect 6846 18830 6914 18945
rect 7449 18943 7691 19013
rect 7449 18909 7527 18943
rect 7561 18909 7637 18943
rect 7671 18909 7691 18943
rect 7725 18945 7745 18979
rect 7779 18945 7855 18979
rect 7889 18945 7967 18979
rect 7725 18875 7967 18945
rect 8320 18943 8390 19144
rect 8320 18909 8339 18943
rect 8373 18909 8390 18943
rect 8320 18894 8390 18909
rect 8686 18979 8754 18996
rect 8686 18945 8703 18979
rect 8737 18945 8754 18979
rect 7265 18849 7323 18866
rect 5425 18782 5443 18816
rect 5477 18782 6075 18816
rect 6109 18782 6127 18816
rect 5425 18721 6127 18782
rect 6162 18816 7231 18830
rect 6162 18782 6179 18816
rect 6213 18782 7179 18816
rect 7213 18782 7231 18816
rect 6162 18721 7231 18782
rect 7265 18815 7277 18849
rect 7311 18815 7323 18849
rect 7265 18721 7323 18815
rect 7449 18816 7967 18875
rect 8686 18830 8754 18945
rect 9424 18943 9494 19144
rect 9424 18909 9443 18943
rect 9477 18909 9494 18943
rect 9424 18894 9494 18909
rect 9790 18979 9858 18996
rect 9790 18945 9807 18979
rect 9841 18945 9858 18979
rect 9790 18830 9858 18945
rect 10528 18943 10598 19144
rect 10528 18909 10547 18943
rect 10581 18909 10598 18943
rect 10528 18894 10598 18909
rect 10894 18979 10962 18996
rect 10894 18945 10911 18979
rect 10945 18945 10962 18979
rect 10894 18830 10962 18945
rect 11632 18943 11702 19144
rect 12417 19126 12429 19160
rect 12463 19126 12475 19160
rect 12417 19067 12475 19126
rect 12417 19033 12429 19067
rect 12463 19033 12475 19067
rect 12417 18998 12475 19033
rect 12601 19189 13119 19231
rect 12601 19155 12619 19189
rect 12653 19155 13067 19189
rect 13101 19155 13119 19189
rect 12601 19087 13119 19155
rect 13154 19189 14223 19231
rect 13154 19155 13171 19189
rect 13205 19155 14171 19189
rect 14205 19155 14223 19189
rect 13154 19144 14223 19155
rect 14258 19189 15327 19231
rect 14258 19155 14275 19189
rect 14309 19155 15275 19189
rect 15309 19155 15327 19189
rect 14258 19144 15327 19155
rect 15362 19189 16431 19231
rect 15362 19155 15379 19189
rect 15413 19155 16379 19189
rect 16413 19155 16431 19189
rect 15362 19144 16431 19155
rect 16466 19189 17535 19231
rect 16466 19155 16483 19189
rect 16517 19155 17483 19189
rect 17517 19155 17535 19189
rect 16466 19144 17535 19155
rect 17569 19160 17627 19231
rect 12601 19053 12619 19087
rect 12653 19053 13067 19087
rect 13101 19053 13119 19087
rect 12601 19013 13119 19053
rect 11632 18909 11651 18943
rect 11685 18909 11702 18943
rect 11632 18894 11702 18909
rect 11998 18979 12066 18996
rect 11998 18945 12015 18979
rect 12049 18945 12066 18979
rect 11998 18830 12066 18945
rect 12601 18943 12843 19013
rect 12601 18909 12679 18943
rect 12713 18909 12789 18943
rect 12823 18909 12843 18943
rect 12877 18945 12897 18979
rect 12931 18945 13007 18979
rect 13041 18945 13119 18979
rect 12877 18875 13119 18945
rect 13472 18943 13542 19144
rect 13472 18909 13491 18943
rect 13525 18909 13542 18943
rect 13472 18894 13542 18909
rect 13838 18979 13906 18996
rect 13838 18945 13855 18979
rect 13889 18945 13906 18979
rect 12417 18849 12475 18866
rect 7449 18782 7467 18816
rect 7501 18782 7915 18816
rect 7949 18782 7967 18816
rect 7449 18721 7967 18782
rect 8002 18816 9071 18830
rect 8002 18782 8019 18816
rect 8053 18782 9019 18816
rect 9053 18782 9071 18816
rect 8002 18721 9071 18782
rect 9106 18816 10175 18830
rect 9106 18782 9123 18816
rect 9157 18782 10123 18816
rect 10157 18782 10175 18816
rect 9106 18721 10175 18782
rect 10210 18816 11279 18830
rect 10210 18782 10227 18816
rect 10261 18782 11227 18816
rect 11261 18782 11279 18816
rect 10210 18721 11279 18782
rect 11314 18816 12383 18830
rect 11314 18782 11331 18816
rect 11365 18782 12331 18816
rect 12365 18782 12383 18816
rect 11314 18721 12383 18782
rect 12417 18815 12429 18849
rect 12463 18815 12475 18849
rect 12417 18721 12475 18815
rect 12601 18816 13119 18875
rect 13838 18830 13906 18945
rect 14576 18943 14646 19144
rect 14576 18909 14595 18943
rect 14629 18909 14646 18943
rect 14576 18894 14646 18909
rect 14942 18979 15010 18996
rect 14942 18945 14959 18979
rect 14993 18945 15010 18979
rect 14942 18830 15010 18945
rect 15680 18943 15750 19144
rect 15680 18909 15699 18943
rect 15733 18909 15750 18943
rect 15680 18894 15750 18909
rect 16046 18979 16114 18996
rect 16046 18945 16063 18979
rect 16097 18945 16114 18979
rect 16046 18830 16114 18945
rect 16784 18943 16854 19144
rect 17569 19126 17581 19160
rect 17615 19126 17627 19160
rect 17754 19189 18823 19231
rect 17754 19155 17771 19189
rect 17805 19155 18771 19189
rect 18805 19155 18823 19189
rect 17754 19144 18823 19155
rect 18858 19189 19927 19231
rect 18858 19155 18875 19189
rect 18909 19155 19875 19189
rect 19909 19155 19927 19189
rect 18858 19144 19927 19155
rect 19961 19189 20203 19231
rect 19961 19155 19979 19189
rect 20013 19155 20151 19189
rect 20185 19155 20203 19189
rect 17569 19067 17627 19126
rect 17569 19033 17581 19067
rect 17615 19033 17627 19067
rect 17569 18998 17627 19033
rect 16784 18909 16803 18943
rect 16837 18909 16854 18943
rect 16784 18894 16854 18909
rect 17150 18979 17218 18996
rect 17150 18945 17167 18979
rect 17201 18945 17218 18979
rect 17150 18830 17218 18945
rect 18072 18943 18142 19144
rect 18072 18909 18091 18943
rect 18125 18909 18142 18943
rect 18072 18894 18142 18909
rect 18438 18979 18506 18996
rect 18438 18945 18455 18979
rect 18489 18945 18506 18979
rect 17569 18849 17627 18866
rect 12601 18782 12619 18816
rect 12653 18782 13067 18816
rect 13101 18782 13119 18816
rect 12601 18721 13119 18782
rect 13154 18816 14223 18830
rect 13154 18782 13171 18816
rect 13205 18782 14171 18816
rect 14205 18782 14223 18816
rect 13154 18721 14223 18782
rect 14258 18816 15327 18830
rect 14258 18782 14275 18816
rect 14309 18782 15275 18816
rect 15309 18782 15327 18816
rect 14258 18721 15327 18782
rect 15362 18816 16431 18830
rect 15362 18782 15379 18816
rect 15413 18782 16379 18816
rect 16413 18782 16431 18816
rect 15362 18721 16431 18782
rect 16466 18816 17535 18830
rect 16466 18782 16483 18816
rect 16517 18782 17483 18816
rect 17517 18782 17535 18816
rect 16466 18721 17535 18782
rect 17569 18815 17581 18849
rect 17615 18815 17627 18849
rect 18438 18830 18506 18945
rect 19176 18943 19246 19144
rect 19961 19094 20203 19155
rect 19961 19060 19979 19094
rect 20013 19060 20151 19094
rect 20185 19060 20203 19094
rect 19961 19013 20203 19060
rect 19176 18909 19195 18943
rect 19229 18909 19246 18943
rect 19176 18894 19246 18909
rect 19542 18979 19610 18996
rect 19542 18945 19559 18979
rect 19593 18945 19610 18979
rect 19542 18830 19610 18945
rect 19961 18939 20065 19013
rect 19961 18905 20011 18939
rect 20045 18905 20065 18939
rect 20099 18945 20119 18979
rect 20153 18945 20203 18979
rect 20099 18871 20203 18945
rect 17569 18721 17627 18815
rect 17754 18816 18823 18830
rect 17754 18782 17771 18816
rect 17805 18782 18771 18816
rect 18805 18782 18823 18816
rect 17754 18721 18823 18782
rect 18858 18816 19927 18830
rect 18858 18782 18875 18816
rect 18909 18782 19875 18816
rect 19909 18782 19927 18816
rect 18858 18721 19927 18782
rect 19961 18818 20203 18871
rect 19961 18784 19979 18818
rect 20013 18784 20151 18818
rect 20185 18784 20203 18818
rect 19961 18721 20203 18784
rect 4948 18687 4977 18721
rect 5011 18687 5069 18721
rect 5103 18687 5161 18721
rect 5195 18687 5253 18721
rect 5287 18687 5345 18721
rect 5379 18687 5437 18721
rect 5471 18687 5529 18721
rect 5563 18687 5621 18721
rect 5655 18687 5713 18721
rect 5747 18687 5805 18721
rect 5839 18687 5897 18721
rect 5931 18687 5989 18721
rect 6023 18687 6081 18721
rect 6115 18687 6173 18721
rect 6207 18687 6265 18721
rect 6299 18687 6357 18721
rect 6391 18687 6449 18721
rect 6483 18687 6541 18721
rect 6575 18687 6633 18721
rect 6667 18687 6725 18721
rect 6759 18687 6817 18721
rect 6851 18687 6909 18721
rect 6943 18687 7001 18721
rect 7035 18687 7093 18721
rect 7127 18687 7185 18721
rect 7219 18687 7277 18721
rect 7311 18687 7369 18721
rect 7403 18687 7461 18721
rect 7495 18687 7553 18721
rect 7587 18687 7645 18721
rect 7679 18687 7737 18721
rect 7771 18687 7829 18721
rect 7863 18687 7921 18721
rect 7955 18687 8013 18721
rect 8047 18687 8105 18721
rect 8139 18687 8197 18721
rect 8231 18687 8289 18721
rect 8323 18687 8381 18721
rect 8415 18687 8473 18721
rect 8507 18687 8565 18721
rect 8599 18687 8657 18721
rect 8691 18687 8749 18721
rect 8783 18687 8841 18721
rect 8875 18687 8933 18721
rect 8967 18687 9025 18721
rect 9059 18687 9117 18721
rect 9151 18687 9209 18721
rect 9243 18687 9301 18721
rect 9335 18687 9393 18721
rect 9427 18687 9485 18721
rect 9519 18687 9577 18721
rect 9611 18687 9669 18721
rect 9703 18687 9761 18721
rect 9795 18687 9853 18721
rect 9887 18687 9945 18721
rect 9979 18687 10037 18721
rect 10071 18687 10129 18721
rect 10163 18687 10221 18721
rect 10255 18687 10313 18721
rect 10347 18687 10405 18721
rect 10439 18687 10497 18721
rect 10531 18687 10589 18721
rect 10623 18687 10681 18721
rect 10715 18687 10773 18721
rect 10807 18687 10865 18721
rect 10899 18687 10957 18721
rect 10991 18687 11049 18721
rect 11083 18687 11141 18721
rect 11175 18687 11233 18721
rect 11267 18687 11325 18721
rect 11359 18687 11417 18721
rect 11451 18687 11509 18721
rect 11543 18687 11601 18721
rect 11635 18687 11693 18721
rect 11727 18687 11785 18721
rect 11819 18687 11877 18721
rect 11911 18687 11969 18721
rect 12003 18687 12061 18721
rect 12095 18687 12153 18721
rect 12187 18687 12245 18721
rect 12279 18687 12337 18721
rect 12371 18687 12429 18721
rect 12463 18687 12521 18721
rect 12555 18687 12613 18721
rect 12647 18687 12705 18721
rect 12739 18687 12797 18721
rect 12831 18687 12889 18721
rect 12923 18687 12981 18721
rect 13015 18687 13073 18721
rect 13107 18687 13165 18721
rect 13199 18687 13257 18721
rect 13291 18687 13349 18721
rect 13383 18687 13441 18721
rect 13475 18687 13533 18721
rect 13567 18687 13625 18721
rect 13659 18687 13717 18721
rect 13751 18687 13809 18721
rect 13843 18687 13901 18721
rect 13935 18687 13993 18721
rect 14027 18687 14085 18721
rect 14119 18687 14177 18721
rect 14211 18687 14269 18721
rect 14303 18687 14361 18721
rect 14395 18687 14453 18721
rect 14487 18687 14545 18721
rect 14579 18687 14637 18721
rect 14671 18687 14729 18721
rect 14763 18687 14821 18721
rect 14855 18687 14913 18721
rect 14947 18687 15005 18721
rect 15039 18687 15097 18721
rect 15131 18687 15189 18721
rect 15223 18687 15281 18721
rect 15315 18687 15373 18721
rect 15407 18687 15465 18721
rect 15499 18687 15557 18721
rect 15591 18687 15649 18721
rect 15683 18687 15741 18721
rect 15775 18687 15833 18721
rect 15867 18687 15925 18721
rect 15959 18687 16017 18721
rect 16051 18687 16109 18721
rect 16143 18687 16201 18721
rect 16235 18687 16293 18721
rect 16327 18687 16385 18721
rect 16419 18687 16477 18721
rect 16511 18687 16569 18721
rect 16603 18687 16661 18721
rect 16695 18687 16753 18721
rect 16787 18687 16845 18721
rect 16879 18687 16937 18721
rect 16971 18687 17029 18721
rect 17063 18687 17121 18721
rect 17155 18687 17213 18721
rect 17247 18687 17305 18721
rect 17339 18687 17397 18721
rect 17431 18687 17489 18721
rect 17523 18687 17581 18721
rect 17615 18687 17673 18721
rect 17707 18687 17765 18721
rect 17799 18687 17857 18721
rect 17891 18687 17949 18721
rect 17983 18687 18041 18721
rect 18075 18687 18133 18721
rect 18167 18687 18225 18721
rect 18259 18687 18317 18721
rect 18351 18687 18409 18721
rect 18443 18687 18501 18721
rect 18535 18687 18593 18721
rect 18627 18687 18685 18721
rect 18719 18687 18777 18721
rect 18811 18687 18869 18721
rect 18903 18687 18961 18721
rect 18995 18687 19053 18721
rect 19087 18687 19145 18721
rect 19179 18687 19237 18721
rect 19271 18687 19329 18721
rect 19363 18687 19421 18721
rect 19455 18687 19513 18721
rect 19547 18687 19605 18721
rect 19639 18687 19697 18721
rect 19731 18687 19789 18721
rect 19823 18687 19881 18721
rect 19915 18687 19973 18721
rect 20007 18687 20065 18721
rect 20099 18687 20157 18721
rect 20191 18687 20220 18721
rect 4965 18624 5207 18687
rect 4965 18590 4983 18624
rect 5017 18590 5155 18624
rect 5189 18590 5207 18624
rect 4965 18537 5207 18590
rect 5426 18626 6495 18687
rect 5426 18592 5443 18626
rect 5477 18592 6443 18626
rect 6477 18592 6495 18626
rect 5426 18578 6495 18592
rect 6530 18626 7599 18687
rect 6530 18592 6547 18626
rect 6581 18592 7547 18626
rect 7581 18592 7599 18626
rect 6530 18578 7599 18592
rect 7634 18626 8703 18687
rect 7634 18592 7651 18626
rect 7685 18592 8651 18626
rect 8685 18592 8703 18626
rect 7634 18578 8703 18592
rect 8738 18626 9807 18687
rect 8738 18592 8755 18626
rect 8789 18592 9755 18626
rect 9789 18592 9807 18626
rect 8738 18578 9807 18592
rect 9841 18593 9899 18687
rect 4965 18463 5069 18537
rect 4965 18429 5015 18463
rect 5049 18429 5069 18463
rect 5103 18469 5123 18503
rect 5157 18469 5207 18503
rect 5103 18395 5207 18469
rect 4965 18348 5207 18395
rect 4965 18314 4983 18348
rect 5017 18314 5155 18348
rect 5189 18314 5207 18348
rect 4965 18253 5207 18314
rect 5744 18499 5814 18514
rect 5744 18465 5763 18499
rect 5797 18465 5814 18499
rect 5744 18264 5814 18465
rect 6110 18463 6178 18578
rect 6110 18429 6127 18463
rect 6161 18429 6178 18463
rect 6110 18412 6178 18429
rect 6848 18499 6918 18514
rect 6848 18465 6867 18499
rect 6901 18465 6918 18499
rect 6848 18264 6918 18465
rect 7214 18463 7282 18578
rect 7214 18429 7231 18463
rect 7265 18429 7282 18463
rect 7214 18412 7282 18429
rect 7952 18499 8022 18514
rect 7952 18465 7971 18499
rect 8005 18465 8022 18499
rect 7952 18264 8022 18465
rect 8318 18463 8386 18578
rect 8318 18429 8335 18463
rect 8369 18429 8386 18463
rect 8318 18412 8386 18429
rect 9056 18499 9126 18514
rect 9056 18465 9075 18499
rect 9109 18465 9126 18499
rect 9056 18264 9126 18465
rect 9422 18463 9490 18578
rect 9841 18559 9853 18593
rect 9887 18559 9899 18593
rect 9841 18542 9899 18559
rect 10025 18626 10543 18687
rect 10025 18592 10043 18626
rect 10077 18592 10491 18626
rect 10525 18592 10543 18626
rect 10025 18533 10543 18592
rect 10578 18626 11647 18687
rect 10578 18592 10595 18626
rect 10629 18592 11595 18626
rect 11629 18592 11647 18626
rect 10578 18578 11647 18592
rect 11682 18626 12751 18687
rect 11682 18592 11699 18626
rect 11733 18592 12699 18626
rect 12733 18592 12751 18626
rect 11682 18578 12751 18592
rect 12786 18626 13855 18687
rect 12786 18592 12803 18626
rect 12837 18592 13803 18626
rect 13837 18592 13855 18626
rect 12786 18578 13855 18592
rect 13890 18626 14959 18687
rect 13890 18592 13907 18626
rect 13941 18592 14907 18626
rect 14941 18592 14959 18626
rect 13890 18578 14959 18592
rect 14993 18593 15051 18687
rect 9422 18429 9439 18463
rect 9473 18429 9490 18463
rect 9422 18412 9490 18429
rect 10025 18465 10103 18499
rect 10137 18465 10213 18499
rect 10247 18465 10267 18499
rect 9841 18375 9899 18410
rect 9841 18341 9853 18375
rect 9887 18341 9899 18375
rect 9841 18282 9899 18341
rect 4965 18219 4983 18253
rect 5017 18219 5155 18253
rect 5189 18219 5207 18253
rect 4965 18177 5207 18219
rect 5426 18253 6495 18264
rect 5426 18219 5443 18253
rect 5477 18219 6443 18253
rect 6477 18219 6495 18253
rect 5426 18177 6495 18219
rect 6530 18253 7599 18264
rect 6530 18219 6547 18253
rect 6581 18219 7547 18253
rect 7581 18219 7599 18253
rect 6530 18177 7599 18219
rect 7634 18253 8703 18264
rect 7634 18219 7651 18253
rect 7685 18219 8651 18253
rect 8685 18219 8703 18253
rect 7634 18177 8703 18219
rect 8738 18253 9807 18264
rect 8738 18219 8755 18253
rect 8789 18219 9755 18253
rect 9789 18219 9807 18253
rect 8738 18177 9807 18219
rect 9841 18248 9853 18282
rect 9887 18248 9899 18282
rect 9841 18177 9899 18248
rect 10025 18395 10267 18465
rect 10301 18463 10543 18533
rect 10301 18429 10321 18463
rect 10355 18429 10431 18463
rect 10465 18429 10543 18463
rect 10896 18499 10966 18514
rect 10896 18465 10915 18499
rect 10949 18465 10966 18499
rect 10025 18355 10543 18395
rect 10025 18321 10043 18355
rect 10077 18321 10491 18355
rect 10525 18321 10543 18355
rect 10025 18253 10543 18321
rect 10896 18264 10966 18465
rect 11262 18463 11330 18578
rect 11262 18429 11279 18463
rect 11313 18429 11330 18463
rect 11262 18412 11330 18429
rect 12000 18499 12070 18514
rect 12000 18465 12019 18499
rect 12053 18465 12070 18499
rect 12000 18264 12070 18465
rect 12366 18463 12434 18578
rect 12366 18429 12383 18463
rect 12417 18429 12434 18463
rect 12366 18412 12434 18429
rect 13104 18499 13174 18514
rect 13104 18465 13123 18499
rect 13157 18465 13174 18499
rect 13104 18264 13174 18465
rect 13470 18463 13538 18578
rect 13470 18429 13487 18463
rect 13521 18429 13538 18463
rect 13470 18412 13538 18429
rect 14208 18499 14278 18514
rect 14208 18465 14227 18499
rect 14261 18465 14278 18499
rect 14208 18264 14278 18465
rect 14574 18463 14642 18578
rect 14993 18559 15005 18593
rect 15039 18559 15051 18593
rect 14993 18542 15051 18559
rect 15177 18619 15511 18687
rect 15177 18585 15195 18619
rect 15229 18585 15459 18619
rect 15493 18585 15511 18619
rect 15177 18533 15511 18585
rect 15546 18626 16615 18687
rect 15546 18592 15563 18626
rect 15597 18592 16563 18626
rect 16597 18592 16615 18626
rect 15546 18578 16615 18592
rect 16650 18626 17719 18687
rect 16650 18592 16667 18626
rect 16701 18592 17667 18626
rect 17701 18592 17719 18626
rect 16650 18578 17719 18592
rect 17754 18626 18823 18687
rect 17754 18592 17771 18626
rect 17805 18592 18771 18626
rect 18805 18592 18823 18626
rect 17754 18578 18823 18592
rect 18858 18626 19927 18687
rect 18858 18592 18875 18626
rect 18909 18592 19875 18626
rect 19909 18592 19927 18626
rect 18858 18578 19927 18592
rect 19961 18624 20203 18687
rect 19961 18590 19979 18624
rect 20013 18590 20151 18624
rect 20185 18590 20203 18624
rect 14574 18429 14591 18463
rect 14625 18429 14642 18463
rect 14574 18412 14642 18429
rect 15177 18465 15197 18499
rect 15231 18465 15327 18499
rect 14993 18375 15051 18410
rect 14993 18341 15005 18375
rect 15039 18341 15051 18375
rect 14993 18282 15051 18341
rect 10025 18219 10043 18253
rect 10077 18219 10491 18253
rect 10525 18219 10543 18253
rect 10025 18177 10543 18219
rect 10578 18253 11647 18264
rect 10578 18219 10595 18253
rect 10629 18219 11595 18253
rect 11629 18219 11647 18253
rect 10578 18177 11647 18219
rect 11682 18253 12751 18264
rect 11682 18219 11699 18253
rect 11733 18219 12699 18253
rect 12733 18219 12751 18253
rect 11682 18177 12751 18219
rect 12786 18253 13855 18264
rect 12786 18219 12803 18253
rect 12837 18219 13803 18253
rect 13837 18219 13855 18253
rect 12786 18177 13855 18219
rect 13890 18253 14959 18264
rect 13890 18219 13907 18253
rect 13941 18219 14907 18253
rect 14941 18219 14959 18253
rect 13890 18177 14959 18219
rect 14993 18248 15005 18282
rect 15039 18248 15051 18282
rect 14993 18177 15051 18248
rect 15177 18395 15327 18465
rect 15361 18463 15511 18533
rect 15361 18429 15457 18463
rect 15491 18429 15511 18463
rect 15864 18499 15934 18514
rect 15864 18465 15883 18499
rect 15917 18465 15934 18499
rect 15177 18355 15511 18395
rect 15177 18321 15195 18355
rect 15229 18321 15459 18355
rect 15493 18321 15511 18355
rect 15177 18253 15511 18321
rect 15864 18264 15934 18465
rect 16230 18463 16298 18578
rect 16230 18429 16247 18463
rect 16281 18429 16298 18463
rect 16230 18412 16298 18429
rect 16968 18499 17038 18514
rect 16968 18465 16987 18499
rect 17021 18465 17038 18499
rect 16968 18264 17038 18465
rect 17334 18463 17402 18578
rect 17334 18429 17351 18463
rect 17385 18429 17402 18463
rect 17334 18412 17402 18429
rect 18072 18499 18142 18514
rect 18072 18465 18091 18499
rect 18125 18465 18142 18499
rect 18072 18264 18142 18465
rect 18438 18463 18506 18578
rect 18438 18429 18455 18463
rect 18489 18429 18506 18463
rect 18438 18412 18506 18429
rect 19176 18499 19246 18514
rect 19176 18465 19195 18499
rect 19229 18465 19246 18499
rect 19176 18264 19246 18465
rect 19542 18463 19610 18578
rect 19961 18537 20203 18590
rect 19542 18429 19559 18463
rect 19593 18429 19610 18463
rect 19542 18412 19610 18429
rect 19961 18469 20011 18503
rect 20045 18469 20065 18503
rect 19961 18395 20065 18469
rect 20099 18463 20203 18537
rect 20099 18429 20119 18463
rect 20153 18429 20203 18463
rect 19961 18348 20203 18395
rect 19961 18314 19979 18348
rect 20013 18314 20151 18348
rect 20185 18314 20203 18348
rect 15177 18219 15195 18253
rect 15229 18219 15459 18253
rect 15493 18219 15511 18253
rect 15177 18177 15511 18219
rect 15546 18253 16615 18264
rect 15546 18219 15563 18253
rect 15597 18219 16563 18253
rect 16597 18219 16615 18253
rect 15546 18177 16615 18219
rect 16650 18253 17719 18264
rect 16650 18219 16667 18253
rect 16701 18219 17667 18253
rect 17701 18219 17719 18253
rect 16650 18177 17719 18219
rect 17754 18253 18823 18264
rect 17754 18219 17771 18253
rect 17805 18219 18771 18253
rect 18805 18219 18823 18253
rect 17754 18177 18823 18219
rect 18858 18253 19927 18264
rect 18858 18219 18875 18253
rect 18909 18219 19875 18253
rect 19909 18219 19927 18253
rect 18858 18177 19927 18219
rect 19961 18253 20203 18314
rect 19961 18219 19979 18253
rect 20013 18219 20151 18253
rect 20185 18219 20203 18253
rect 19961 18177 20203 18219
rect 4948 18143 4977 18177
rect 5011 18143 5069 18177
rect 5103 18143 5161 18177
rect 5195 18143 5253 18177
rect 5287 18143 5345 18177
rect 5379 18143 5437 18177
rect 5471 18143 5529 18177
rect 5563 18143 5621 18177
rect 5655 18143 5713 18177
rect 5747 18143 5805 18177
rect 5839 18143 5897 18177
rect 5931 18143 5989 18177
rect 6023 18143 6081 18177
rect 6115 18143 6173 18177
rect 6207 18143 6265 18177
rect 6299 18143 6357 18177
rect 6391 18143 6449 18177
rect 6483 18143 6541 18177
rect 6575 18143 6633 18177
rect 6667 18143 6725 18177
rect 6759 18143 6817 18177
rect 6851 18143 6909 18177
rect 6943 18143 7001 18177
rect 7035 18143 7093 18177
rect 7127 18143 7185 18177
rect 7219 18143 7277 18177
rect 7311 18143 7369 18177
rect 7403 18143 7461 18177
rect 7495 18143 7553 18177
rect 7587 18143 7645 18177
rect 7679 18143 7737 18177
rect 7771 18143 7829 18177
rect 7863 18143 7921 18177
rect 7955 18143 8013 18177
rect 8047 18143 8105 18177
rect 8139 18143 8197 18177
rect 8231 18143 8289 18177
rect 8323 18143 8381 18177
rect 8415 18143 8473 18177
rect 8507 18143 8565 18177
rect 8599 18143 8657 18177
rect 8691 18143 8749 18177
rect 8783 18143 8841 18177
rect 8875 18143 8933 18177
rect 8967 18143 9025 18177
rect 9059 18143 9117 18177
rect 9151 18143 9209 18177
rect 9243 18143 9301 18177
rect 9335 18143 9393 18177
rect 9427 18143 9485 18177
rect 9519 18143 9577 18177
rect 9611 18143 9669 18177
rect 9703 18143 9761 18177
rect 9795 18143 9853 18177
rect 9887 18143 9945 18177
rect 9979 18143 10037 18177
rect 10071 18143 10129 18177
rect 10163 18143 10221 18177
rect 10255 18143 10313 18177
rect 10347 18143 10405 18177
rect 10439 18143 10497 18177
rect 10531 18143 10589 18177
rect 10623 18143 10681 18177
rect 10715 18143 10773 18177
rect 10807 18143 10865 18177
rect 10899 18143 10957 18177
rect 10991 18143 11049 18177
rect 11083 18143 11141 18177
rect 11175 18143 11233 18177
rect 11267 18143 11325 18177
rect 11359 18143 11417 18177
rect 11451 18143 11509 18177
rect 11543 18143 11601 18177
rect 11635 18143 11693 18177
rect 11727 18143 11785 18177
rect 11819 18143 11877 18177
rect 11911 18143 11969 18177
rect 12003 18143 12061 18177
rect 12095 18143 12153 18177
rect 12187 18143 12245 18177
rect 12279 18143 12337 18177
rect 12371 18143 12429 18177
rect 12463 18143 12521 18177
rect 12555 18143 12613 18177
rect 12647 18143 12705 18177
rect 12739 18143 12797 18177
rect 12831 18143 12889 18177
rect 12923 18143 12981 18177
rect 13015 18143 13073 18177
rect 13107 18143 13165 18177
rect 13199 18143 13257 18177
rect 13291 18143 13349 18177
rect 13383 18143 13441 18177
rect 13475 18143 13533 18177
rect 13567 18143 13625 18177
rect 13659 18143 13717 18177
rect 13751 18143 13809 18177
rect 13843 18143 13901 18177
rect 13935 18143 13993 18177
rect 14027 18143 14085 18177
rect 14119 18143 14177 18177
rect 14211 18143 14269 18177
rect 14303 18143 14361 18177
rect 14395 18143 14453 18177
rect 14487 18143 14545 18177
rect 14579 18143 14637 18177
rect 14671 18143 14729 18177
rect 14763 18143 14821 18177
rect 14855 18143 14913 18177
rect 14947 18143 15005 18177
rect 15039 18143 15097 18177
rect 15131 18143 15189 18177
rect 15223 18143 15281 18177
rect 15315 18143 15373 18177
rect 15407 18143 15465 18177
rect 15499 18143 15557 18177
rect 15591 18143 15649 18177
rect 15683 18143 15741 18177
rect 15775 18143 15833 18177
rect 15867 18143 15925 18177
rect 15959 18143 16017 18177
rect 16051 18143 16109 18177
rect 16143 18143 16201 18177
rect 16235 18143 16293 18177
rect 16327 18143 16385 18177
rect 16419 18143 16477 18177
rect 16511 18143 16569 18177
rect 16603 18143 16661 18177
rect 16695 18143 16753 18177
rect 16787 18143 16845 18177
rect 16879 18143 16937 18177
rect 16971 18143 17029 18177
rect 17063 18143 17121 18177
rect 17155 18143 17213 18177
rect 17247 18143 17305 18177
rect 17339 18143 17397 18177
rect 17431 18143 17489 18177
rect 17523 18143 17581 18177
rect 17615 18143 17673 18177
rect 17707 18143 17765 18177
rect 17799 18143 17857 18177
rect 17891 18143 17949 18177
rect 17983 18143 18041 18177
rect 18075 18143 18133 18177
rect 18167 18143 18225 18177
rect 18259 18143 18317 18177
rect 18351 18143 18409 18177
rect 18443 18143 18501 18177
rect 18535 18143 18593 18177
rect 18627 18143 18685 18177
rect 18719 18143 18777 18177
rect 18811 18143 18869 18177
rect 18903 18143 18961 18177
rect 18995 18143 19053 18177
rect 19087 18143 19145 18177
rect 19179 18143 19237 18177
rect 19271 18143 19329 18177
rect 19363 18143 19421 18177
rect 19455 18143 19513 18177
rect 19547 18143 19605 18177
rect 19639 18143 19697 18177
rect 19731 18143 19789 18177
rect 19823 18143 19881 18177
rect 19915 18143 19973 18177
rect 20007 18143 20065 18177
rect 20099 18143 20157 18177
rect 20191 18143 20220 18177
rect 4965 18101 5207 18143
rect 4965 18067 4983 18101
rect 5017 18067 5155 18101
rect 5189 18067 5207 18101
rect 4965 18006 5207 18067
rect 4965 17972 4983 18006
rect 5017 17972 5155 18006
rect 5189 17972 5207 18006
rect 4965 17925 5207 17972
rect 4965 17857 5015 17891
rect 5049 17857 5069 17891
rect 4965 17783 5069 17857
rect 5103 17851 5207 17925
rect 5103 17817 5123 17851
rect 5157 17817 5207 17851
rect 5425 18101 6127 18143
rect 5425 18067 5443 18101
rect 5477 18067 6075 18101
rect 6109 18067 6127 18101
rect 5425 17999 6127 18067
rect 6162 18101 7231 18143
rect 6162 18067 6179 18101
rect 6213 18067 7179 18101
rect 7213 18067 7231 18101
rect 6162 18056 7231 18067
rect 7265 18072 7323 18143
rect 5425 17965 5443 17999
rect 5477 17965 6075 17999
rect 6109 17965 6127 17999
rect 5425 17925 6127 17965
rect 5425 17855 5763 17925
rect 5425 17821 5503 17855
rect 5537 17821 5606 17855
rect 5640 17821 5709 17855
rect 5743 17821 5763 17855
rect 5797 17857 5817 17891
rect 5851 17857 5916 17891
rect 5950 17857 6015 17891
rect 6049 17857 6127 17891
rect 5797 17787 6127 17857
rect 6480 17855 6550 18056
rect 7265 18038 7277 18072
rect 7311 18038 7323 18072
rect 7265 17979 7323 18038
rect 7265 17945 7277 17979
rect 7311 17945 7323 17979
rect 7265 17910 7323 17945
rect 7449 18101 7967 18143
rect 7449 18067 7467 18101
rect 7501 18067 7915 18101
rect 7949 18067 7967 18101
rect 7449 17999 7967 18067
rect 8002 18101 9071 18143
rect 8002 18067 8019 18101
rect 8053 18067 9019 18101
rect 9053 18067 9071 18101
rect 8002 18056 9071 18067
rect 9106 18101 10175 18143
rect 9106 18067 9123 18101
rect 9157 18067 10123 18101
rect 10157 18067 10175 18101
rect 9106 18056 10175 18067
rect 10210 18101 11279 18143
rect 10210 18067 10227 18101
rect 10261 18067 11227 18101
rect 11261 18067 11279 18101
rect 10210 18056 11279 18067
rect 11314 18101 12383 18143
rect 11314 18067 11331 18101
rect 11365 18067 12331 18101
rect 12365 18067 12383 18101
rect 11314 18056 12383 18067
rect 12417 18072 12475 18143
rect 7449 17965 7467 17999
rect 7501 17965 7915 17999
rect 7949 17965 7967 17999
rect 7449 17925 7967 17965
rect 6480 17821 6499 17855
rect 6533 17821 6550 17855
rect 6480 17806 6550 17821
rect 6846 17891 6914 17908
rect 6846 17857 6863 17891
rect 6897 17857 6914 17891
rect 4965 17730 5207 17783
rect 4965 17696 4983 17730
rect 5017 17696 5155 17730
rect 5189 17696 5207 17730
rect 4965 17633 5207 17696
rect 5425 17728 6127 17787
rect 6846 17742 6914 17857
rect 7449 17855 7691 17925
rect 7449 17821 7527 17855
rect 7561 17821 7637 17855
rect 7671 17821 7691 17855
rect 7725 17857 7745 17891
rect 7779 17857 7855 17891
rect 7889 17857 7967 17891
rect 7725 17787 7967 17857
rect 8320 17855 8390 18056
rect 8320 17821 8339 17855
rect 8373 17821 8390 17855
rect 8320 17806 8390 17821
rect 8686 17891 8754 17908
rect 8686 17857 8703 17891
rect 8737 17857 8754 17891
rect 7265 17761 7323 17778
rect 5425 17694 5443 17728
rect 5477 17694 6075 17728
rect 6109 17694 6127 17728
rect 5425 17633 6127 17694
rect 6162 17728 7231 17742
rect 6162 17694 6179 17728
rect 6213 17694 7179 17728
rect 7213 17694 7231 17728
rect 6162 17633 7231 17694
rect 7265 17727 7277 17761
rect 7311 17727 7323 17761
rect 7265 17633 7323 17727
rect 7449 17728 7967 17787
rect 8686 17742 8754 17857
rect 9424 17855 9494 18056
rect 9424 17821 9443 17855
rect 9477 17821 9494 17855
rect 9424 17806 9494 17821
rect 9790 17891 9858 17908
rect 9790 17857 9807 17891
rect 9841 17857 9858 17891
rect 9790 17742 9858 17857
rect 10528 17855 10598 18056
rect 10528 17821 10547 17855
rect 10581 17821 10598 17855
rect 10528 17806 10598 17821
rect 10894 17891 10962 17908
rect 10894 17857 10911 17891
rect 10945 17857 10962 17891
rect 10894 17742 10962 17857
rect 11632 17855 11702 18056
rect 12417 18038 12429 18072
rect 12463 18038 12475 18072
rect 12417 17979 12475 18038
rect 12417 17945 12429 17979
rect 12463 17945 12475 17979
rect 12417 17910 12475 17945
rect 12601 18101 13119 18143
rect 12601 18067 12619 18101
rect 12653 18067 13067 18101
rect 13101 18067 13119 18101
rect 12601 17999 13119 18067
rect 13154 18101 14223 18143
rect 13154 18067 13171 18101
rect 13205 18067 14171 18101
rect 14205 18067 14223 18101
rect 13154 18056 14223 18067
rect 14258 18101 15327 18143
rect 14258 18067 14275 18101
rect 14309 18067 15275 18101
rect 15309 18067 15327 18101
rect 14258 18056 15327 18067
rect 15362 18101 16431 18143
rect 15362 18067 15379 18101
rect 15413 18067 16379 18101
rect 16413 18067 16431 18101
rect 15362 18056 16431 18067
rect 16466 18101 17535 18143
rect 16466 18067 16483 18101
rect 16517 18067 17483 18101
rect 17517 18067 17535 18101
rect 16466 18056 17535 18067
rect 17569 18072 17627 18143
rect 12601 17965 12619 17999
rect 12653 17965 13067 17999
rect 13101 17965 13119 17999
rect 12601 17925 13119 17965
rect 11632 17821 11651 17855
rect 11685 17821 11702 17855
rect 11632 17806 11702 17821
rect 11998 17891 12066 17908
rect 11998 17857 12015 17891
rect 12049 17857 12066 17891
rect 11998 17742 12066 17857
rect 12601 17855 12843 17925
rect 12601 17821 12679 17855
rect 12713 17821 12789 17855
rect 12823 17821 12843 17855
rect 12877 17857 12897 17891
rect 12931 17857 13007 17891
rect 13041 17857 13119 17891
rect 12877 17787 13119 17857
rect 13472 17855 13542 18056
rect 13472 17821 13491 17855
rect 13525 17821 13542 17855
rect 13472 17806 13542 17821
rect 13838 17891 13906 17908
rect 13838 17857 13855 17891
rect 13889 17857 13906 17891
rect 12417 17761 12475 17778
rect 7449 17694 7467 17728
rect 7501 17694 7915 17728
rect 7949 17694 7967 17728
rect 7449 17633 7967 17694
rect 8002 17728 9071 17742
rect 8002 17694 8019 17728
rect 8053 17694 9019 17728
rect 9053 17694 9071 17728
rect 8002 17633 9071 17694
rect 9106 17728 10175 17742
rect 9106 17694 9123 17728
rect 9157 17694 10123 17728
rect 10157 17694 10175 17728
rect 9106 17633 10175 17694
rect 10210 17728 11279 17742
rect 10210 17694 10227 17728
rect 10261 17694 11227 17728
rect 11261 17694 11279 17728
rect 10210 17633 11279 17694
rect 11314 17728 12383 17742
rect 11314 17694 11331 17728
rect 11365 17694 12331 17728
rect 12365 17694 12383 17728
rect 11314 17633 12383 17694
rect 12417 17727 12429 17761
rect 12463 17727 12475 17761
rect 12417 17633 12475 17727
rect 12601 17728 13119 17787
rect 13838 17742 13906 17857
rect 14576 17855 14646 18056
rect 14576 17821 14595 17855
rect 14629 17821 14646 17855
rect 14576 17806 14646 17821
rect 14942 17891 15010 17908
rect 14942 17857 14959 17891
rect 14993 17857 15010 17891
rect 14942 17742 15010 17857
rect 15680 17855 15750 18056
rect 15680 17821 15699 17855
rect 15733 17821 15750 17855
rect 15680 17806 15750 17821
rect 16046 17891 16114 17908
rect 16046 17857 16063 17891
rect 16097 17857 16114 17891
rect 16046 17742 16114 17857
rect 16784 17855 16854 18056
rect 17569 18038 17581 18072
rect 17615 18038 17627 18072
rect 17754 18101 18823 18143
rect 17754 18067 17771 18101
rect 17805 18067 18771 18101
rect 18805 18067 18823 18101
rect 17754 18056 18823 18067
rect 18858 18101 19927 18143
rect 18858 18067 18875 18101
rect 18909 18067 19875 18101
rect 19909 18067 19927 18101
rect 18858 18056 19927 18067
rect 19961 18101 20203 18143
rect 19961 18067 19979 18101
rect 20013 18067 20151 18101
rect 20185 18067 20203 18101
rect 17569 17979 17627 18038
rect 17569 17945 17581 17979
rect 17615 17945 17627 17979
rect 17569 17910 17627 17945
rect 16784 17821 16803 17855
rect 16837 17821 16854 17855
rect 16784 17806 16854 17821
rect 17150 17891 17218 17908
rect 17150 17857 17167 17891
rect 17201 17857 17218 17891
rect 17150 17742 17218 17857
rect 18072 17855 18142 18056
rect 18072 17821 18091 17855
rect 18125 17821 18142 17855
rect 18072 17806 18142 17821
rect 18438 17891 18506 17908
rect 18438 17857 18455 17891
rect 18489 17857 18506 17891
rect 17569 17761 17627 17778
rect 12601 17694 12619 17728
rect 12653 17694 13067 17728
rect 13101 17694 13119 17728
rect 12601 17633 13119 17694
rect 13154 17728 14223 17742
rect 13154 17694 13171 17728
rect 13205 17694 14171 17728
rect 14205 17694 14223 17728
rect 13154 17633 14223 17694
rect 14258 17728 15327 17742
rect 14258 17694 14275 17728
rect 14309 17694 15275 17728
rect 15309 17694 15327 17728
rect 14258 17633 15327 17694
rect 15362 17728 16431 17742
rect 15362 17694 15379 17728
rect 15413 17694 16379 17728
rect 16413 17694 16431 17728
rect 15362 17633 16431 17694
rect 16466 17728 17535 17742
rect 16466 17694 16483 17728
rect 16517 17694 17483 17728
rect 17517 17694 17535 17728
rect 16466 17633 17535 17694
rect 17569 17727 17581 17761
rect 17615 17727 17627 17761
rect 18438 17742 18506 17857
rect 19176 17855 19246 18056
rect 19961 18006 20203 18067
rect 19961 17972 19979 18006
rect 20013 17972 20151 18006
rect 20185 17972 20203 18006
rect 19961 17925 20203 17972
rect 19176 17821 19195 17855
rect 19229 17821 19246 17855
rect 19176 17806 19246 17821
rect 19542 17891 19610 17908
rect 19542 17857 19559 17891
rect 19593 17857 19610 17891
rect 19542 17742 19610 17857
rect 19961 17851 20065 17925
rect 19961 17817 20011 17851
rect 20045 17817 20065 17851
rect 20099 17857 20119 17891
rect 20153 17857 20203 17891
rect 20099 17783 20203 17857
rect 17569 17633 17627 17727
rect 17754 17728 18823 17742
rect 17754 17694 17771 17728
rect 17805 17694 18771 17728
rect 18805 17694 18823 17728
rect 17754 17633 18823 17694
rect 18858 17728 19927 17742
rect 18858 17694 18875 17728
rect 18909 17694 19875 17728
rect 19909 17694 19927 17728
rect 18858 17633 19927 17694
rect 19961 17730 20203 17783
rect 19961 17696 19979 17730
rect 20013 17696 20151 17730
rect 20185 17696 20203 17730
rect 19961 17633 20203 17696
rect 4948 17599 4977 17633
rect 5011 17599 5069 17633
rect 5103 17599 5161 17633
rect 5195 17599 5253 17633
rect 5287 17599 5345 17633
rect 5379 17599 5437 17633
rect 5471 17599 5529 17633
rect 5563 17599 5621 17633
rect 5655 17599 5713 17633
rect 5747 17599 5805 17633
rect 5839 17599 5897 17633
rect 5931 17599 5989 17633
rect 6023 17599 6081 17633
rect 6115 17599 6173 17633
rect 6207 17599 6265 17633
rect 6299 17599 6357 17633
rect 6391 17599 6449 17633
rect 6483 17599 6541 17633
rect 6575 17599 6633 17633
rect 6667 17599 6725 17633
rect 6759 17599 6817 17633
rect 6851 17599 6909 17633
rect 6943 17599 7001 17633
rect 7035 17599 7093 17633
rect 7127 17599 7185 17633
rect 7219 17599 7277 17633
rect 7311 17599 7369 17633
rect 7403 17599 7461 17633
rect 7495 17599 7553 17633
rect 7587 17599 7645 17633
rect 7679 17599 7737 17633
rect 7771 17599 7829 17633
rect 7863 17599 7921 17633
rect 7955 17599 8013 17633
rect 8047 17599 8105 17633
rect 8139 17599 8197 17633
rect 8231 17599 8289 17633
rect 8323 17599 8381 17633
rect 8415 17599 8473 17633
rect 8507 17599 8565 17633
rect 8599 17599 8657 17633
rect 8691 17599 8749 17633
rect 8783 17599 8841 17633
rect 8875 17599 8933 17633
rect 8967 17599 9025 17633
rect 9059 17599 9117 17633
rect 9151 17599 9209 17633
rect 9243 17599 9301 17633
rect 9335 17599 9393 17633
rect 9427 17599 9485 17633
rect 9519 17599 9577 17633
rect 9611 17599 9669 17633
rect 9703 17599 9761 17633
rect 9795 17599 9853 17633
rect 9887 17599 9945 17633
rect 9979 17599 10037 17633
rect 10071 17599 10129 17633
rect 10163 17599 10221 17633
rect 10255 17599 10313 17633
rect 10347 17599 10405 17633
rect 10439 17599 10497 17633
rect 10531 17599 10589 17633
rect 10623 17599 10681 17633
rect 10715 17599 10773 17633
rect 10807 17599 10865 17633
rect 10899 17599 10957 17633
rect 10991 17599 11049 17633
rect 11083 17599 11141 17633
rect 11175 17599 11233 17633
rect 11267 17599 11325 17633
rect 11359 17599 11417 17633
rect 11451 17599 11509 17633
rect 11543 17599 11601 17633
rect 11635 17599 11693 17633
rect 11727 17599 11785 17633
rect 11819 17599 11877 17633
rect 11911 17599 11969 17633
rect 12003 17599 12061 17633
rect 12095 17599 12153 17633
rect 12187 17599 12245 17633
rect 12279 17599 12337 17633
rect 12371 17599 12429 17633
rect 12463 17599 12521 17633
rect 12555 17599 12613 17633
rect 12647 17599 12705 17633
rect 12739 17599 12797 17633
rect 12831 17599 12889 17633
rect 12923 17599 12981 17633
rect 13015 17599 13073 17633
rect 13107 17599 13165 17633
rect 13199 17599 13257 17633
rect 13291 17599 13349 17633
rect 13383 17599 13441 17633
rect 13475 17599 13533 17633
rect 13567 17599 13625 17633
rect 13659 17599 13717 17633
rect 13751 17599 13809 17633
rect 13843 17599 13901 17633
rect 13935 17599 13993 17633
rect 14027 17599 14085 17633
rect 14119 17599 14177 17633
rect 14211 17599 14269 17633
rect 14303 17599 14361 17633
rect 14395 17599 14453 17633
rect 14487 17599 14545 17633
rect 14579 17599 14637 17633
rect 14671 17599 14729 17633
rect 14763 17599 14821 17633
rect 14855 17599 14913 17633
rect 14947 17599 15005 17633
rect 15039 17599 15097 17633
rect 15131 17599 15189 17633
rect 15223 17599 15281 17633
rect 15315 17599 15373 17633
rect 15407 17599 15465 17633
rect 15499 17599 15557 17633
rect 15591 17599 15649 17633
rect 15683 17599 15741 17633
rect 15775 17599 15833 17633
rect 15867 17599 15925 17633
rect 15959 17599 16017 17633
rect 16051 17599 16109 17633
rect 16143 17599 16201 17633
rect 16235 17599 16293 17633
rect 16327 17599 16385 17633
rect 16419 17599 16477 17633
rect 16511 17599 16569 17633
rect 16603 17599 16661 17633
rect 16695 17599 16753 17633
rect 16787 17599 16845 17633
rect 16879 17599 16937 17633
rect 16971 17599 17029 17633
rect 17063 17599 17121 17633
rect 17155 17599 17213 17633
rect 17247 17599 17305 17633
rect 17339 17599 17397 17633
rect 17431 17599 17489 17633
rect 17523 17599 17581 17633
rect 17615 17599 17673 17633
rect 17707 17599 17765 17633
rect 17799 17599 17857 17633
rect 17891 17599 17949 17633
rect 17983 17599 18041 17633
rect 18075 17599 18133 17633
rect 18167 17599 18225 17633
rect 18259 17599 18317 17633
rect 18351 17599 18409 17633
rect 18443 17599 18501 17633
rect 18535 17599 18593 17633
rect 18627 17599 18685 17633
rect 18719 17599 18777 17633
rect 18811 17599 18869 17633
rect 18903 17599 18961 17633
rect 18995 17599 19053 17633
rect 19087 17599 19145 17633
rect 19179 17599 19237 17633
rect 19271 17599 19329 17633
rect 19363 17599 19421 17633
rect 19455 17599 19513 17633
rect 19547 17599 19605 17633
rect 19639 17599 19697 17633
rect 19731 17599 19789 17633
rect 19823 17599 19881 17633
rect 19915 17599 19973 17633
rect 20007 17599 20065 17633
rect 20099 17599 20157 17633
rect 20191 17599 20220 17633
rect 4965 17536 5207 17599
rect 4965 17502 4983 17536
rect 5017 17502 5155 17536
rect 5189 17502 5207 17536
rect 4965 17449 5207 17502
rect 5426 17538 6495 17599
rect 5426 17504 5443 17538
rect 5477 17504 6443 17538
rect 6477 17504 6495 17538
rect 5426 17490 6495 17504
rect 6530 17538 7599 17599
rect 6530 17504 6547 17538
rect 6581 17504 7547 17538
rect 7581 17504 7599 17538
rect 6530 17490 7599 17504
rect 7634 17538 8703 17599
rect 7634 17504 7651 17538
rect 7685 17504 8651 17538
rect 8685 17504 8703 17538
rect 7634 17490 8703 17504
rect 8738 17538 9807 17599
rect 8738 17504 8755 17538
rect 8789 17504 9755 17538
rect 9789 17504 9807 17538
rect 8738 17490 9807 17504
rect 9841 17505 9899 17599
rect 4965 17375 5069 17449
rect 4965 17341 5015 17375
rect 5049 17341 5069 17375
rect 5103 17381 5123 17415
rect 5157 17381 5207 17415
rect 5103 17307 5207 17381
rect 4965 17260 5207 17307
rect 4965 17226 4983 17260
rect 5017 17226 5155 17260
rect 5189 17226 5207 17260
rect 4965 17165 5207 17226
rect 5744 17411 5814 17426
rect 5744 17377 5763 17411
rect 5797 17377 5814 17411
rect 5744 17176 5814 17377
rect 6110 17375 6178 17490
rect 6110 17341 6127 17375
rect 6161 17341 6178 17375
rect 6110 17324 6178 17341
rect 6848 17411 6918 17426
rect 6848 17377 6867 17411
rect 6901 17377 6918 17411
rect 6848 17176 6918 17377
rect 7214 17375 7282 17490
rect 7214 17341 7231 17375
rect 7265 17341 7282 17375
rect 7214 17324 7282 17341
rect 7952 17411 8022 17426
rect 7952 17377 7971 17411
rect 8005 17377 8022 17411
rect 7952 17176 8022 17377
rect 8318 17375 8386 17490
rect 8318 17341 8335 17375
rect 8369 17341 8386 17375
rect 8318 17324 8386 17341
rect 9056 17411 9126 17426
rect 9056 17377 9075 17411
rect 9109 17377 9126 17411
rect 9056 17176 9126 17377
rect 9422 17375 9490 17490
rect 9841 17471 9853 17505
rect 9887 17471 9899 17505
rect 9841 17454 9899 17471
rect 10025 17538 10543 17599
rect 10025 17504 10043 17538
rect 10077 17504 10491 17538
rect 10525 17504 10543 17538
rect 10025 17445 10543 17504
rect 10578 17538 11647 17599
rect 10578 17504 10595 17538
rect 10629 17504 11595 17538
rect 11629 17504 11647 17538
rect 10578 17490 11647 17504
rect 11682 17538 12751 17599
rect 11682 17504 11699 17538
rect 11733 17504 12699 17538
rect 12733 17504 12751 17538
rect 11682 17490 12751 17504
rect 12786 17538 13855 17599
rect 12786 17504 12803 17538
rect 12837 17504 13803 17538
rect 13837 17504 13855 17538
rect 12786 17490 13855 17504
rect 13890 17538 14959 17599
rect 13890 17504 13907 17538
rect 13941 17504 14907 17538
rect 14941 17504 14959 17538
rect 13890 17490 14959 17504
rect 14993 17505 15051 17599
rect 9422 17341 9439 17375
rect 9473 17341 9490 17375
rect 9422 17324 9490 17341
rect 10025 17377 10103 17411
rect 10137 17377 10213 17411
rect 10247 17377 10267 17411
rect 9841 17287 9899 17322
rect 9841 17253 9853 17287
rect 9887 17253 9899 17287
rect 9841 17194 9899 17253
rect 4965 17131 4983 17165
rect 5017 17131 5155 17165
rect 5189 17131 5207 17165
rect 4965 17089 5207 17131
rect 5426 17165 6495 17176
rect 5426 17131 5443 17165
rect 5477 17131 6443 17165
rect 6477 17131 6495 17165
rect 5426 17089 6495 17131
rect 6530 17165 7599 17176
rect 6530 17131 6547 17165
rect 6581 17131 7547 17165
rect 7581 17131 7599 17165
rect 6530 17089 7599 17131
rect 7634 17165 8703 17176
rect 7634 17131 7651 17165
rect 7685 17131 8651 17165
rect 8685 17131 8703 17165
rect 7634 17089 8703 17131
rect 8738 17165 9807 17176
rect 8738 17131 8755 17165
rect 8789 17131 9755 17165
rect 9789 17131 9807 17165
rect 8738 17089 9807 17131
rect 9841 17160 9853 17194
rect 9887 17160 9899 17194
rect 9841 17089 9899 17160
rect 10025 17307 10267 17377
rect 10301 17375 10543 17445
rect 10301 17341 10321 17375
rect 10355 17341 10431 17375
rect 10465 17341 10543 17375
rect 10896 17411 10966 17426
rect 10896 17377 10915 17411
rect 10949 17377 10966 17411
rect 10025 17267 10543 17307
rect 10025 17233 10043 17267
rect 10077 17233 10491 17267
rect 10525 17233 10543 17267
rect 10025 17165 10543 17233
rect 10896 17176 10966 17377
rect 11262 17375 11330 17490
rect 11262 17341 11279 17375
rect 11313 17341 11330 17375
rect 11262 17324 11330 17341
rect 12000 17411 12070 17426
rect 12000 17377 12019 17411
rect 12053 17377 12070 17411
rect 12000 17176 12070 17377
rect 12366 17375 12434 17490
rect 12366 17341 12383 17375
rect 12417 17341 12434 17375
rect 12366 17324 12434 17341
rect 13104 17411 13174 17426
rect 13104 17377 13123 17411
rect 13157 17377 13174 17411
rect 13104 17176 13174 17377
rect 13470 17375 13538 17490
rect 13470 17341 13487 17375
rect 13521 17341 13538 17375
rect 13470 17324 13538 17341
rect 14208 17411 14278 17426
rect 14208 17377 14227 17411
rect 14261 17377 14278 17411
rect 14208 17176 14278 17377
rect 14574 17375 14642 17490
rect 14993 17471 15005 17505
rect 15039 17471 15051 17505
rect 14993 17454 15051 17471
rect 15177 17531 15511 17599
rect 15177 17497 15195 17531
rect 15229 17497 15459 17531
rect 15493 17497 15511 17531
rect 15177 17445 15511 17497
rect 15546 17538 16615 17599
rect 15546 17504 15563 17538
rect 15597 17504 16563 17538
rect 16597 17504 16615 17538
rect 15546 17490 16615 17504
rect 16650 17538 17719 17599
rect 16650 17504 16667 17538
rect 16701 17504 17667 17538
rect 17701 17504 17719 17538
rect 16650 17490 17719 17504
rect 17754 17538 18823 17599
rect 17754 17504 17771 17538
rect 17805 17504 18771 17538
rect 18805 17504 18823 17538
rect 17754 17490 18823 17504
rect 18858 17538 19927 17599
rect 18858 17504 18875 17538
rect 18909 17504 19875 17538
rect 19909 17504 19927 17538
rect 18858 17490 19927 17504
rect 19961 17536 20203 17599
rect 19961 17502 19979 17536
rect 20013 17502 20151 17536
rect 20185 17502 20203 17536
rect 14574 17341 14591 17375
rect 14625 17341 14642 17375
rect 14574 17324 14642 17341
rect 15177 17377 15197 17411
rect 15231 17377 15327 17411
rect 14993 17287 15051 17322
rect 14993 17253 15005 17287
rect 15039 17253 15051 17287
rect 14993 17194 15051 17253
rect 10025 17131 10043 17165
rect 10077 17131 10491 17165
rect 10525 17131 10543 17165
rect 10025 17089 10543 17131
rect 10578 17165 11647 17176
rect 10578 17131 10595 17165
rect 10629 17131 11595 17165
rect 11629 17131 11647 17165
rect 10578 17089 11647 17131
rect 11682 17165 12751 17176
rect 11682 17131 11699 17165
rect 11733 17131 12699 17165
rect 12733 17131 12751 17165
rect 11682 17089 12751 17131
rect 12786 17165 13855 17176
rect 12786 17131 12803 17165
rect 12837 17131 13803 17165
rect 13837 17131 13855 17165
rect 12786 17089 13855 17131
rect 13890 17165 14959 17176
rect 13890 17131 13907 17165
rect 13941 17131 14907 17165
rect 14941 17131 14959 17165
rect 13890 17089 14959 17131
rect 14993 17160 15005 17194
rect 15039 17160 15051 17194
rect 14993 17089 15051 17160
rect 15177 17307 15327 17377
rect 15361 17375 15511 17445
rect 15361 17341 15457 17375
rect 15491 17341 15511 17375
rect 15864 17411 15934 17426
rect 15864 17377 15883 17411
rect 15917 17377 15934 17411
rect 15177 17267 15511 17307
rect 15177 17233 15195 17267
rect 15229 17233 15459 17267
rect 15493 17233 15511 17267
rect 15177 17165 15511 17233
rect 15864 17176 15934 17377
rect 16230 17375 16298 17490
rect 16230 17341 16247 17375
rect 16281 17341 16298 17375
rect 16230 17324 16298 17341
rect 16968 17411 17038 17426
rect 16968 17377 16987 17411
rect 17021 17377 17038 17411
rect 16968 17176 17038 17377
rect 17334 17375 17402 17490
rect 17334 17341 17351 17375
rect 17385 17341 17402 17375
rect 17334 17324 17402 17341
rect 18072 17411 18142 17426
rect 18072 17377 18091 17411
rect 18125 17377 18142 17411
rect 18072 17176 18142 17377
rect 18438 17375 18506 17490
rect 18438 17341 18455 17375
rect 18489 17341 18506 17375
rect 18438 17324 18506 17341
rect 19176 17411 19246 17426
rect 19176 17377 19195 17411
rect 19229 17377 19246 17411
rect 19176 17176 19246 17377
rect 19542 17375 19610 17490
rect 19961 17449 20203 17502
rect 19542 17341 19559 17375
rect 19593 17341 19610 17375
rect 19542 17324 19610 17341
rect 19961 17381 20011 17415
rect 20045 17381 20065 17415
rect 19961 17307 20065 17381
rect 20099 17375 20203 17449
rect 20099 17341 20119 17375
rect 20153 17341 20203 17375
rect 19961 17260 20203 17307
rect 19961 17226 19979 17260
rect 20013 17226 20151 17260
rect 20185 17226 20203 17260
rect 15177 17131 15195 17165
rect 15229 17131 15459 17165
rect 15493 17131 15511 17165
rect 15177 17089 15511 17131
rect 15546 17165 16615 17176
rect 15546 17131 15563 17165
rect 15597 17131 16563 17165
rect 16597 17131 16615 17165
rect 15546 17089 16615 17131
rect 16650 17165 17719 17176
rect 16650 17131 16667 17165
rect 16701 17131 17667 17165
rect 17701 17131 17719 17165
rect 16650 17089 17719 17131
rect 17754 17165 18823 17176
rect 17754 17131 17771 17165
rect 17805 17131 18771 17165
rect 18805 17131 18823 17165
rect 17754 17089 18823 17131
rect 18858 17165 19927 17176
rect 18858 17131 18875 17165
rect 18909 17131 19875 17165
rect 19909 17131 19927 17165
rect 18858 17089 19927 17131
rect 19961 17165 20203 17226
rect 19961 17131 19979 17165
rect 20013 17131 20151 17165
rect 20185 17131 20203 17165
rect 19961 17089 20203 17131
rect 4948 17055 4977 17089
rect 5011 17055 5069 17089
rect 5103 17055 5161 17089
rect 5195 17055 5253 17089
rect 5287 17055 5345 17089
rect 5379 17055 5437 17089
rect 5471 17055 5529 17089
rect 5563 17055 5621 17089
rect 5655 17055 5713 17089
rect 5747 17055 5805 17089
rect 5839 17055 5897 17089
rect 5931 17055 5989 17089
rect 6023 17055 6081 17089
rect 6115 17055 6173 17089
rect 6207 17055 6265 17089
rect 6299 17055 6357 17089
rect 6391 17055 6449 17089
rect 6483 17055 6541 17089
rect 6575 17055 6633 17089
rect 6667 17055 6725 17089
rect 6759 17055 6817 17089
rect 6851 17055 6909 17089
rect 6943 17055 7001 17089
rect 7035 17055 7093 17089
rect 7127 17055 7185 17089
rect 7219 17055 7277 17089
rect 7311 17055 7369 17089
rect 7403 17055 7461 17089
rect 7495 17055 7553 17089
rect 7587 17055 7645 17089
rect 7679 17055 7737 17089
rect 7771 17055 7829 17089
rect 7863 17055 7921 17089
rect 7955 17055 8013 17089
rect 8047 17055 8105 17089
rect 8139 17055 8197 17089
rect 8231 17055 8289 17089
rect 8323 17055 8381 17089
rect 8415 17055 8473 17089
rect 8507 17055 8565 17089
rect 8599 17055 8657 17089
rect 8691 17055 8749 17089
rect 8783 17055 8841 17089
rect 8875 17055 8933 17089
rect 8967 17055 9025 17089
rect 9059 17055 9117 17089
rect 9151 17055 9209 17089
rect 9243 17055 9301 17089
rect 9335 17055 9393 17089
rect 9427 17055 9485 17089
rect 9519 17055 9577 17089
rect 9611 17055 9669 17089
rect 9703 17055 9761 17089
rect 9795 17055 9853 17089
rect 9887 17055 9945 17089
rect 9979 17055 10037 17089
rect 10071 17055 10129 17089
rect 10163 17055 10221 17089
rect 10255 17055 10313 17089
rect 10347 17055 10405 17089
rect 10439 17055 10497 17089
rect 10531 17055 10589 17089
rect 10623 17055 10681 17089
rect 10715 17055 10773 17089
rect 10807 17055 10865 17089
rect 10899 17055 10957 17089
rect 10991 17055 11049 17089
rect 11083 17055 11141 17089
rect 11175 17055 11233 17089
rect 11267 17055 11325 17089
rect 11359 17055 11417 17089
rect 11451 17055 11509 17089
rect 11543 17055 11601 17089
rect 11635 17055 11693 17089
rect 11727 17055 11785 17089
rect 11819 17055 11877 17089
rect 11911 17055 11969 17089
rect 12003 17055 12061 17089
rect 12095 17055 12153 17089
rect 12187 17055 12245 17089
rect 12279 17055 12337 17089
rect 12371 17055 12429 17089
rect 12463 17055 12521 17089
rect 12555 17055 12613 17089
rect 12647 17055 12705 17089
rect 12739 17055 12797 17089
rect 12831 17055 12889 17089
rect 12923 17055 12981 17089
rect 13015 17055 13073 17089
rect 13107 17055 13165 17089
rect 13199 17055 13257 17089
rect 13291 17055 13349 17089
rect 13383 17055 13441 17089
rect 13475 17055 13533 17089
rect 13567 17055 13625 17089
rect 13659 17055 13717 17089
rect 13751 17055 13809 17089
rect 13843 17055 13901 17089
rect 13935 17055 13993 17089
rect 14027 17055 14085 17089
rect 14119 17055 14177 17089
rect 14211 17055 14269 17089
rect 14303 17055 14361 17089
rect 14395 17055 14453 17089
rect 14487 17055 14545 17089
rect 14579 17055 14637 17089
rect 14671 17055 14729 17089
rect 14763 17055 14821 17089
rect 14855 17055 14913 17089
rect 14947 17055 15005 17089
rect 15039 17055 15097 17089
rect 15131 17055 15189 17089
rect 15223 17055 15281 17089
rect 15315 17055 15373 17089
rect 15407 17055 15465 17089
rect 15499 17055 15557 17089
rect 15591 17055 15649 17089
rect 15683 17055 15741 17089
rect 15775 17055 15833 17089
rect 15867 17055 15925 17089
rect 15959 17055 16017 17089
rect 16051 17055 16109 17089
rect 16143 17055 16201 17089
rect 16235 17055 16293 17089
rect 16327 17055 16385 17089
rect 16419 17055 16477 17089
rect 16511 17055 16569 17089
rect 16603 17055 16661 17089
rect 16695 17055 16753 17089
rect 16787 17055 16845 17089
rect 16879 17055 16937 17089
rect 16971 17055 17029 17089
rect 17063 17055 17121 17089
rect 17155 17055 17213 17089
rect 17247 17055 17305 17089
rect 17339 17055 17397 17089
rect 17431 17055 17489 17089
rect 17523 17055 17581 17089
rect 17615 17055 17673 17089
rect 17707 17055 17765 17089
rect 17799 17055 17857 17089
rect 17891 17055 17949 17089
rect 17983 17055 18041 17089
rect 18075 17055 18133 17089
rect 18167 17055 18225 17089
rect 18259 17055 18317 17089
rect 18351 17055 18409 17089
rect 18443 17055 18501 17089
rect 18535 17055 18593 17089
rect 18627 17055 18685 17089
rect 18719 17055 18777 17089
rect 18811 17055 18869 17089
rect 18903 17055 18961 17089
rect 18995 17055 19053 17089
rect 19087 17055 19145 17089
rect 19179 17055 19237 17089
rect 19271 17055 19329 17089
rect 19363 17055 19421 17089
rect 19455 17055 19513 17089
rect 19547 17055 19605 17089
rect 19639 17055 19697 17089
rect 19731 17055 19789 17089
rect 19823 17055 19881 17089
rect 19915 17055 19973 17089
rect 20007 17055 20065 17089
rect 20099 17055 20157 17089
rect 20191 17055 20220 17089
rect 4965 17013 5207 17055
rect 4965 16979 4983 17013
rect 5017 16979 5155 17013
rect 5189 16979 5207 17013
rect 4965 16918 5207 16979
rect 4965 16884 4983 16918
rect 5017 16884 5155 16918
rect 5189 16884 5207 16918
rect 4965 16837 5207 16884
rect 4965 16769 5015 16803
rect 5049 16769 5069 16803
rect 4965 16695 5069 16769
rect 5103 16763 5207 16837
rect 5103 16729 5123 16763
rect 5157 16729 5207 16763
rect 5425 17013 6127 17055
rect 5425 16979 5443 17013
rect 5477 16979 6075 17013
rect 6109 16979 6127 17013
rect 5425 16911 6127 16979
rect 6162 17013 7231 17055
rect 6162 16979 6179 17013
rect 6213 16979 7179 17013
rect 7213 16979 7231 17013
rect 6162 16968 7231 16979
rect 7265 16984 7323 17055
rect 5425 16877 5443 16911
rect 5477 16877 6075 16911
rect 6109 16877 6127 16911
rect 5425 16837 6127 16877
rect 5425 16767 5763 16837
rect 5425 16733 5503 16767
rect 5537 16733 5606 16767
rect 5640 16733 5709 16767
rect 5743 16733 5763 16767
rect 5797 16769 5817 16803
rect 5851 16769 5916 16803
rect 5950 16769 6015 16803
rect 6049 16769 6127 16803
rect 5797 16699 6127 16769
rect 6480 16767 6550 16968
rect 7265 16950 7277 16984
rect 7311 16950 7323 16984
rect 7265 16891 7323 16950
rect 7265 16857 7277 16891
rect 7311 16857 7323 16891
rect 7265 16822 7323 16857
rect 7449 17013 7967 17055
rect 7449 16979 7467 17013
rect 7501 16979 7915 17013
rect 7949 16979 7967 17013
rect 7449 16911 7967 16979
rect 8002 17013 9071 17055
rect 8002 16979 8019 17013
rect 8053 16979 9019 17013
rect 9053 16979 9071 17013
rect 8002 16968 9071 16979
rect 9106 17013 10175 17055
rect 9106 16979 9123 17013
rect 9157 16979 10123 17013
rect 10157 16979 10175 17013
rect 9106 16968 10175 16979
rect 10210 17013 11279 17055
rect 10210 16979 10227 17013
rect 10261 16979 11227 17013
rect 11261 16979 11279 17013
rect 10210 16968 11279 16979
rect 11314 17013 12383 17055
rect 11314 16979 11331 17013
rect 11365 16979 12331 17013
rect 12365 16979 12383 17013
rect 11314 16968 12383 16979
rect 12417 16984 12475 17055
rect 7449 16877 7467 16911
rect 7501 16877 7915 16911
rect 7949 16877 7967 16911
rect 7449 16837 7967 16877
rect 6480 16733 6499 16767
rect 6533 16733 6550 16767
rect 6480 16718 6550 16733
rect 6846 16803 6914 16820
rect 6846 16769 6863 16803
rect 6897 16769 6914 16803
rect 4965 16642 5207 16695
rect 4965 16608 4983 16642
rect 5017 16608 5155 16642
rect 5189 16608 5207 16642
rect 4965 16545 5207 16608
rect 5425 16640 6127 16699
rect 6846 16654 6914 16769
rect 7449 16767 7691 16837
rect 7449 16733 7527 16767
rect 7561 16733 7637 16767
rect 7671 16733 7691 16767
rect 7725 16769 7745 16803
rect 7779 16769 7855 16803
rect 7889 16769 7967 16803
rect 7725 16699 7967 16769
rect 8320 16767 8390 16968
rect 8320 16733 8339 16767
rect 8373 16733 8390 16767
rect 8320 16718 8390 16733
rect 8686 16803 8754 16820
rect 8686 16769 8703 16803
rect 8737 16769 8754 16803
rect 7265 16673 7323 16690
rect 5425 16606 5443 16640
rect 5477 16606 6075 16640
rect 6109 16606 6127 16640
rect 5425 16545 6127 16606
rect 6162 16640 7231 16654
rect 6162 16606 6179 16640
rect 6213 16606 7179 16640
rect 7213 16606 7231 16640
rect 6162 16545 7231 16606
rect 7265 16639 7277 16673
rect 7311 16639 7323 16673
rect 7265 16545 7323 16639
rect 7449 16640 7967 16699
rect 8686 16654 8754 16769
rect 9424 16767 9494 16968
rect 9424 16733 9443 16767
rect 9477 16733 9494 16767
rect 9424 16718 9494 16733
rect 9790 16803 9858 16820
rect 9790 16769 9807 16803
rect 9841 16769 9858 16803
rect 9790 16654 9858 16769
rect 10528 16767 10598 16968
rect 10528 16733 10547 16767
rect 10581 16733 10598 16767
rect 10528 16718 10598 16733
rect 10894 16803 10962 16820
rect 10894 16769 10911 16803
rect 10945 16769 10962 16803
rect 10894 16654 10962 16769
rect 11632 16767 11702 16968
rect 12417 16950 12429 16984
rect 12463 16950 12475 16984
rect 12417 16891 12475 16950
rect 12417 16857 12429 16891
rect 12463 16857 12475 16891
rect 12417 16822 12475 16857
rect 12601 17013 13119 17055
rect 12601 16979 12619 17013
rect 12653 16979 13067 17013
rect 13101 16979 13119 17013
rect 12601 16911 13119 16979
rect 13154 17013 14223 17055
rect 13154 16979 13171 17013
rect 13205 16979 14171 17013
rect 14205 16979 14223 17013
rect 13154 16968 14223 16979
rect 14258 17013 15327 17055
rect 14258 16979 14275 17013
rect 14309 16979 15275 17013
rect 15309 16979 15327 17013
rect 14258 16968 15327 16979
rect 15362 17013 16431 17055
rect 15362 16979 15379 17013
rect 15413 16979 16379 17013
rect 16413 16979 16431 17013
rect 15362 16968 16431 16979
rect 16466 17013 17535 17055
rect 16466 16979 16483 17013
rect 16517 16979 17483 17013
rect 17517 16979 17535 17013
rect 16466 16968 17535 16979
rect 17569 16984 17627 17055
rect 12601 16877 12619 16911
rect 12653 16877 13067 16911
rect 13101 16877 13119 16911
rect 12601 16837 13119 16877
rect 11632 16733 11651 16767
rect 11685 16733 11702 16767
rect 11632 16718 11702 16733
rect 11998 16803 12066 16820
rect 11998 16769 12015 16803
rect 12049 16769 12066 16803
rect 11998 16654 12066 16769
rect 12601 16767 12843 16837
rect 12601 16733 12679 16767
rect 12713 16733 12789 16767
rect 12823 16733 12843 16767
rect 12877 16769 12897 16803
rect 12931 16769 13007 16803
rect 13041 16769 13119 16803
rect 12877 16699 13119 16769
rect 13472 16767 13542 16968
rect 13472 16733 13491 16767
rect 13525 16733 13542 16767
rect 13472 16718 13542 16733
rect 13838 16803 13906 16820
rect 13838 16769 13855 16803
rect 13889 16769 13906 16803
rect 12417 16673 12475 16690
rect 7449 16606 7467 16640
rect 7501 16606 7915 16640
rect 7949 16606 7967 16640
rect 7449 16545 7967 16606
rect 8002 16640 9071 16654
rect 8002 16606 8019 16640
rect 8053 16606 9019 16640
rect 9053 16606 9071 16640
rect 8002 16545 9071 16606
rect 9106 16640 10175 16654
rect 9106 16606 9123 16640
rect 9157 16606 10123 16640
rect 10157 16606 10175 16640
rect 9106 16545 10175 16606
rect 10210 16640 11279 16654
rect 10210 16606 10227 16640
rect 10261 16606 11227 16640
rect 11261 16606 11279 16640
rect 10210 16545 11279 16606
rect 11314 16640 12383 16654
rect 11314 16606 11331 16640
rect 11365 16606 12331 16640
rect 12365 16606 12383 16640
rect 11314 16545 12383 16606
rect 12417 16639 12429 16673
rect 12463 16639 12475 16673
rect 12417 16545 12475 16639
rect 12601 16640 13119 16699
rect 13838 16654 13906 16769
rect 14576 16767 14646 16968
rect 14576 16733 14595 16767
rect 14629 16733 14646 16767
rect 14576 16718 14646 16733
rect 14942 16803 15010 16820
rect 14942 16769 14959 16803
rect 14993 16769 15010 16803
rect 14942 16654 15010 16769
rect 15680 16767 15750 16968
rect 15680 16733 15699 16767
rect 15733 16733 15750 16767
rect 15680 16718 15750 16733
rect 16046 16803 16114 16820
rect 16046 16769 16063 16803
rect 16097 16769 16114 16803
rect 16046 16654 16114 16769
rect 16784 16767 16854 16968
rect 17569 16950 17581 16984
rect 17615 16950 17627 16984
rect 17754 17013 18823 17055
rect 17754 16979 17771 17013
rect 17805 16979 18771 17013
rect 18805 16979 18823 17013
rect 17754 16968 18823 16979
rect 18858 17013 19927 17055
rect 18858 16979 18875 17013
rect 18909 16979 19875 17013
rect 19909 16979 19927 17013
rect 18858 16968 19927 16979
rect 19961 17013 20203 17055
rect 19961 16979 19979 17013
rect 20013 16979 20151 17013
rect 20185 16979 20203 17013
rect 17569 16891 17627 16950
rect 17569 16857 17581 16891
rect 17615 16857 17627 16891
rect 17569 16822 17627 16857
rect 16784 16733 16803 16767
rect 16837 16733 16854 16767
rect 16784 16718 16854 16733
rect 17150 16803 17218 16820
rect 17150 16769 17167 16803
rect 17201 16769 17218 16803
rect 17150 16654 17218 16769
rect 18072 16767 18142 16968
rect 18072 16733 18091 16767
rect 18125 16733 18142 16767
rect 18072 16718 18142 16733
rect 18438 16803 18506 16820
rect 18438 16769 18455 16803
rect 18489 16769 18506 16803
rect 17569 16673 17627 16690
rect 12601 16606 12619 16640
rect 12653 16606 13067 16640
rect 13101 16606 13119 16640
rect 12601 16545 13119 16606
rect 13154 16640 14223 16654
rect 13154 16606 13171 16640
rect 13205 16606 14171 16640
rect 14205 16606 14223 16640
rect 13154 16545 14223 16606
rect 14258 16640 15327 16654
rect 14258 16606 14275 16640
rect 14309 16606 15275 16640
rect 15309 16606 15327 16640
rect 14258 16545 15327 16606
rect 15362 16640 16431 16654
rect 15362 16606 15379 16640
rect 15413 16606 16379 16640
rect 16413 16606 16431 16640
rect 15362 16545 16431 16606
rect 16466 16640 17535 16654
rect 16466 16606 16483 16640
rect 16517 16606 17483 16640
rect 17517 16606 17535 16640
rect 16466 16545 17535 16606
rect 17569 16639 17581 16673
rect 17615 16639 17627 16673
rect 18438 16654 18506 16769
rect 19176 16767 19246 16968
rect 19961 16918 20203 16979
rect 19961 16884 19979 16918
rect 20013 16884 20151 16918
rect 20185 16884 20203 16918
rect 19961 16837 20203 16884
rect 19176 16733 19195 16767
rect 19229 16733 19246 16767
rect 19176 16718 19246 16733
rect 19542 16803 19610 16820
rect 19542 16769 19559 16803
rect 19593 16769 19610 16803
rect 19542 16654 19610 16769
rect 19961 16763 20065 16837
rect 19961 16729 20011 16763
rect 20045 16729 20065 16763
rect 20099 16769 20119 16803
rect 20153 16769 20203 16803
rect 20099 16695 20203 16769
rect 17569 16545 17627 16639
rect 17754 16640 18823 16654
rect 17754 16606 17771 16640
rect 17805 16606 18771 16640
rect 18805 16606 18823 16640
rect 17754 16545 18823 16606
rect 18858 16640 19927 16654
rect 18858 16606 18875 16640
rect 18909 16606 19875 16640
rect 19909 16606 19927 16640
rect 18858 16545 19927 16606
rect 19961 16642 20203 16695
rect 19961 16608 19979 16642
rect 20013 16608 20151 16642
rect 20185 16608 20203 16642
rect 19961 16545 20203 16608
rect 4948 16511 4977 16545
rect 5011 16511 5069 16545
rect 5103 16511 5161 16545
rect 5195 16511 5253 16545
rect 5287 16511 5345 16545
rect 5379 16511 5437 16545
rect 5471 16511 5529 16545
rect 5563 16511 5621 16545
rect 5655 16511 5713 16545
rect 5747 16511 5805 16545
rect 5839 16511 5897 16545
rect 5931 16511 5989 16545
rect 6023 16511 6081 16545
rect 6115 16511 6173 16545
rect 6207 16511 6265 16545
rect 6299 16511 6357 16545
rect 6391 16511 6449 16545
rect 6483 16511 6541 16545
rect 6575 16511 6633 16545
rect 6667 16511 6725 16545
rect 6759 16511 6817 16545
rect 6851 16511 6909 16545
rect 6943 16511 7001 16545
rect 7035 16511 7093 16545
rect 7127 16511 7185 16545
rect 7219 16511 7277 16545
rect 7311 16511 7369 16545
rect 7403 16511 7461 16545
rect 7495 16511 7553 16545
rect 7587 16511 7645 16545
rect 7679 16511 7737 16545
rect 7771 16511 7829 16545
rect 7863 16511 7921 16545
rect 7955 16511 8013 16545
rect 8047 16511 8105 16545
rect 8139 16511 8197 16545
rect 8231 16511 8289 16545
rect 8323 16511 8381 16545
rect 8415 16511 8473 16545
rect 8507 16511 8565 16545
rect 8599 16511 8657 16545
rect 8691 16511 8749 16545
rect 8783 16511 8841 16545
rect 8875 16511 8933 16545
rect 8967 16511 9025 16545
rect 9059 16511 9117 16545
rect 9151 16511 9209 16545
rect 9243 16511 9301 16545
rect 9335 16511 9393 16545
rect 9427 16511 9485 16545
rect 9519 16511 9577 16545
rect 9611 16511 9669 16545
rect 9703 16511 9761 16545
rect 9795 16511 9853 16545
rect 9887 16511 9945 16545
rect 9979 16511 10037 16545
rect 10071 16511 10129 16545
rect 10163 16511 10221 16545
rect 10255 16511 10313 16545
rect 10347 16511 10405 16545
rect 10439 16511 10497 16545
rect 10531 16511 10589 16545
rect 10623 16511 10681 16545
rect 10715 16511 10773 16545
rect 10807 16511 10865 16545
rect 10899 16511 10957 16545
rect 10991 16511 11049 16545
rect 11083 16511 11141 16545
rect 11175 16511 11233 16545
rect 11267 16511 11325 16545
rect 11359 16511 11417 16545
rect 11451 16511 11509 16545
rect 11543 16511 11601 16545
rect 11635 16511 11693 16545
rect 11727 16511 11785 16545
rect 11819 16511 11877 16545
rect 11911 16511 11969 16545
rect 12003 16511 12061 16545
rect 12095 16511 12153 16545
rect 12187 16511 12245 16545
rect 12279 16511 12337 16545
rect 12371 16511 12429 16545
rect 12463 16511 12521 16545
rect 12555 16511 12613 16545
rect 12647 16511 12705 16545
rect 12739 16511 12797 16545
rect 12831 16511 12889 16545
rect 12923 16511 12981 16545
rect 13015 16511 13073 16545
rect 13107 16511 13165 16545
rect 13199 16511 13257 16545
rect 13291 16511 13349 16545
rect 13383 16511 13441 16545
rect 13475 16511 13533 16545
rect 13567 16511 13625 16545
rect 13659 16511 13717 16545
rect 13751 16511 13809 16545
rect 13843 16511 13901 16545
rect 13935 16511 13993 16545
rect 14027 16511 14085 16545
rect 14119 16511 14177 16545
rect 14211 16511 14269 16545
rect 14303 16511 14361 16545
rect 14395 16511 14453 16545
rect 14487 16511 14545 16545
rect 14579 16511 14637 16545
rect 14671 16511 14729 16545
rect 14763 16511 14821 16545
rect 14855 16511 14913 16545
rect 14947 16511 15005 16545
rect 15039 16511 15097 16545
rect 15131 16511 15189 16545
rect 15223 16511 15281 16545
rect 15315 16511 15373 16545
rect 15407 16511 15465 16545
rect 15499 16511 15557 16545
rect 15591 16511 15649 16545
rect 15683 16511 15741 16545
rect 15775 16511 15833 16545
rect 15867 16511 15925 16545
rect 15959 16511 16017 16545
rect 16051 16511 16109 16545
rect 16143 16511 16201 16545
rect 16235 16511 16293 16545
rect 16327 16511 16385 16545
rect 16419 16511 16477 16545
rect 16511 16511 16569 16545
rect 16603 16511 16661 16545
rect 16695 16511 16753 16545
rect 16787 16511 16845 16545
rect 16879 16511 16937 16545
rect 16971 16511 17029 16545
rect 17063 16511 17121 16545
rect 17155 16511 17213 16545
rect 17247 16511 17305 16545
rect 17339 16511 17397 16545
rect 17431 16511 17489 16545
rect 17523 16511 17581 16545
rect 17615 16511 17673 16545
rect 17707 16511 17765 16545
rect 17799 16511 17857 16545
rect 17891 16511 17949 16545
rect 17983 16511 18041 16545
rect 18075 16511 18133 16545
rect 18167 16511 18225 16545
rect 18259 16511 18317 16545
rect 18351 16511 18409 16545
rect 18443 16511 18501 16545
rect 18535 16511 18593 16545
rect 18627 16511 18685 16545
rect 18719 16511 18777 16545
rect 18811 16511 18869 16545
rect 18903 16511 18961 16545
rect 18995 16511 19053 16545
rect 19087 16511 19145 16545
rect 19179 16511 19237 16545
rect 19271 16511 19329 16545
rect 19363 16511 19421 16545
rect 19455 16511 19513 16545
rect 19547 16511 19605 16545
rect 19639 16511 19697 16545
rect 19731 16511 19789 16545
rect 19823 16511 19881 16545
rect 19915 16511 19973 16545
rect 20007 16511 20065 16545
rect 20099 16511 20157 16545
rect 20191 16511 20220 16545
rect 4965 16448 5207 16511
rect 4965 16414 4983 16448
rect 5017 16414 5155 16448
rect 5189 16414 5207 16448
rect 4965 16361 5207 16414
rect 5426 16450 6495 16511
rect 5426 16416 5443 16450
rect 5477 16416 6443 16450
rect 6477 16416 6495 16450
rect 5426 16402 6495 16416
rect 6530 16450 7599 16511
rect 6530 16416 6547 16450
rect 6581 16416 7547 16450
rect 7581 16416 7599 16450
rect 6530 16402 7599 16416
rect 7634 16450 8703 16511
rect 7634 16416 7651 16450
rect 7685 16416 8651 16450
rect 8685 16416 8703 16450
rect 7634 16402 8703 16416
rect 8738 16450 9807 16511
rect 8738 16416 8755 16450
rect 8789 16416 9755 16450
rect 9789 16416 9807 16450
rect 8738 16402 9807 16416
rect 9841 16417 9899 16511
rect 4965 16287 5069 16361
rect 4965 16253 5015 16287
rect 5049 16253 5069 16287
rect 5103 16293 5123 16327
rect 5157 16293 5207 16327
rect 5103 16219 5207 16293
rect 4965 16172 5207 16219
rect 4965 16138 4983 16172
rect 5017 16138 5155 16172
rect 5189 16138 5207 16172
rect 4965 16077 5207 16138
rect 5744 16323 5814 16338
rect 5744 16289 5763 16323
rect 5797 16289 5814 16323
rect 5744 16088 5814 16289
rect 6110 16287 6178 16402
rect 6110 16253 6127 16287
rect 6161 16253 6178 16287
rect 6110 16236 6178 16253
rect 6848 16323 6918 16338
rect 6848 16289 6867 16323
rect 6901 16289 6918 16323
rect 6848 16088 6918 16289
rect 7214 16287 7282 16402
rect 7214 16253 7231 16287
rect 7265 16253 7282 16287
rect 7214 16236 7282 16253
rect 7952 16323 8022 16338
rect 7952 16289 7971 16323
rect 8005 16289 8022 16323
rect 7952 16088 8022 16289
rect 8318 16287 8386 16402
rect 8318 16253 8335 16287
rect 8369 16253 8386 16287
rect 8318 16236 8386 16253
rect 9056 16323 9126 16338
rect 9056 16289 9075 16323
rect 9109 16289 9126 16323
rect 9056 16088 9126 16289
rect 9422 16287 9490 16402
rect 9841 16383 9853 16417
rect 9887 16383 9899 16417
rect 9841 16366 9899 16383
rect 10025 16450 10543 16511
rect 10025 16416 10043 16450
rect 10077 16416 10491 16450
rect 10525 16416 10543 16450
rect 10025 16357 10543 16416
rect 10578 16450 11647 16511
rect 10578 16416 10595 16450
rect 10629 16416 11595 16450
rect 11629 16416 11647 16450
rect 10578 16402 11647 16416
rect 11682 16450 12751 16511
rect 11682 16416 11699 16450
rect 11733 16416 12699 16450
rect 12733 16416 12751 16450
rect 11682 16402 12751 16416
rect 12786 16450 13855 16511
rect 12786 16416 12803 16450
rect 12837 16416 13803 16450
rect 13837 16416 13855 16450
rect 12786 16402 13855 16416
rect 13890 16450 14959 16511
rect 13890 16416 13907 16450
rect 13941 16416 14907 16450
rect 14941 16416 14959 16450
rect 13890 16402 14959 16416
rect 14993 16417 15051 16511
rect 9422 16253 9439 16287
rect 9473 16253 9490 16287
rect 9422 16236 9490 16253
rect 10025 16289 10103 16323
rect 10137 16289 10213 16323
rect 10247 16289 10267 16323
rect 9841 16199 9899 16234
rect 9841 16165 9853 16199
rect 9887 16165 9899 16199
rect 9841 16106 9899 16165
rect 4965 16043 4983 16077
rect 5017 16043 5155 16077
rect 5189 16043 5207 16077
rect 4965 16001 5207 16043
rect 5426 16077 6495 16088
rect 5426 16043 5443 16077
rect 5477 16043 6443 16077
rect 6477 16043 6495 16077
rect 5426 16001 6495 16043
rect 6530 16077 7599 16088
rect 6530 16043 6547 16077
rect 6581 16043 7547 16077
rect 7581 16043 7599 16077
rect 6530 16001 7599 16043
rect 7634 16077 8703 16088
rect 7634 16043 7651 16077
rect 7685 16043 8651 16077
rect 8685 16043 8703 16077
rect 7634 16001 8703 16043
rect 8738 16077 9807 16088
rect 8738 16043 8755 16077
rect 8789 16043 9755 16077
rect 9789 16043 9807 16077
rect 8738 16001 9807 16043
rect 9841 16072 9853 16106
rect 9887 16072 9899 16106
rect 9841 16001 9899 16072
rect 10025 16219 10267 16289
rect 10301 16287 10543 16357
rect 10301 16253 10321 16287
rect 10355 16253 10431 16287
rect 10465 16253 10543 16287
rect 10896 16323 10966 16338
rect 10896 16289 10915 16323
rect 10949 16289 10966 16323
rect 10025 16179 10543 16219
rect 10025 16145 10043 16179
rect 10077 16145 10491 16179
rect 10525 16145 10543 16179
rect 10025 16077 10543 16145
rect 10896 16088 10966 16289
rect 11262 16287 11330 16402
rect 11262 16253 11279 16287
rect 11313 16253 11330 16287
rect 11262 16236 11330 16253
rect 12000 16323 12070 16338
rect 12000 16289 12019 16323
rect 12053 16289 12070 16323
rect 12000 16088 12070 16289
rect 12366 16287 12434 16402
rect 12366 16253 12383 16287
rect 12417 16253 12434 16287
rect 12366 16236 12434 16253
rect 13104 16323 13174 16338
rect 13104 16289 13123 16323
rect 13157 16289 13174 16323
rect 13104 16088 13174 16289
rect 13470 16287 13538 16402
rect 13470 16253 13487 16287
rect 13521 16253 13538 16287
rect 13470 16236 13538 16253
rect 14208 16323 14278 16338
rect 14208 16289 14227 16323
rect 14261 16289 14278 16323
rect 14208 16088 14278 16289
rect 14574 16287 14642 16402
rect 14993 16383 15005 16417
rect 15039 16383 15051 16417
rect 14993 16366 15051 16383
rect 15177 16443 15511 16511
rect 15177 16409 15195 16443
rect 15229 16409 15459 16443
rect 15493 16409 15511 16443
rect 15177 16357 15511 16409
rect 15546 16450 16615 16511
rect 15546 16416 15563 16450
rect 15597 16416 16563 16450
rect 16597 16416 16615 16450
rect 15546 16402 16615 16416
rect 16650 16450 17719 16511
rect 16650 16416 16667 16450
rect 16701 16416 17667 16450
rect 17701 16416 17719 16450
rect 16650 16402 17719 16416
rect 17754 16450 18823 16511
rect 17754 16416 17771 16450
rect 17805 16416 18771 16450
rect 18805 16416 18823 16450
rect 17754 16402 18823 16416
rect 18858 16450 19927 16511
rect 18858 16416 18875 16450
rect 18909 16416 19875 16450
rect 19909 16416 19927 16450
rect 18858 16402 19927 16416
rect 19961 16448 20203 16511
rect 19961 16414 19979 16448
rect 20013 16414 20151 16448
rect 20185 16414 20203 16448
rect 14574 16253 14591 16287
rect 14625 16253 14642 16287
rect 14574 16236 14642 16253
rect 15177 16289 15197 16323
rect 15231 16289 15327 16323
rect 14993 16199 15051 16234
rect 14993 16165 15005 16199
rect 15039 16165 15051 16199
rect 14993 16106 15051 16165
rect 10025 16043 10043 16077
rect 10077 16043 10491 16077
rect 10525 16043 10543 16077
rect 10025 16001 10543 16043
rect 10578 16077 11647 16088
rect 10578 16043 10595 16077
rect 10629 16043 11595 16077
rect 11629 16043 11647 16077
rect 10578 16001 11647 16043
rect 11682 16077 12751 16088
rect 11682 16043 11699 16077
rect 11733 16043 12699 16077
rect 12733 16043 12751 16077
rect 11682 16001 12751 16043
rect 12786 16077 13855 16088
rect 12786 16043 12803 16077
rect 12837 16043 13803 16077
rect 13837 16043 13855 16077
rect 12786 16001 13855 16043
rect 13890 16077 14959 16088
rect 13890 16043 13907 16077
rect 13941 16043 14907 16077
rect 14941 16043 14959 16077
rect 13890 16001 14959 16043
rect 14993 16072 15005 16106
rect 15039 16072 15051 16106
rect 14993 16001 15051 16072
rect 15177 16219 15327 16289
rect 15361 16287 15511 16357
rect 15361 16253 15457 16287
rect 15491 16253 15511 16287
rect 15864 16323 15934 16338
rect 15864 16289 15883 16323
rect 15917 16289 15934 16323
rect 15177 16179 15511 16219
rect 15177 16145 15195 16179
rect 15229 16145 15459 16179
rect 15493 16145 15511 16179
rect 15177 16077 15511 16145
rect 15864 16088 15934 16289
rect 16230 16287 16298 16402
rect 16230 16253 16247 16287
rect 16281 16253 16298 16287
rect 16230 16236 16298 16253
rect 16968 16323 17038 16338
rect 16968 16289 16987 16323
rect 17021 16289 17038 16323
rect 16968 16088 17038 16289
rect 17334 16287 17402 16402
rect 17334 16253 17351 16287
rect 17385 16253 17402 16287
rect 17334 16236 17402 16253
rect 18072 16323 18142 16338
rect 18072 16289 18091 16323
rect 18125 16289 18142 16323
rect 18072 16088 18142 16289
rect 18438 16287 18506 16402
rect 18438 16253 18455 16287
rect 18489 16253 18506 16287
rect 18438 16236 18506 16253
rect 19176 16323 19246 16338
rect 19176 16289 19195 16323
rect 19229 16289 19246 16323
rect 19176 16088 19246 16289
rect 19542 16287 19610 16402
rect 19961 16361 20203 16414
rect 19542 16253 19559 16287
rect 19593 16253 19610 16287
rect 19542 16236 19610 16253
rect 19961 16293 20011 16327
rect 20045 16293 20065 16327
rect 19961 16219 20065 16293
rect 20099 16287 20203 16361
rect 20099 16253 20119 16287
rect 20153 16253 20203 16287
rect 19961 16172 20203 16219
rect 19961 16138 19979 16172
rect 20013 16138 20151 16172
rect 20185 16138 20203 16172
rect 15177 16043 15195 16077
rect 15229 16043 15459 16077
rect 15493 16043 15511 16077
rect 15177 16001 15511 16043
rect 15546 16077 16615 16088
rect 15546 16043 15563 16077
rect 15597 16043 16563 16077
rect 16597 16043 16615 16077
rect 15546 16001 16615 16043
rect 16650 16077 17719 16088
rect 16650 16043 16667 16077
rect 16701 16043 17667 16077
rect 17701 16043 17719 16077
rect 16650 16001 17719 16043
rect 17754 16077 18823 16088
rect 17754 16043 17771 16077
rect 17805 16043 18771 16077
rect 18805 16043 18823 16077
rect 17754 16001 18823 16043
rect 18858 16077 19927 16088
rect 18858 16043 18875 16077
rect 18909 16043 19875 16077
rect 19909 16043 19927 16077
rect 18858 16001 19927 16043
rect 19961 16077 20203 16138
rect 19961 16043 19979 16077
rect 20013 16043 20151 16077
rect 20185 16043 20203 16077
rect 19961 16001 20203 16043
rect 4948 15967 4977 16001
rect 5011 15967 5069 16001
rect 5103 15967 5161 16001
rect 5195 15967 5253 16001
rect 5287 15967 5345 16001
rect 5379 15967 5437 16001
rect 5471 15967 5529 16001
rect 5563 15967 5621 16001
rect 5655 15967 5713 16001
rect 5747 15967 5805 16001
rect 5839 15967 5897 16001
rect 5931 15967 5989 16001
rect 6023 15967 6081 16001
rect 6115 15967 6173 16001
rect 6207 15967 6265 16001
rect 6299 15967 6357 16001
rect 6391 15967 6449 16001
rect 6483 15967 6541 16001
rect 6575 15967 6633 16001
rect 6667 15967 6725 16001
rect 6759 15967 6817 16001
rect 6851 15967 6909 16001
rect 6943 15967 7001 16001
rect 7035 15967 7093 16001
rect 7127 15967 7185 16001
rect 7219 15967 7277 16001
rect 7311 15967 7369 16001
rect 7403 15967 7461 16001
rect 7495 15967 7553 16001
rect 7587 15967 7645 16001
rect 7679 15967 7737 16001
rect 7771 15967 7829 16001
rect 7863 15967 7921 16001
rect 7955 15967 8013 16001
rect 8047 15967 8105 16001
rect 8139 15967 8197 16001
rect 8231 15967 8289 16001
rect 8323 15967 8381 16001
rect 8415 15967 8473 16001
rect 8507 15967 8565 16001
rect 8599 15967 8657 16001
rect 8691 15967 8749 16001
rect 8783 15967 8841 16001
rect 8875 15967 8933 16001
rect 8967 15967 9025 16001
rect 9059 15967 9117 16001
rect 9151 15967 9209 16001
rect 9243 15967 9301 16001
rect 9335 15967 9393 16001
rect 9427 15967 9485 16001
rect 9519 15967 9577 16001
rect 9611 15967 9669 16001
rect 9703 15967 9761 16001
rect 9795 15967 9853 16001
rect 9887 15967 9945 16001
rect 9979 15967 10037 16001
rect 10071 15967 10129 16001
rect 10163 15967 10221 16001
rect 10255 15967 10313 16001
rect 10347 15967 10405 16001
rect 10439 15967 10497 16001
rect 10531 15967 10589 16001
rect 10623 15967 10681 16001
rect 10715 15967 10773 16001
rect 10807 15967 10865 16001
rect 10899 15967 10957 16001
rect 10991 15967 11049 16001
rect 11083 15967 11141 16001
rect 11175 15967 11233 16001
rect 11267 15967 11325 16001
rect 11359 15967 11417 16001
rect 11451 15967 11509 16001
rect 11543 15967 11601 16001
rect 11635 15967 11693 16001
rect 11727 15967 11785 16001
rect 11819 15967 11877 16001
rect 11911 15967 11969 16001
rect 12003 15967 12061 16001
rect 12095 15967 12153 16001
rect 12187 15967 12245 16001
rect 12279 15967 12337 16001
rect 12371 15967 12429 16001
rect 12463 15967 12521 16001
rect 12555 15967 12613 16001
rect 12647 15967 12705 16001
rect 12739 15967 12797 16001
rect 12831 15967 12889 16001
rect 12923 15967 12981 16001
rect 13015 15967 13073 16001
rect 13107 15967 13165 16001
rect 13199 15967 13257 16001
rect 13291 15967 13349 16001
rect 13383 15967 13441 16001
rect 13475 15967 13533 16001
rect 13567 15967 13625 16001
rect 13659 15967 13717 16001
rect 13751 15967 13809 16001
rect 13843 15967 13901 16001
rect 13935 15967 13993 16001
rect 14027 15967 14085 16001
rect 14119 15967 14177 16001
rect 14211 15967 14269 16001
rect 14303 15967 14361 16001
rect 14395 15967 14453 16001
rect 14487 15967 14545 16001
rect 14579 15967 14637 16001
rect 14671 15967 14729 16001
rect 14763 15967 14821 16001
rect 14855 15967 14913 16001
rect 14947 15967 15005 16001
rect 15039 15967 15097 16001
rect 15131 15967 15189 16001
rect 15223 15967 15281 16001
rect 15315 15967 15373 16001
rect 15407 15967 15465 16001
rect 15499 15967 15557 16001
rect 15591 15967 15649 16001
rect 15683 15967 15741 16001
rect 15775 15967 15833 16001
rect 15867 15967 15925 16001
rect 15959 15967 16017 16001
rect 16051 15967 16109 16001
rect 16143 15967 16201 16001
rect 16235 15967 16293 16001
rect 16327 15967 16385 16001
rect 16419 15967 16477 16001
rect 16511 15967 16569 16001
rect 16603 15967 16661 16001
rect 16695 15967 16753 16001
rect 16787 15967 16845 16001
rect 16879 15967 16937 16001
rect 16971 15967 17029 16001
rect 17063 15967 17121 16001
rect 17155 15967 17213 16001
rect 17247 15967 17305 16001
rect 17339 15967 17397 16001
rect 17431 15967 17489 16001
rect 17523 15967 17581 16001
rect 17615 15967 17673 16001
rect 17707 15967 17765 16001
rect 17799 15967 17857 16001
rect 17891 15967 17949 16001
rect 17983 15967 18041 16001
rect 18075 15967 18133 16001
rect 18167 15967 18225 16001
rect 18259 15967 18317 16001
rect 18351 15967 18409 16001
rect 18443 15967 18501 16001
rect 18535 15967 18593 16001
rect 18627 15967 18685 16001
rect 18719 15967 18777 16001
rect 18811 15967 18869 16001
rect 18903 15967 18961 16001
rect 18995 15967 19053 16001
rect 19087 15967 19145 16001
rect 19179 15967 19237 16001
rect 19271 15967 19329 16001
rect 19363 15967 19421 16001
rect 19455 15967 19513 16001
rect 19547 15967 19605 16001
rect 19639 15967 19697 16001
rect 19731 15967 19789 16001
rect 19823 15967 19881 16001
rect 19915 15967 19973 16001
rect 20007 15967 20065 16001
rect 20099 15967 20157 16001
rect 20191 15967 20220 16001
rect 4965 15925 5207 15967
rect 4965 15891 4983 15925
rect 5017 15891 5155 15925
rect 5189 15891 5207 15925
rect 4965 15830 5207 15891
rect 4965 15796 4983 15830
rect 5017 15796 5155 15830
rect 5189 15796 5207 15830
rect 4965 15749 5207 15796
rect 4965 15681 5015 15715
rect 5049 15681 5069 15715
rect 4965 15607 5069 15681
rect 5103 15675 5207 15749
rect 5103 15641 5123 15675
rect 5157 15641 5207 15675
rect 5425 15925 6127 15967
rect 5425 15891 5443 15925
rect 5477 15891 6075 15925
rect 6109 15891 6127 15925
rect 5425 15823 6127 15891
rect 6162 15925 7231 15967
rect 6162 15891 6179 15925
rect 6213 15891 7179 15925
rect 7213 15891 7231 15925
rect 6162 15880 7231 15891
rect 7265 15896 7323 15967
rect 5425 15789 5443 15823
rect 5477 15789 6075 15823
rect 6109 15789 6127 15823
rect 5425 15749 6127 15789
rect 5425 15679 5763 15749
rect 5425 15645 5503 15679
rect 5537 15645 5606 15679
rect 5640 15645 5709 15679
rect 5743 15645 5763 15679
rect 5797 15681 5817 15715
rect 5851 15681 5916 15715
rect 5950 15681 6015 15715
rect 6049 15681 6127 15715
rect 5797 15611 6127 15681
rect 6480 15679 6550 15880
rect 7265 15862 7277 15896
rect 7311 15862 7323 15896
rect 7265 15803 7323 15862
rect 7265 15769 7277 15803
rect 7311 15769 7323 15803
rect 7265 15734 7323 15769
rect 7449 15925 7967 15967
rect 7449 15891 7467 15925
rect 7501 15891 7915 15925
rect 7949 15891 7967 15925
rect 7449 15823 7967 15891
rect 8002 15925 9071 15967
rect 8002 15891 8019 15925
rect 8053 15891 9019 15925
rect 9053 15891 9071 15925
rect 8002 15880 9071 15891
rect 9106 15925 10175 15967
rect 9106 15891 9123 15925
rect 9157 15891 10123 15925
rect 10157 15891 10175 15925
rect 9106 15880 10175 15891
rect 10210 15925 11279 15967
rect 10210 15891 10227 15925
rect 10261 15891 11227 15925
rect 11261 15891 11279 15925
rect 10210 15880 11279 15891
rect 11314 15925 12383 15967
rect 11314 15891 11331 15925
rect 11365 15891 12331 15925
rect 12365 15891 12383 15925
rect 11314 15880 12383 15891
rect 12417 15896 12475 15967
rect 7449 15789 7467 15823
rect 7501 15789 7915 15823
rect 7949 15789 7967 15823
rect 7449 15749 7967 15789
rect 6480 15645 6499 15679
rect 6533 15645 6550 15679
rect 6480 15630 6550 15645
rect 6846 15715 6914 15732
rect 6846 15681 6863 15715
rect 6897 15681 6914 15715
rect 4965 15554 5207 15607
rect 4965 15520 4983 15554
rect 5017 15520 5155 15554
rect 5189 15520 5207 15554
rect 4965 15457 5207 15520
rect 5425 15552 6127 15611
rect 6846 15566 6914 15681
rect 7449 15679 7691 15749
rect 7449 15645 7527 15679
rect 7561 15645 7637 15679
rect 7671 15645 7691 15679
rect 7725 15681 7745 15715
rect 7779 15681 7855 15715
rect 7889 15681 7967 15715
rect 7725 15611 7967 15681
rect 8320 15679 8390 15880
rect 8320 15645 8339 15679
rect 8373 15645 8390 15679
rect 8320 15630 8390 15645
rect 8686 15715 8754 15732
rect 8686 15681 8703 15715
rect 8737 15681 8754 15715
rect 7265 15585 7323 15602
rect 5425 15518 5443 15552
rect 5477 15518 6075 15552
rect 6109 15518 6127 15552
rect 5425 15457 6127 15518
rect 6162 15552 7231 15566
rect 6162 15518 6179 15552
rect 6213 15518 7179 15552
rect 7213 15518 7231 15552
rect 6162 15457 7231 15518
rect 7265 15551 7277 15585
rect 7311 15551 7323 15585
rect 7265 15457 7323 15551
rect 7449 15552 7967 15611
rect 8686 15566 8754 15681
rect 9424 15679 9494 15880
rect 9424 15645 9443 15679
rect 9477 15645 9494 15679
rect 9424 15630 9494 15645
rect 9790 15715 9858 15732
rect 9790 15681 9807 15715
rect 9841 15681 9858 15715
rect 9790 15566 9858 15681
rect 10528 15679 10598 15880
rect 10528 15645 10547 15679
rect 10581 15645 10598 15679
rect 10528 15630 10598 15645
rect 10894 15715 10962 15732
rect 10894 15681 10911 15715
rect 10945 15681 10962 15715
rect 10894 15566 10962 15681
rect 11632 15679 11702 15880
rect 12417 15862 12429 15896
rect 12463 15862 12475 15896
rect 12417 15803 12475 15862
rect 12417 15769 12429 15803
rect 12463 15769 12475 15803
rect 12417 15734 12475 15769
rect 12601 15925 13119 15967
rect 12601 15891 12619 15925
rect 12653 15891 13067 15925
rect 13101 15891 13119 15925
rect 12601 15823 13119 15891
rect 13154 15925 14223 15967
rect 13154 15891 13171 15925
rect 13205 15891 14171 15925
rect 14205 15891 14223 15925
rect 13154 15880 14223 15891
rect 14258 15925 15327 15967
rect 14258 15891 14275 15925
rect 14309 15891 15275 15925
rect 15309 15891 15327 15925
rect 14258 15880 15327 15891
rect 15362 15925 16431 15967
rect 15362 15891 15379 15925
rect 15413 15891 16379 15925
rect 16413 15891 16431 15925
rect 15362 15880 16431 15891
rect 16466 15925 17535 15967
rect 16466 15891 16483 15925
rect 16517 15891 17483 15925
rect 17517 15891 17535 15925
rect 16466 15880 17535 15891
rect 17569 15896 17627 15967
rect 12601 15789 12619 15823
rect 12653 15789 13067 15823
rect 13101 15789 13119 15823
rect 12601 15749 13119 15789
rect 11632 15645 11651 15679
rect 11685 15645 11702 15679
rect 11632 15630 11702 15645
rect 11998 15715 12066 15732
rect 11998 15681 12015 15715
rect 12049 15681 12066 15715
rect 11998 15566 12066 15681
rect 12601 15679 12843 15749
rect 12601 15645 12679 15679
rect 12713 15645 12789 15679
rect 12823 15645 12843 15679
rect 12877 15681 12897 15715
rect 12931 15681 13007 15715
rect 13041 15681 13119 15715
rect 12877 15611 13119 15681
rect 13472 15679 13542 15880
rect 13472 15645 13491 15679
rect 13525 15645 13542 15679
rect 13472 15630 13542 15645
rect 13838 15715 13906 15732
rect 13838 15681 13855 15715
rect 13889 15681 13906 15715
rect 12417 15585 12475 15602
rect 7449 15518 7467 15552
rect 7501 15518 7915 15552
rect 7949 15518 7967 15552
rect 7449 15457 7967 15518
rect 8002 15552 9071 15566
rect 8002 15518 8019 15552
rect 8053 15518 9019 15552
rect 9053 15518 9071 15552
rect 8002 15457 9071 15518
rect 9106 15552 10175 15566
rect 9106 15518 9123 15552
rect 9157 15518 10123 15552
rect 10157 15518 10175 15552
rect 9106 15457 10175 15518
rect 10210 15552 11279 15566
rect 10210 15518 10227 15552
rect 10261 15518 11227 15552
rect 11261 15518 11279 15552
rect 10210 15457 11279 15518
rect 11314 15552 12383 15566
rect 11314 15518 11331 15552
rect 11365 15518 12331 15552
rect 12365 15518 12383 15552
rect 11314 15457 12383 15518
rect 12417 15551 12429 15585
rect 12463 15551 12475 15585
rect 12417 15457 12475 15551
rect 12601 15552 13119 15611
rect 13838 15566 13906 15681
rect 14576 15679 14646 15880
rect 14576 15645 14595 15679
rect 14629 15645 14646 15679
rect 14576 15630 14646 15645
rect 14942 15715 15010 15732
rect 14942 15681 14959 15715
rect 14993 15681 15010 15715
rect 14942 15566 15010 15681
rect 15680 15679 15750 15880
rect 15680 15645 15699 15679
rect 15733 15645 15750 15679
rect 15680 15630 15750 15645
rect 16046 15715 16114 15732
rect 16046 15681 16063 15715
rect 16097 15681 16114 15715
rect 16046 15566 16114 15681
rect 16784 15679 16854 15880
rect 17569 15862 17581 15896
rect 17615 15862 17627 15896
rect 17754 15925 18823 15967
rect 17754 15891 17771 15925
rect 17805 15891 18771 15925
rect 18805 15891 18823 15925
rect 17754 15880 18823 15891
rect 18858 15925 19927 15967
rect 18858 15891 18875 15925
rect 18909 15891 19875 15925
rect 19909 15891 19927 15925
rect 18858 15880 19927 15891
rect 19961 15925 20203 15967
rect 19961 15891 19979 15925
rect 20013 15891 20151 15925
rect 20185 15891 20203 15925
rect 17569 15803 17627 15862
rect 17569 15769 17581 15803
rect 17615 15769 17627 15803
rect 17569 15734 17627 15769
rect 16784 15645 16803 15679
rect 16837 15645 16854 15679
rect 16784 15630 16854 15645
rect 17150 15715 17218 15732
rect 17150 15681 17167 15715
rect 17201 15681 17218 15715
rect 17150 15566 17218 15681
rect 18072 15679 18142 15880
rect 18072 15645 18091 15679
rect 18125 15645 18142 15679
rect 18072 15630 18142 15645
rect 18438 15715 18506 15732
rect 18438 15681 18455 15715
rect 18489 15681 18506 15715
rect 17569 15585 17627 15602
rect 12601 15518 12619 15552
rect 12653 15518 13067 15552
rect 13101 15518 13119 15552
rect 12601 15457 13119 15518
rect 13154 15552 14223 15566
rect 13154 15518 13171 15552
rect 13205 15518 14171 15552
rect 14205 15518 14223 15552
rect 13154 15457 14223 15518
rect 14258 15552 15327 15566
rect 14258 15518 14275 15552
rect 14309 15518 15275 15552
rect 15309 15518 15327 15552
rect 14258 15457 15327 15518
rect 15362 15552 16431 15566
rect 15362 15518 15379 15552
rect 15413 15518 16379 15552
rect 16413 15518 16431 15552
rect 15362 15457 16431 15518
rect 16466 15552 17535 15566
rect 16466 15518 16483 15552
rect 16517 15518 17483 15552
rect 17517 15518 17535 15552
rect 16466 15457 17535 15518
rect 17569 15551 17581 15585
rect 17615 15551 17627 15585
rect 18438 15566 18506 15681
rect 19176 15679 19246 15880
rect 19961 15830 20203 15891
rect 19961 15796 19979 15830
rect 20013 15796 20151 15830
rect 20185 15796 20203 15830
rect 19961 15749 20203 15796
rect 19176 15645 19195 15679
rect 19229 15645 19246 15679
rect 19176 15630 19246 15645
rect 19542 15715 19610 15732
rect 19542 15681 19559 15715
rect 19593 15681 19610 15715
rect 19542 15566 19610 15681
rect 19961 15675 20065 15749
rect 19961 15641 20011 15675
rect 20045 15641 20065 15675
rect 20099 15681 20119 15715
rect 20153 15681 20203 15715
rect 20099 15607 20203 15681
rect 17569 15457 17627 15551
rect 17754 15552 18823 15566
rect 17754 15518 17771 15552
rect 17805 15518 18771 15552
rect 18805 15518 18823 15552
rect 17754 15457 18823 15518
rect 18858 15552 19927 15566
rect 18858 15518 18875 15552
rect 18909 15518 19875 15552
rect 19909 15518 19927 15552
rect 18858 15457 19927 15518
rect 19961 15554 20203 15607
rect 19961 15520 19979 15554
rect 20013 15520 20151 15554
rect 20185 15520 20203 15554
rect 19961 15457 20203 15520
rect 4948 15423 4977 15457
rect 5011 15423 5069 15457
rect 5103 15423 5161 15457
rect 5195 15423 5253 15457
rect 5287 15423 5345 15457
rect 5379 15423 5437 15457
rect 5471 15423 5529 15457
rect 5563 15423 5621 15457
rect 5655 15423 5713 15457
rect 5747 15423 5805 15457
rect 5839 15423 5897 15457
rect 5931 15423 5989 15457
rect 6023 15423 6081 15457
rect 6115 15423 6173 15457
rect 6207 15423 6265 15457
rect 6299 15423 6357 15457
rect 6391 15423 6449 15457
rect 6483 15423 6541 15457
rect 6575 15423 6633 15457
rect 6667 15423 6725 15457
rect 6759 15423 6817 15457
rect 6851 15423 6909 15457
rect 6943 15423 7001 15457
rect 7035 15423 7093 15457
rect 7127 15423 7185 15457
rect 7219 15423 7277 15457
rect 7311 15423 7369 15457
rect 7403 15423 7461 15457
rect 7495 15423 7553 15457
rect 7587 15423 7645 15457
rect 7679 15423 7737 15457
rect 7771 15423 7829 15457
rect 7863 15423 7921 15457
rect 7955 15423 8013 15457
rect 8047 15423 8105 15457
rect 8139 15423 8197 15457
rect 8231 15423 8289 15457
rect 8323 15423 8381 15457
rect 8415 15423 8473 15457
rect 8507 15423 8565 15457
rect 8599 15423 8657 15457
rect 8691 15423 8749 15457
rect 8783 15423 8841 15457
rect 8875 15423 8933 15457
rect 8967 15423 9025 15457
rect 9059 15423 9117 15457
rect 9151 15423 9209 15457
rect 9243 15423 9301 15457
rect 9335 15423 9393 15457
rect 9427 15423 9485 15457
rect 9519 15423 9577 15457
rect 9611 15423 9669 15457
rect 9703 15423 9761 15457
rect 9795 15423 9853 15457
rect 9887 15423 9945 15457
rect 9979 15423 10037 15457
rect 10071 15423 10129 15457
rect 10163 15423 10221 15457
rect 10255 15423 10313 15457
rect 10347 15423 10405 15457
rect 10439 15423 10497 15457
rect 10531 15423 10589 15457
rect 10623 15423 10681 15457
rect 10715 15423 10773 15457
rect 10807 15423 10865 15457
rect 10899 15423 10957 15457
rect 10991 15423 11049 15457
rect 11083 15423 11141 15457
rect 11175 15423 11233 15457
rect 11267 15423 11325 15457
rect 11359 15423 11417 15457
rect 11451 15423 11509 15457
rect 11543 15423 11601 15457
rect 11635 15423 11693 15457
rect 11727 15423 11785 15457
rect 11819 15423 11877 15457
rect 11911 15423 11969 15457
rect 12003 15423 12061 15457
rect 12095 15423 12153 15457
rect 12187 15423 12245 15457
rect 12279 15423 12337 15457
rect 12371 15423 12429 15457
rect 12463 15423 12521 15457
rect 12555 15423 12613 15457
rect 12647 15423 12705 15457
rect 12739 15423 12797 15457
rect 12831 15423 12889 15457
rect 12923 15423 12981 15457
rect 13015 15423 13073 15457
rect 13107 15423 13165 15457
rect 13199 15423 13257 15457
rect 13291 15423 13349 15457
rect 13383 15423 13441 15457
rect 13475 15423 13533 15457
rect 13567 15423 13625 15457
rect 13659 15423 13717 15457
rect 13751 15423 13809 15457
rect 13843 15423 13901 15457
rect 13935 15423 13993 15457
rect 14027 15423 14085 15457
rect 14119 15423 14177 15457
rect 14211 15423 14269 15457
rect 14303 15423 14361 15457
rect 14395 15423 14453 15457
rect 14487 15423 14545 15457
rect 14579 15423 14637 15457
rect 14671 15423 14729 15457
rect 14763 15423 14821 15457
rect 14855 15423 14913 15457
rect 14947 15423 15005 15457
rect 15039 15423 15097 15457
rect 15131 15423 15189 15457
rect 15223 15423 15281 15457
rect 15315 15423 15373 15457
rect 15407 15423 15465 15457
rect 15499 15423 15557 15457
rect 15591 15423 15649 15457
rect 15683 15423 15741 15457
rect 15775 15423 15833 15457
rect 15867 15423 15925 15457
rect 15959 15423 16017 15457
rect 16051 15423 16109 15457
rect 16143 15423 16201 15457
rect 16235 15423 16293 15457
rect 16327 15423 16385 15457
rect 16419 15423 16477 15457
rect 16511 15423 16569 15457
rect 16603 15423 16661 15457
rect 16695 15423 16753 15457
rect 16787 15423 16845 15457
rect 16879 15423 16937 15457
rect 16971 15423 17029 15457
rect 17063 15423 17121 15457
rect 17155 15423 17213 15457
rect 17247 15423 17305 15457
rect 17339 15423 17397 15457
rect 17431 15423 17489 15457
rect 17523 15423 17581 15457
rect 17615 15423 17673 15457
rect 17707 15423 17765 15457
rect 17799 15423 17857 15457
rect 17891 15423 17949 15457
rect 17983 15423 18041 15457
rect 18075 15423 18133 15457
rect 18167 15423 18225 15457
rect 18259 15423 18317 15457
rect 18351 15423 18409 15457
rect 18443 15423 18501 15457
rect 18535 15423 18593 15457
rect 18627 15423 18685 15457
rect 18719 15423 18777 15457
rect 18811 15423 18869 15457
rect 18903 15423 18961 15457
rect 18995 15423 19053 15457
rect 19087 15423 19145 15457
rect 19179 15423 19237 15457
rect 19271 15423 19329 15457
rect 19363 15423 19421 15457
rect 19455 15423 19513 15457
rect 19547 15423 19605 15457
rect 19639 15423 19697 15457
rect 19731 15423 19789 15457
rect 19823 15423 19881 15457
rect 19915 15423 19973 15457
rect 20007 15423 20065 15457
rect 20099 15423 20157 15457
rect 20191 15423 20220 15457
rect 4965 15360 5207 15423
rect 4965 15326 4983 15360
rect 5017 15326 5155 15360
rect 5189 15326 5207 15360
rect 4965 15273 5207 15326
rect 5426 15362 6495 15423
rect 5426 15328 5443 15362
rect 5477 15328 6443 15362
rect 6477 15328 6495 15362
rect 5426 15314 6495 15328
rect 6530 15362 7599 15423
rect 6530 15328 6547 15362
rect 6581 15328 7547 15362
rect 7581 15328 7599 15362
rect 6530 15314 7599 15328
rect 7634 15362 8703 15423
rect 7634 15328 7651 15362
rect 7685 15328 8651 15362
rect 8685 15328 8703 15362
rect 7634 15314 8703 15328
rect 8738 15362 9807 15423
rect 8738 15328 8755 15362
rect 8789 15328 9755 15362
rect 9789 15328 9807 15362
rect 8738 15314 9807 15328
rect 9841 15329 9899 15423
rect 4965 15199 5069 15273
rect 4965 15165 5015 15199
rect 5049 15165 5069 15199
rect 5103 15205 5123 15239
rect 5157 15205 5207 15239
rect 5103 15131 5207 15205
rect 4965 15084 5207 15131
rect 4965 15050 4983 15084
rect 5017 15050 5155 15084
rect 5189 15050 5207 15084
rect 4965 14989 5207 15050
rect 5744 15235 5814 15250
rect 5744 15201 5763 15235
rect 5797 15201 5814 15235
rect 5744 15000 5814 15201
rect 6110 15199 6178 15314
rect 6110 15165 6127 15199
rect 6161 15165 6178 15199
rect 6110 15148 6178 15165
rect 6848 15235 6918 15250
rect 6848 15201 6867 15235
rect 6901 15201 6918 15235
rect 6848 15000 6918 15201
rect 7214 15199 7282 15314
rect 7214 15165 7231 15199
rect 7265 15165 7282 15199
rect 7214 15148 7282 15165
rect 7952 15235 8022 15250
rect 7952 15201 7971 15235
rect 8005 15201 8022 15235
rect 7952 15000 8022 15201
rect 8318 15199 8386 15314
rect 8318 15165 8335 15199
rect 8369 15165 8386 15199
rect 8318 15148 8386 15165
rect 9056 15235 9126 15250
rect 9056 15201 9075 15235
rect 9109 15201 9126 15235
rect 9056 15000 9126 15201
rect 9422 15199 9490 15314
rect 9841 15295 9853 15329
rect 9887 15295 9899 15329
rect 9841 15278 9899 15295
rect 10025 15362 10543 15423
rect 10025 15328 10043 15362
rect 10077 15328 10491 15362
rect 10525 15328 10543 15362
rect 10025 15269 10543 15328
rect 10578 15362 11647 15423
rect 10578 15328 10595 15362
rect 10629 15328 11595 15362
rect 11629 15328 11647 15362
rect 10578 15314 11647 15328
rect 11682 15362 12751 15423
rect 11682 15328 11699 15362
rect 11733 15328 12699 15362
rect 12733 15328 12751 15362
rect 11682 15314 12751 15328
rect 12808 15355 12865 15389
rect 12808 15321 12825 15355
rect 12859 15321 12865 15355
rect 12899 15381 12953 15423
rect 12899 15347 12909 15381
rect 12943 15347 12953 15381
rect 12899 15331 12953 15347
rect 13033 15355 13113 15389
rect 9422 15165 9439 15199
rect 9473 15165 9490 15199
rect 9422 15148 9490 15165
rect 10025 15201 10103 15235
rect 10137 15201 10213 15235
rect 10247 15201 10267 15235
rect 9841 15111 9899 15146
rect 9841 15077 9853 15111
rect 9887 15077 9899 15111
rect 9841 15018 9899 15077
rect 4965 14955 4983 14989
rect 5017 14955 5155 14989
rect 5189 14955 5207 14989
rect 4965 14913 5207 14955
rect 5426 14989 6495 15000
rect 5426 14955 5443 14989
rect 5477 14955 6443 14989
rect 6477 14955 6495 14989
rect 5426 14913 6495 14955
rect 6530 14989 7599 15000
rect 6530 14955 6547 14989
rect 6581 14955 7547 14989
rect 7581 14955 7599 14989
rect 6530 14913 7599 14955
rect 7634 14989 8703 15000
rect 7634 14955 7651 14989
rect 7685 14955 8651 14989
rect 8685 14955 8703 14989
rect 7634 14913 8703 14955
rect 8738 14989 9807 15000
rect 8738 14955 8755 14989
rect 8789 14955 9755 14989
rect 9789 14955 9807 14989
rect 8738 14913 9807 14955
rect 9841 14984 9853 15018
rect 9887 14984 9899 15018
rect 9841 14913 9899 14984
rect 10025 15131 10267 15201
rect 10301 15199 10543 15269
rect 10301 15165 10321 15199
rect 10355 15165 10431 15199
rect 10465 15165 10543 15199
rect 10896 15235 10966 15250
rect 10896 15201 10915 15235
rect 10949 15201 10966 15235
rect 10025 15091 10543 15131
rect 10025 15057 10043 15091
rect 10077 15057 10491 15091
rect 10525 15057 10543 15091
rect 10025 14989 10543 15057
rect 10896 15000 10966 15201
rect 11262 15199 11330 15314
rect 11262 15165 11279 15199
rect 11313 15165 11330 15199
rect 11262 15148 11330 15165
rect 12000 15235 12070 15250
rect 12000 15201 12019 15235
rect 12053 15201 12070 15235
rect 12000 15000 12070 15201
rect 12366 15199 12434 15314
rect 12808 15297 12865 15321
rect 13033 15321 13063 15355
rect 13097 15321 13113 15355
rect 12808 15263 12999 15297
rect 12366 15165 12383 15199
rect 12417 15165 12434 15199
rect 12366 15148 12434 15165
rect 12785 15225 12923 15229
rect 12785 15191 12849 15225
rect 12883 15191 12923 15225
rect 12785 15151 12923 15191
rect 12785 15117 12889 15151
rect 12957 15225 12999 15263
rect 12957 15191 12963 15225
rect 12997 15191 12999 15225
rect 12957 15083 12999 15191
rect 12808 15039 12999 15083
rect 13033 15229 13113 15321
rect 13151 15355 13207 15389
rect 13151 15321 13167 15355
rect 13201 15321 13207 15355
rect 13311 15381 13376 15423
rect 13311 15347 13326 15381
rect 13360 15347 13376 15381
rect 13311 15331 13376 15347
rect 13410 15355 13487 15389
rect 13151 15297 13207 15321
rect 13410 15321 13416 15355
rect 13450 15321 13487 15355
rect 13151 15263 13376 15297
rect 13410 15275 13487 15321
rect 13286 15241 13376 15263
rect 13033 15225 13252 15229
rect 13033 15191 13167 15225
rect 13201 15191 13252 15225
rect 13033 15117 13252 15191
rect 13286 15225 13397 15241
rect 13286 15191 13363 15225
rect 13286 15175 13397 15191
rect 12808 15015 12865 15039
rect 10025 14955 10043 14989
rect 10077 14955 10491 14989
rect 10525 14955 10543 14989
rect 10025 14913 10543 14955
rect 10578 14989 11647 15000
rect 10578 14955 10595 14989
rect 10629 14955 11595 14989
rect 11629 14955 11647 14989
rect 10578 14913 11647 14955
rect 11682 14989 12751 15000
rect 11682 14955 11699 14989
rect 11733 14955 12699 14989
rect 12733 14955 12751 14989
rect 11682 14913 12751 14955
rect 12808 14981 12825 15015
rect 12859 14981 12865 15015
rect 13033 15015 13113 15117
rect 13286 15083 13376 15175
rect 13431 15141 13487 15275
rect 13521 15355 13855 15423
rect 13521 15321 13539 15355
rect 13573 15321 13803 15355
rect 13837 15321 13855 15355
rect 13521 15269 13855 15321
rect 13890 15362 14959 15423
rect 13890 15328 13907 15362
rect 13941 15328 14907 15362
rect 14941 15328 14959 15362
rect 13890 15314 14959 15328
rect 14993 15329 15051 15423
rect 12808 14947 12865 14981
rect 12899 14989 12953 15005
rect 12899 14955 12909 14989
rect 12943 14955 12953 14989
rect 12899 14913 12953 14955
rect 13033 14981 13063 15015
rect 13097 14981 13113 15015
rect 13033 14947 13113 14981
rect 13151 15039 13376 15083
rect 13151 15015 13207 15039
rect 13151 14981 13167 15015
rect 13201 14981 13207 15015
rect 13410 15015 13487 15141
rect 13151 14947 13207 14981
rect 13311 14989 13376 15005
rect 13311 14955 13326 14989
rect 13360 14955 13376 14989
rect 13311 14913 13376 14955
rect 13410 14981 13416 15015
rect 13475 14981 13487 15015
rect 13410 14947 13487 14981
rect 13521 15201 13541 15235
rect 13575 15201 13671 15235
rect 13521 15131 13671 15201
rect 13705 15199 13855 15269
rect 13705 15165 13801 15199
rect 13835 15165 13855 15199
rect 14208 15235 14278 15250
rect 14208 15201 14227 15235
rect 14261 15201 14278 15235
rect 13521 15091 13855 15131
rect 13521 15057 13539 15091
rect 13573 15057 13803 15091
rect 13837 15057 13855 15091
rect 13521 14989 13855 15057
rect 14208 15000 14278 15201
rect 14574 15199 14642 15314
rect 14993 15295 15005 15329
rect 15039 15295 15051 15329
rect 14993 15278 15051 15295
rect 15085 15360 15327 15423
rect 15085 15326 15103 15360
rect 15137 15326 15275 15360
rect 15309 15326 15327 15360
rect 15085 15273 15327 15326
rect 14574 15165 14591 15199
rect 14625 15165 14642 15199
rect 14574 15148 14642 15165
rect 15085 15205 15135 15239
rect 15169 15205 15189 15239
rect 14993 15111 15051 15146
rect 14993 15077 15005 15111
rect 15039 15077 15051 15111
rect 14993 15018 15051 15077
rect 13521 14955 13539 14989
rect 13573 14955 13803 14989
rect 13837 14955 13855 14989
rect 13521 14913 13855 14955
rect 13890 14989 14959 15000
rect 13890 14955 13907 14989
rect 13941 14955 14907 14989
rect 14941 14955 14959 14989
rect 13890 14913 14959 14955
rect 14993 14984 15005 15018
rect 15039 14984 15051 15018
rect 14993 14913 15051 14984
rect 15085 15131 15189 15205
rect 15223 15199 15327 15273
rect 15384 15355 15441 15389
rect 15384 15321 15401 15355
rect 15435 15321 15441 15355
rect 15475 15381 15529 15423
rect 15475 15347 15485 15381
rect 15519 15347 15529 15381
rect 15475 15331 15529 15347
rect 15609 15355 15689 15389
rect 15384 15297 15441 15321
rect 15609 15321 15639 15355
rect 15673 15321 15689 15355
rect 15384 15263 15575 15297
rect 15223 15165 15243 15199
rect 15277 15165 15327 15199
rect 15361 15225 15499 15229
rect 15361 15191 15425 15225
rect 15459 15191 15499 15225
rect 15361 15151 15499 15191
rect 15085 15084 15327 15131
rect 15361 15117 15373 15151
rect 15407 15117 15499 15151
rect 15533 15225 15575 15263
rect 15533 15191 15539 15225
rect 15573 15191 15575 15225
rect 15085 15050 15103 15084
rect 15137 15050 15275 15084
rect 15309 15050 15327 15084
rect 15533 15083 15575 15191
rect 15085 14989 15327 15050
rect 15085 14955 15103 14989
rect 15137 14955 15275 14989
rect 15309 14955 15327 14989
rect 15085 14913 15327 14955
rect 15384 15039 15575 15083
rect 15609 15229 15689 15321
rect 15727 15355 15783 15389
rect 15727 15321 15743 15355
rect 15777 15321 15783 15355
rect 15887 15381 15952 15423
rect 15887 15347 15902 15381
rect 15936 15347 15952 15381
rect 15887 15331 15952 15347
rect 15986 15355 16063 15389
rect 15727 15297 15783 15321
rect 15986 15321 15992 15355
rect 16026 15321 16063 15355
rect 15727 15263 15952 15297
rect 15986 15275 16063 15321
rect 15862 15241 15952 15263
rect 15609 15225 15828 15229
rect 15609 15191 15743 15225
rect 15777 15191 15828 15225
rect 15609 15117 15828 15191
rect 15862 15225 15973 15241
rect 15862 15191 15939 15225
rect 15862 15175 15973 15191
rect 15384 15015 15441 15039
rect 15384 14981 15401 15015
rect 15435 14981 15441 15015
rect 15609 15015 15689 15117
rect 15862 15083 15952 15175
rect 16007 15141 16063 15275
rect 16097 15362 16615 15423
rect 16097 15328 16115 15362
rect 16149 15328 16563 15362
rect 16597 15328 16615 15362
rect 16097 15269 16615 15328
rect 16650 15362 17719 15423
rect 16650 15328 16667 15362
rect 16701 15328 17667 15362
rect 17701 15328 17719 15362
rect 16650 15314 17719 15328
rect 17754 15362 18823 15423
rect 17754 15328 17771 15362
rect 17805 15328 18771 15362
rect 18805 15328 18823 15362
rect 17754 15314 18823 15328
rect 18858 15362 19927 15423
rect 18858 15328 18875 15362
rect 18909 15328 19875 15362
rect 19909 15328 19927 15362
rect 18858 15314 19927 15328
rect 19961 15360 20203 15423
rect 19961 15326 19979 15360
rect 20013 15326 20151 15360
rect 20185 15326 20203 15360
rect 15384 14947 15441 14981
rect 15475 14989 15529 15005
rect 15475 14955 15485 14989
rect 15519 14955 15529 14989
rect 15475 14913 15529 14955
rect 15609 14981 15639 15015
rect 15673 14981 15689 15015
rect 15609 14947 15689 14981
rect 15727 15039 15952 15083
rect 15727 15015 15783 15039
rect 15727 14981 15743 15015
rect 15777 14981 15783 15015
rect 15986 15015 16063 15141
rect 15727 14947 15783 14981
rect 15887 14989 15952 15005
rect 15887 14955 15902 14989
rect 15936 14955 15952 14989
rect 15887 14913 15952 14955
rect 15986 14981 15992 15015
rect 16051 14981 16063 15015
rect 15986 14947 16063 14981
rect 16097 15201 16175 15235
rect 16209 15201 16285 15235
rect 16319 15201 16339 15235
rect 16097 15131 16339 15201
rect 16373 15199 16615 15269
rect 16373 15165 16393 15199
rect 16427 15165 16503 15199
rect 16537 15165 16615 15199
rect 16968 15235 17038 15250
rect 16968 15201 16987 15235
rect 17021 15201 17038 15235
rect 16097 15091 16615 15131
rect 16097 15057 16115 15091
rect 16149 15057 16563 15091
rect 16597 15057 16615 15091
rect 16097 14989 16615 15057
rect 16968 15000 17038 15201
rect 17334 15199 17402 15314
rect 17334 15165 17351 15199
rect 17385 15165 17402 15199
rect 17334 15148 17402 15165
rect 18072 15235 18142 15250
rect 18072 15201 18091 15235
rect 18125 15201 18142 15235
rect 18072 15000 18142 15201
rect 18438 15199 18506 15314
rect 18438 15165 18455 15199
rect 18489 15165 18506 15199
rect 18438 15148 18506 15165
rect 19176 15235 19246 15250
rect 19176 15201 19195 15235
rect 19229 15201 19246 15235
rect 19176 15000 19246 15201
rect 19542 15199 19610 15314
rect 19961 15273 20203 15326
rect 19542 15165 19559 15199
rect 19593 15165 19610 15199
rect 19542 15148 19610 15165
rect 19961 15205 20011 15239
rect 20045 15205 20065 15239
rect 19961 15131 20065 15205
rect 20099 15199 20203 15273
rect 20099 15165 20119 15199
rect 20153 15165 20203 15199
rect 19961 15084 20203 15131
rect 19961 15050 19979 15084
rect 20013 15050 20151 15084
rect 20185 15050 20203 15084
rect 16097 14955 16115 14989
rect 16149 14955 16563 14989
rect 16597 14955 16615 14989
rect 16097 14913 16615 14955
rect 16650 14989 17719 15000
rect 16650 14955 16667 14989
rect 16701 14955 17667 14989
rect 17701 14955 17719 14989
rect 16650 14913 17719 14955
rect 17754 14989 18823 15000
rect 17754 14955 17771 14989
rect 17805 14955 18771 14989
rect 18805 14955 18823 14989
rect 17754 14913 18823 14955
rect 18858 14989 19927 15000
rect 18858 14955 18875 14989
rect 18909 14955 19875 14989
rect 19909 14955 19927 14989
rect 18858 14913 19927 14955
rect 19961 14989 20203 15050
rect 19961 14955 19979 14989
rect 20013 14955 20151 14989
rect 20185 14955 20203 14989
rect 19961 14913 20203 14955
rect 4948 14879 4977 14913
rect 5011 14879 5069 14913
rect 5103 14879 5161 14913
rect 5195 14879 5253 14913
rect 5287 14879 5345 14913
rect 5379 14879 5437 14913
rect 5471 14879 5529 14913
rect 5563 14879 5621 14913
rect 5655 14879 5713 14913
rect 5747 14879 5805 14913
rect 5839 14879 5897 14913
rect 5931 14879 5989 14913
rect 6023 14879 6081 14913
rect 6115 14879 6173 14913
rect 6207 14879 6265 14913
rect 6299 14879 6357 14913
rect 6391 14879 6449 14913
rect 6483 14879 6541 14913
rect 6575 14879 6633 14913
rect 6667 14879 6725 14913
rect 6759 14879 6817 14913
rect 6851 14879 6909 14913
rect 6943 14879 7001 14913
rect 7035 14879 7093 14913
rect 7127 14879 7185 14913
rect 7219 14879 7277 14913
rect 7311 14879 7369 14913
rect 7403 14879 7461 14913
rect 7495 14879 7553 14913
rect 7587 14879 7645 14913
rect 7679 14879 7737 14913
rect 7771 14879 7829 14913
rect 7863 14879 7921 14913
rect 7955 14879 8013 14913
rect 8047 14879 8105 14913
rect 8139 14879 8197 14913
rect 8231 14879 8289 14913
rect 8323 14879 8381 14913
rect 8415 14879 8473 14913
rect 8507 14879 8565 14913
rect 8599 14879 8657 14913
rect 8691 14879 8749 14913
rect 8783 14879 8841 14913
rect 8875 14879 8933 14913
rect 8967 14879 9025 14913
rect 9059 14879 9117 14913
rect 9151 14879 9209 14913
rect 9243 14879 9301 14913
rect 9335 14879 9393 14913
rect 9427 14879 9485 14913
rect 9519 14879 9577 14913
rect 9611 14879 9669 14913
rect 9703 14879 9761 14913
rect 9795 14879 9853 14913
rect 9887 14879 9945 14913
rect 9979 14879 10037 14913
rect 10071 14879 10129 14913
rect 10163 14879 10221 14913
rect 10255 14879 10313 14913
rect 10347 14879 10405 14913
rect 10439 14879 10497 14913
rect 10531 14879 10589 14913
rect 10623 14879 10681 14913
rect 10715 14879 10773 14913
rect 10807 14879 10865 14913
rect 10899 14879 10957 14913
rect 10991 14879 11049 14913
rect 11083 14879 11141 14913
rect 11175 14879 11233 14913
rect 11267 14879 11325 14913
rect 11359 14879 11417 14913
rect 11451 14879 11509 14913
rect 11543 14879 11601 14913
rect 11635 14879 11693 14913
rect 11727 14879 11785 14913
rect 11819 14879 11877 14913
rect 11911 14879 11969 14913
rect 12003 14879 12061 14913
rect 12095 14879 12153 14913
rect 12187 14879 12245 14913
rect 12279 14879 12337 14913
rect 12371 14879 12429 14913
rect 12463 14879 12521 14913
rect 12555 14879 12613 14913
rect 12647 14879 12705 14913
rect 12739 14879 12797 14913
rect 12831 14879 12889 14913
rect 12923 14879 12981 14913
rect 13015 14879 13073 14913
rect 13107 14879 13165 14913
rect 13199 14879 13257 14913
rect 13291 14879 13349 14913
rect 13383 14879 13441 14913
rect 13475 14879 13533 14913
rect 13567 14879 13625 14913
rect 13659 14879 13717 14913
rect 13751 14879 13809 14913
rect 13843 14879 13901 14913
rect 13935 14879 13993 14913
rect 14027 14879 14085 14913
rect 14119 14879 14177 14913
rect 14211 14879 14269 14913
rect 14303 14879 14361 14913
rect 14395 14879 14453 14913
rect 14487 14879 14545 14913
rect 14579 14879 14637 14913
rect 14671 14879 14729 14913
rect 14763 14879 14821 14913
rect 14855 14879 14913 14913
rect 14947 14879 15005 14913
rect 15039 14879 15097 14913
rect 15131 14879 15189 14913
rect 15223 14879 15281 14913
rect 15315 14879 15373 14913
rect 15407 14879 15465 14913
rect 15499 14879 15557 14913
rect 15591 14879 15649 14913
rect 15683 14879 15741 14913
rect 15775 14879 15833 14913
rect 15867 14879 15925 14913
rect 15959 14879 16017 14913
rect 16051 14879 16109 14913
rect 16143 14879 16201 14913
rect 16235 14879 16293 14913
rect 16327 14879 16385 14913
rect 16419 14879 16477 14913
rect 16511 14879 16569 14913
rect 16603 14879 16661 14913
rect 16695 14879 16753 14913
rect 16787 14879 16845 14913
rect 16879 14879 16937 14913
rect 16971 14879 17029 14913
rect 17063 14879 17121 14913
rect 17155 14879 17213 14913
rect 17247 14879 17305 14913
rect 17339 14879 17397 14913
rect 17431 14879 17489 14913
rect 17523 14879 17581 14913
rect 17615 14879 17673 14913
rect 17707 14879 17765 14913
rect 17799 14879 17857 14913
rect 17891 14879 17949 14913
rect 17983 14879 18041 14913
rect 18075 14879 18133 14913
rect 18167 14879 18225 14913
rect 18259 14879 18317 14913
rect 18351 14879 18409 14913
rect 18443 14879 18501 14913
rect 18535 14879 18593 14913
rect 18627 14879 18685 14913
rect 18719 14879 18777 14913
rect 18811 14879 18869 14913
rect 18903 14879 18961 14913
rect 18995 14879 19053 14913
rect 19087 14879 19145 14913
rect 19179 14879 19237 14913
rect 19271 14879 19329 14913
rect 19363 14879 19421 14913
rect 19455 14879 19513 14913
rect 19547 14879 19605 14913
rect 19639 14879 19697 14913
rect 19731 14879 19789 14913
rect 19823 14879 19881 14913
rect 19915 14879 19973 14913
rect 20007 14879 20065 14913
rect 20099 14879 20157 14913
rect 20191 14879 20220 14913
rect 4965 14837 5207 14879
rect 4965 14803 4983 14837
rect 5017 14803 5155 14837
rect 5189 14803 5207 14837
rect 4965 14742 5207 14803
rect 4965 14708 4983 14742
rect 5017 14708 5155 14742
rect 5189 14708 5207 14742
rect 4965 14661 5207 14708
rect 4965 14593 5015 14627
rect 5049 14593 5069 14627
rect 4965 14519 5069 14593
rect 5103 14587 5207 14661
rect 5103 14553 5123 14587
rect 5157 14553 5207 14587
rect 5425 14837 6127 14879
rect 5425 14803 5443 14837
rect 5477 14803 6075 14837
rect 6109 14803 6127 14837
rect 5425 14735 6127 14803
rect 6162 14837 7231 14879
rect 6162 14803 6179 14837
rect 6213 14803 7179 14837
rect 7213 14803 7231 14837
rect 6162 14792 7231 14803
rect 7265 14808 7323 14879
rect 5425 14701 5443 14735
rect 5477 14701 6075 14735
rect 6109 14701 6127 14735
rect 5425 14661 6127 14701
rect 5425 14591 5763 14661
rect 5425 14557 5503 14591
rect 5537 14557 5606 14591
rect 5640 14557 5709 14591
rect 5743 14557 5763 14591
rect 5797 14593 5817 14627
rect 5851 14593 5916 14627
rect 5950 14593 6015 14627
rect 6049 14593 6127 14627
rect 5797 14523 6127 14593
rect 6480 14591 6550 14792
rect 7265 14774 7277 14808
rect 7311 14774 7323 14808
rect 7358 14837 8427 14879
rect 7358 14803 7375 14837
rect 7409 14803 8375 14837
rect 8409 14803 8427 14837
rect 7358 14792 8427 14803
rect 8462 14837 9531 14879
rect 8462 14803 8479 14837
rect 8513 14803 9479 14837
rect 9513 14803 9531 14837
rect 8462 14792 9531 14803
rect 9566 14837 10635 14879
rect 9566 14803 9583 14837
rect 9617 14803 10583 14837
rect 10617 14803 10635 14837
rect 9566 14792 10635 14803
rect 7265 14715 7323 14774
rect 7265 14681 7277 14715
rect 7311 14681 7323 14715
rect 7265 14646 7323 14681
rect 6480 14557 6499 14591
rect 6533 14557 6550 14591
rect 6480 14542 6550 14557
rect 6846 14627 6914 14644
rect 6846 14593 6863 14627
rect 6897 14593 6914 14627
rect 4965 14466 5207 14519
rect 4965 14432 4983 14466
rect 5017 14432 5155 14466
rect 5189 14432 5207 14466
rect 4965 14369 5207 14432
rect 5425 14464 6127 14523
rect 6846 14478 6914 14593
rect 7676 14591 7746 14792
rect 7676 14557 7695 14591
rect 7729 14557 7746 14591
rect 7676 14542 7746 14557
rect 8042 14627 8110 14644
rect 8042 14593 8059 14627
rect 8093 14593 8110 14627
rect 7265 14497 7323 14514
rect 5425 14430 5443 14464
rect 5477 14430 6075 14464
rect 6109 14430 6127 14464
rect 5425 14369 6127 14430
rect 6162 14464 7231 14478
rect 6162 14430 6179 14464
rect 6213 14430 7179 14464
rect 7213 14430 7231 14464
rect 6162 14369 7231 14430
rect 7265 14463 7277 14497
rect 7311 14463 7323 14497
rect 8042 14478 8110 14593
rect 8780 14591 8850 14792
rect 8780 14557 8799 14591
rect 8833 14557 8850 14591
rect 8780 14542 8850 14557
rect 9146 14627 9214 14644
rect 9146 14593 9163 14627
rect 9197 14593 9214 14627
rect 9146 14478 9214 14593
rect 9884 14591 9954 14792
rect 10669 14777 10772 14809
rect 10669 14743 10733 14777
rect 10767 14743 10772 14777
rect 10669 14727 10772 14743
rect 10819 14777 10853 14879
rect 10819 14727 10853 14743
rect 10887 14811 11293 14845
rect 9884 14557 9903 14591
rect 9937 14557 9954 14591
rect 9884 14542 9954 14557
rect 10250 14627 10318 14644
rect 10250 14593 10267 14627
rect 10301 14593 10318 14627
rect 10250 14478 10318 14593
rect 10669 14565 10737 14727
rect 10887 14678 10921 14811
rect 11000 14743 11016 14777
rect 11050 14743 11091 14777
rect 11125 14743 11225 14777
rect 10771 14644 10787 14678
rect 10821 14675 10921 14678
rect 10821 14644 10865 14675
rect 10771 14641 10865 14644
rect 10899 14641 10921 14675
rect 10771 14640 10921 14641
rect 10955 14678 11157 14709
rect 10989 14675 11157 14678
rect 10989 14644 10993 14675
rect 10669 14531 10865 14565
rect 10899 14531 10915 14565
rect 7265 14369 7323 14463
rect 7358 14464 8427 14478
rect 7358 14430 7375 14464
rect 7409 14430 8375 14464
rect 8409 14430 8427 14464
rect 7358 14369 8427 14430
rect 8462 14464 9531 14478
rect 8462 14430 8479 14464
rect 8513 14430 9479 14464
rect 9513 14430 9531 14464
rect 8462 14369 9531 14430
rect 9566 14464 10635 14478
rect 9566 14430 9583 14464
rect 9617 14430 10583 14464
rect 10617 14430 10635 14464
rect 9566 14369 10635 14430
rect 10724 14460 10773 14531
rect 10724 14426 10733 14460
rect 10767 14426 10773 14460
rect 10724 14410 10773 14426
rect 10817 14460 10919 14476
rect 10851 14426 10885 14460
rect 10817 14369 10919 14426
rect 10955 14471 10993 14644
rect 10955 14437 10957 14471
rect 10991 14437 10993 14471
rect 10955 14403 10993 14437
rect 11027 14607 11082 14635
rect 11027 14573 11049 14607
rect 11027 14565 11082 14573
rect 11061 14531 11082 14565
rect 11027 14403 11082 14531
rect 11123 14565 11157 14675
rect 11123 14515 11157 14531
rect 11191 14517 11225 14743
rect 11259 14617 11293 14811
rect 11327 14837 11361 14879
rect 11327 14769 11361 14803
rect 11327 14701 11361 14735
rect 11327 14651 11361 14667
rect 11395 14837 11462 14845
rect 11395 14803 11411 14837
rect 11445 14803 11462 14837
rect 11395 14769 11462 14803
rect 11395 14735 11411 14769
rect 11445 14735 11462 14769
rect 11395 14701 11462 14735
rect 11395 14667 11411 14701
rect 11445 14667 11462 14701
rect 11395 14651 11462 14667
rect 11259 14601 11298 14617
rect 11259 14567 11264 14601
rect 11259 14551 11298 14567
rect 11343 14601 11394 14617
rect 11343 14567 11360 14601
rect 11343 14551 11394 14567
rect 11343 14517 11377 14551
rect 11428 14517 11462 14651
rect 11681 14837 12383 14879
rect 11681 14803 11699 14837
rect 11733 14803 12331 14837
rect 12365 14803 12383 14837
rect 11681 14735 12383 14803
rect 11681 14701 11699 14735
rect 11733 14701 12331 14735
rect 12365 14701 12383 14735
rect 11681 14661 12383 14701
rect 12417 14808 12475 14879
rect 12417 14774 12429 14808
rect 12463 14774 12475 14808
rect 12417 14715 12475 14774
rect 12417 14681 12429 14715
rect 12463 14681 12475 14715
rect 11681 14591 12019 14661
rect 12417 14646 12475 14681
rect 12693 14777 12796 14809
rect 12693 14743 12757 14777
rect 12791 14743 12796 14777
rect 12693 14727 12796 14743
rect 12843 14777 12877 14879
rect 12843 14727 12877 14743
rect 12911 14811 13317 14845
rect 11681 14557 11759 14591
rect 11793 14557 11862 14591
rect 11896 14557 11965 14591
rect 11999 14557 12019 14591
rect 12053 14593 12073 14627
rect 12107 14593 12172 14627
rect 12206 14593 12271 14627
rect 12305 14593 12383 14627
rect 12053 14523 12383 14593
rect 12693 14565 12761 14727
rect 12911 14678 12945 14811
rect 13024 14743 13040 14777
rect 13074 14743 13115 14777
rect 13149 14743 13249 14777
rect 12795 14644 12811 14678
rect 12845 14675 12945 14678
rect 12845 14644 12889 14675
rect 12795 14641 12889 14644
rect 12923 14641 12945 14675
rect 12795 14640 12945 14641
rect 12979 14678 13181 14709
rect 13013 14675 13181 14678
rect 13013 14644 13017 14675
rect 12693 14531 12889 14565
rect 12923 14531 12939 14565
rect 11191 14483 11377 14517
rect 11191 14476 11226 14483
rect 11120 14460 11226 14476
rect 11154 14426 11226 14460
rect 11411 14471 11462 14517
rect 11411 14464 11417 14471
rect 11120 14403 11226 14426
rect 11311 14445 11377 14449
rect 11311 14411 11327 14445
rect 11361 14411 11377 14445
rect 11311 14369 11377 14411
rect 11451 14437 11462 14471
rect 11445 14430 11462 14437
rect 11411 14403 11462 14430
rect 11681 14464 12383 14523
rect 11681 14430 11699 14464
rect 11733 14430 12331 14464
rect 12365 14430 12383 14464
rect 11681 14369 12383 14430
rect 12417 14497 12475 14514
rect 12417 14463 12429 14497
rect 12463 14463 12475 14497
rect 12417 14369 12475 14463
rect 12748 14460 12797 14531
rect 12748 14426 12757 14460
rect 12791 14426 12797 14460
rect 12748 14410 12797 14426
rect 12841 14460 12943 14476
rect 12875 14426 12909 14460
rect 12841 14369 12943 14426
rect 12979 14471 13017 14644
rect 12979 14437 12981 14471
rect 13015 14437 13017 14471
rect 12979 14403 13017 14437
rect 13051 14607 13106 14635
rect 13051 14573 13073 14607
rect 13051 14565 13106 14573
rect 13085 14531 13106 14565
rect 13051 14403 13106 14531
rect 13147 14565 13181 14675
rect 13147 14515 13181 14531
rect 13215 14517 13249 14743
rect 13283 14617 13317 14811
rect 13351 14837 13385 14879
rect 13351 14769 13385 14803
rect 13351 14701 13385 14735
rect 13351 14651 13385 14667
rect 13419 14837 13486 14845
rect 13419 14803 13435 14837
rect 13469 14803 13486 14837
rect 13419 14769 13486 14803
rect 13419 14735 13435 14769
rect 13469 14735 13486 14769
rect 13419 14701 13486 14735
rect 13419 14667 13435 14701
rect 13469 14667 13486 14701
rect 13419 14651 13486 14667
rect 13283 14601 13322 14617
rect 13283 14567 13288 14601
rect 13283 14551 13322 14567
rect 13367 14601 13418 14617
rect 13367 14567 13384 14601
rect 13367 14551 13418 14567
rect 13367 14517 13401 14551
rect 13452 14517 13486 14651
rect 13521 14837 14223 14879
rect 13521 14803 13539 14837
rect 13573 14803 14171 14837
rect 14205 14803 14223 14837
rect 13521 14735 14223 14803
rect 13521 14701 13539 14735
rect 13573 14701 14171 14735
rect 14205 14701 14223 14735
rect 13521 14661 14223 14701
rect 14275 14829 14309 14845
rect 14275 14761 14309 14795
rect 14345 14829 14411 14879
rect 14345 14795 14361 14829
rect 14395 14795 14411 14829
rect 14345 14761 14411 14795
rect 14345 14727 14361 14761
rect 14395 14727 14411 14761
rect 14445 14829 14499 14845
rect 14445 14795 14447 14829
rect 14481 14795 14499 14829
rect 14619 14837 14680 14879
rect 14445 14748 14499 14795
rect 14275 14693 14309 14727
rect 14445 14714 14447 14748
rect 14481 14743 14499 14748
rect 14445 14709 14453 14714
rect 14487 14709 14499 14743
rect 13521 14591 13859 14661
rect 14275 14659 14408 14693
rect 14445 14664 14499 14709
rect 14374 14630 14408 14659
rect 13521 14557 13599 14591
rect 13633 14557 13702 14591
rect 13736 14557 13805 14591
rect 13839 14557 13859 14591
rect 13893 14593 13913 14627
rect 13947 14593 14012 14627
rect 14046 14593 14111 14627
rect 14145 14593 14223 14627
rect 13893 14523 14223 14593
rect 14261 14607 14327 14623
rect 14261 14573 14269 14607
rect 14303 14601 14327 14607
rect 14261 14567 14277 14573
rect 14311 14567 14327 14601
rect 14261 14549 14327 14567
rect 14374 14614 14431 14630
rect 14374 14580 14397 14614
rect 14374 14564 14431 14580
rect 13215 14483 13401 14517
rect 13215 14476 13250 14483
rect 13144 14460 13250 14476
rect 13178 14426 13250 14460
rect 13435 14471 13486 14517
rect 13435 14464 13441 14471
rect 13144 14403 13250 14426
rect 13335 14445 13401 14449
rect 13335 14411 13351 14445
rect 13385 14411 13401 14445
rect 13335 14369 13401 14411
rect 13475 14437 13486 14471
rect 13469 14430 13486 14437
rect 13435 14403 13486 14430
rect 13521 14464 14223 14523
rect 14374 14513 14408 14564
rect 13521 14430 13539 14464
rect 13573 14430 14171 14464
rect 14205 14430 14223 14464
rect 13521 14369 14223 14430
rect 14275 14479 14408 14513
rect 14465 14504 14499 14664
rect 14275 14458 14309 14479
rect 14447 14475 14499 14504
rect 14275 14403 14309 14424
rect 14345 14411 14361 14445
rect 14395 14411 14411 14445
rect 14345 14369 14411 14411
rect 14481 14441 14499 14475
rect 14447 14403 14499 14441
rect 14534 14801 14585 14817
rect 14534 14767 14551 14801
rect 14534 14733 14585 14767
rect 14534 14699 14551 14733
rect 14534 14641 14585 14699
rect 14619 14803 14635 14837
rect 14669 14803 14680 14837
rect 14748 14837 14814 14879
rect 14748 14803 14764 14837
rect 14798 14803 14814 14837
rect 14918 14837 14968 14879
rect 14850 14811 14884 14827
rect 14619 14769 14680 14803
rect 14918 14803 14934 14837
rect 14918 14787 14968 14803
rect 15002 14836 15176 14845
rect 15002 14802 15126 14836
rect 15160 14802 15176 14836
rect 14850 14769 14884 14777
rect 14619 14735 14635 14769
rect 14669 14735 14680 14769
rect 14619 14651 14680 14735
rect 14724 14735 14884 14769
rect 15002 14777 15176 14802
rect 15223 14829 15257 14845
rect 14534 14511 14576 14641
rect 14724 14617 14758 14735
rect 15002 14701 15036 14777
rect 15223 14753 15257 14795
rect 15291 14837 15365 14879
rect 15291 14803 15311 14837
rect 15345 14803 15365 14837
rect 15492 14827 15558 14879
rect 15673 14835 15809 14845
rect 15291 14787 15365 14803
rect 15424 14811 15458 14827
rect 15492 14793 15508 14827
rect 15542 14793 15558 14827
rect 15605 14811 15639 14827
rect 15424 14759 15458 14777
rect 15605 14759 15639 14777
rect 14792 14667 14808 14701
rect 14842 14667 15036 14701
rect 15070 14717 15117 14743
rect 15070 14683 15086 14717
rect 15151 14709 15162 14743
rect 15223 14719 15335 14753
rect 15424 14725 15639 14759
rect 15673 14801 15759 14835
rect 15793 14801 15809 14835
rect 15673 14779 15809 14801
rect 15852 14829 15902 14845
rect 15886 14795 15902 14829
rect 15852 14779 15902 14795
rect 15936 14837 15986 14879
rect 15970 14803 15986 14837
rect 15936 14787 15986 14803
rect 15120 14685 15162 14709
rect 15301 14691 15335 14719
rect 15120 14683 15263 14685
rect 15002 14649 15036 14667
rect 15128 14651 15263 14683
rect 14610 14611 14758 14617
rect 14610 14601 14793 14611
rect 14644 14567 14793 14601
rect 14610 14551 14793 14567
rect 14728 14516 14793 14551
rect 14534 14495 14585 14511
rect 14534 14471 14551 14495
rect 14534 14437 14545 14471
rect 14729 14461 14793 14516
rect 14827 14602 14935 14633
rect 15002 14615 15083 14649
rect 14827 14593 14901 14602
rect 14827 14559 14885 14593
rect 14919 14559 14935 14568
rect 14971 14565 15015 14581
rect 14827 14539 14875 14559
rect 14827 14505 14841 14539
rect 14971 14531 14981 14565
rect 14971 14525 15015 14531
rect 14827 14479 14875 14505
rect 14909 14491 15015 14525
rect 14579 14437 14585 14461
rect 14534 14405 14585 14437
rect 14619 14445 14680 14461
rect 14619 14411 14635 14445
rect 14669 14411 14680 14445
rect 14729 14427 14759 14461
rect 14909 14445 14943 14491
rect 15049 14459 15083 14615
rect 15117 14607 15187 14617
rect 15151 14591 15187 14607
rect 15117 14557 15125 14573
rect 15159 14557 15187 14591
rect 15117 14493 15187 14557
rect 15221 14543 15263 14651
rect 15255 14509 15263 14543
rect 15221 14493 15263 14509
rect 15301 14657 15551 14691
rect 15585 14657 15601 14691
rect 15301 14519 15335 14657
rect 15673 14623 15707 14779
rect 15868 14753 15902 14779
rect 15369 14603 15707 14623
rect 15403 14589 15707 14603
rect 15741 14743 15834 14745
rect 15775 14717 15834 14743
rect 15868 14719 15947 14753
rect 15775 14709 15800 14717
rect 15741 14683 15800 14709
rect 15741 14667 15834 14683
rect 15369 14553 15403 14569
rect 15437 14521 15465 14555
rect 15499 14539 15595 14555
rect 14793 14427 14943 14445
rect 14729 14411 14943 14427
rect 14977 14441 15015 14457
rect 14619 14369 14680 14411
rect 15011 14407 15015 14441
rect 14977 14369 15015 14407
rect 15049 14445 15239 14459
rect 15049 14411 15189 14445
rect 15223 14411 15239 14445
rect 15301 14441 15353 14519
rect 15437 14505 15489 14521
rect 15523 14505 15561 14539
rect 15049 14403 15239 14411
rect 15283 14407 15299 14441
rect 15333 14407 15353 14441
rect 15395 14445 15461 14461
rect 15395 14411 15411 14445
rect 15445 14411 15461 14445
rect 15636 14447 15670 14589
rect 15741 14549 15775 14667
rect 15704 14515 15720 14549
rect 15754 14515 15775 14549
rect 15704 14505 15775 14515
rect 15809 14607 15879 14629
rect 15809 14573 15833 14607
rect 15867 14573 15879 14607
rect 15809 14555 15879 14573
rect 15809 14521 15822 14555
rect 15856 14521 15879 14555
rect 15809 14505 15879 14521
rect 15913 14447 15947 14719
rect 16020 14685 16085 14842
rect 16119 14829 16153 14845
rect 16119 14761 16153 14795
rect 16187 14813 16253 14879
rect 16187 14779 16203 14813
rect 16237 14779 16253 14813
rect 16287 14829 16338 14845
rect 16321 14795 16338 14829
rect 16287 14761 16338 14795
rect 16466 14837 17535 14879
rect 16466 14803 16483 14837
rect 16517 14803 17483 14837
rect 17517 14803 17535 14837
rect 16466 14792 17535 14803
rect 17569 14808 17627 14879
rect 15981 14662 16073 14685
rect 16015 14628 16073 14662
rect 15981 14539 16073 14628
rect 15981 14505 16017 14539
rect 16051 14505 16073 14539
rect 15981 14475 16073 14505
rect 15636 14413 15757 14447
rect 15791 14413 15807 14447
rect 15848 14413 15864 14447
rect 15898 14413 15947 14447
rect 16119 14471 16153 14709
rect 16188 14727 16287 14745
rect 16321 14727 16338 14761
rect 16188 14711 16338 14727
rect 16188 14616 16234 14711
rect 16222 14607 16234 14616
rect 16188 14573 16200 14582
rect 16188 14513 16234 14573
rect 16268 14607 16338 14677
rect 16268 14601 16293 14607
rect 16268 14567 16290 14601
rect 16327 14573 16338 14607
rect 16324 14567 16338 14573
rect 16268 14547 16338 14567
rect 16784 14591 16854 14792
rect 17569 14774 17581 14808
rect 17615 14774 17627 14808
rect 17754 14837 18823 14879
rect 17754 14803 17771 14837
rect 17805 14803 18771 14837
rect 18805 14803 18823 14837
rect 17754 14792 18823 14803
rect 18858 14837 19927 14879
rect 18858 14803 18875 14837
rect 18909 14803 19875 14837
rect 19909 14803 19927 14837
rect 18858 14792 19927 14803
rect 19961 14837 20203 14879
rect 19961 14803 19979 14837
rect 20013 14803 20151 14837
rect 20185 14803 20203 14837
rect 17569 14715 17627 14774
rect 17569 14681 17581 14715
rect 17615 14681 17627 14715
rect 17569 14646 17627 14681
rect 16784 14557 16803 14591
rect 16837 14557 16854 14591
rect 16784 14542 16854 14557
rect 17150 14627 17218 14644
rect 17150 14593 17167 14627
rect 17201 14593 17218 14627
rect 16188 14479 16338 14513
rect 15395 14369 15461 14411
rect 15981 14407 15997 14441
rect 16031 14407 16047 14441
rect 16287 14471 16338 14479
rect 17150 14478 17218 14593
rect 18072 14591 18142 14792
rect 18072 14557 18091 14591
rect 18125 14557 18142 14591
rect 18072 14542 18142 14557
rect 18438 14627 18506 14644
rect 18438 14593 18455 14627
rect 18489 14593 18506 14627
rect 17569 14497 17627 14514
rect 16119 14421 16153 14437
rect 15981 14369 16047 14407
rect 16187 14411 16203 14445
rect 16237 14411 16253 14445
rect 16321 14437 16338 14471
rect 16287 14421 16338 14437
rect 16466 14464 17535 14478
rect 16466 14430 16483 14464
rect 16517 14430 17483 14464
rect 17517 14430 17535 14464
rect 16187 14369 16253 14411
rect 16466 14369 17535 14430
rect 17569 14463 17581 14497
rect 17615 14463 17627 14497
rect 18438 14478 18506 14593
rect 19176 14591 19246 14792
rect 19961 14742 20203 14803
rect 19961 14708 19979 14742
rect 20013 14708 20151 14742
rect 20185 14708 20203 14742
rect 19961 14661 20203 14708
rect 19176 14557 19195 14591
rect 19229 14557 19246 14591
rect 19176 14542 19246 14557
rect 19542 14627 19610 14644
rect 19542 14593 19559 14627
rect 19593 14593 19610 14627
rect 19542 14478 19610 14593
rect 19961 14587 20065 14661
rect 19961 14553 20011 14587
rect 20045 14553 20065 14587
rect 20099 14593 20119 14627
rect 20153 14593 20203 14627
rect 20099 14519 20203 14593
rect 17569 14369 17627 14463
rect 17754 14464 18823 14478
rect 17754 14430 17771 14464
rect 17805 14430 18771 14464
rect 18805 14430 18823 14464
rect 17754 14369 18823 14430
rect 18858 14464 19927 14478
rect 18858 14430 18875 14464
rect 18909 14430 19875 14464
rect 19909 14430 19927 14464
rect 18858 14369 19927 14430
rect 19961 14466 20203 14519
rect 19961 14432 19979 14466
rect 20013 14432 20151 14466
rect 20185 14432 20203 14466
rect 19961 14369 20203 14432
rect 4948 14335 4977 14369
rect 5011 14335 5069 14369
rect 5103 14335 5161 14369
rect 5195 14335 5253 14369
rect 5287 14335 5345 14369
rect 5379 14335 5437 14369
rect 5471 14335 5529 14369
rect 5563 14335 5621 14369
rect 5655 14335 5713 14369
rect 5747 14335 5805 14369
rect 5839 14335 5897 14369
rect 5931 14335 5989 14369
rect 6023 14335 6081 14369
rect 6115 14335 6173 14369
rect 6207 14335 6265 14369
rect 6299 14335 6357 14369
rect 6391 14335 6449 14369
rect 6483 14335 6541 14369
rect 6575 14335 6633 14369
rect 6667 14335 6725 14369
rect 6759 14335 6817 14369
rect 6851 14335 6909 14369
rect 6943 14335 7001 14369
rect 7035 14335 7093 14369
rect 7127 14335 7185 14369
rect 7219 14335 7277 14369
rect 7311 14335 7369 14369
rect 7403 14335 7461 14369
rect 7495 14335 7553 14369
rect 7587 14335 7645 14369
rect 7679 14335 7737 14369
rect 7771 14335 7829 14369
rect 7863 14335 7921 14369
rect 7955 14335 8013 14369
rect 8047 14335 8105 14369
rect 8139 14335 8197 14369
rect 8231 14335 8289 14369
rect 8323 14335 8381 14369
rect 8415 14335 8473 14369
rect 8507 14335 8565 14369
rect 8599 14335 8657 14369
rect 8691 14335 8749 14369
rect 8783 14335 8841 14369
rect 8875 14335 8933 14369
rect 8967 14335 9025 14369
rect 9059 14335 9117 14369
rect 9151 14335 9209 14369
rect 9243 14335 9301 14369
rect 9335 14335 9393 14369
rect 9427 14335 9485 14369
rect 9519 14335 9577 14369
rect 9611 14335 9669 14369
rect 9703 14335 9761 14369
rect 9795 14335 9853 14369
rect 9887 14335 9945 14369
rect 9979 14335 10037 14369
rect 10071 14335 10129 14369
rect 10163 14335 10221 14369
rect 10255 14335 10313 14369
rect 10347 14335 10405 14369
rect 10439 14335 10497 14369
rect 10531 14335 10589 14369
rect 10623 14335 10681 14369
rect 10715 14335 10773 14369
rect 10807 14335 10865 14369
rect 10899 14335 10957 14369
rect 10991 14335 11049 14369
rect 11083 14335 11141 14369
rect 11175 14335 11233 14369
rect 11267 14335 11325 14369
rect 11359 14335 11417 14369
rect 11451 14335 11509 14369
rect 11543 14335 11601 14369
rect 11635 14335 11693 14369
rect 11727 14335 11785 14369
rect 11819 14335 11877 14369
rect 11911 14335 11969 14369
rect 12003 14335 12061 14369
rect 12095 14335 12153 14369
rect 12187 14335 12245 14369
rect 12279 14335 12337 14369
rect 12371 14335 12429 14369
rect 12463 14335 12521 14369
rect 12555 14335 12613 14369
rect 12647 14335 12705 14369
rect 12739 14335 12797 14369
rect 12831 14335 12889 14369
rect 12923 14335 12981 14369
rect 13015 14335 13073 14369
rect 13107 14335 13165 14369
rect 13199 14335 13257 14369
rect 13291 14335 13349 14369
rect 13383 14335 13441 14369
rect 13475 14335 13533 14369
rect 13567 14335 13625 14369
rect 13659 14335 13717 14369
rect 13751 14335 13809 14369
rect 13843 14335 13901 14369
rect 13935 14335 13993 14369
rect 14027 14335 14085 14369
rect 14119 14335 14177 14369
rect 14211 14335 14269 14369
rect 14303 14335 14361 14369
rect 14395 14335 14453 14369
rect 14487 14335 14545 14369
rect 14579 14335 14637 14369
rect 14671 14335 14729 14369
rect 14763 14335 14821 14369
rect 14855 14335 14913 14369
rect 14947 14335 15005 14369
rect 15039 14335 15097 14369
rect 15131 14335 15189 14369
rect 15223 14335 15281 14369
rect 15315 14335 15373 14369
rect 15407 14335 15465 14369
rect 15499 14335 15557 14369
rect 15591 14335 15649 14369
rect 15683 14335 15741 14369
rect 15775 14335 15833 14369
rect 15867 14335 15925 14369
rect 15959 14335 16017 14369
rect 16051 14335 16109 14369
rect 16143 14335 16201 14369
rect 16235 14335 16293 14369
rect 16327 14335 16385 14369
rect 16419 14335 16477 14369
rect 16511 14335 16569 14369
rect 16603 14335 16661 14369
rect 16695 14335 16753 14369
rect 16787 14335 16845 14369
rect 16879 14335 16937 14369
rect 16971 14335 17029 14369
rect 17063 14335 17121 14369
rect 17155 14335 17213 14369
rect 17247 14335 17305 14369
rect 17339 14335 17397 14369
rect 17431 14335 17489 14369
rect 17523 14335 17581 14369
rect 17615 14335 17673 14369
rect 17707 14335 17765 14369
rect 17799 14335 17857 14369
rect 17891 14335 17949 14369
rect 17983 14335 18041 14369
rect 18075 14335 18133 14369
rect 18167 14335 18225 14369
rect 18259 14335 18317 14369
rect 18351 14335 18409 14369
rect 18443 14335 18501 14369
rect 18535 14335 18593 14369
rect 18627 14335 18685 14369
rect 18719 14335 18777 14369
rect 18811 14335 18869 14369
rect 18903 14335 18961 14369
rect 18995 14335 19053 14369
rect 19087 14335 19145 14369
rect 19179 14335 19237 14369
rect 19271 14335 19329 14369
rect 19363 14335 19421 14369
rect 19455 14335 19513 14369
rect 19547 14335 19605 14369
rect 19639 14335 19697 14369
rect 19731 14335 19789 14369
rect 19823 14335 19881 14369
rect 19915 14335 19973 14369
rect 20007 14335 20065 14369
rect 20099 14335 20157 14369
rect 20191 14335 20220 14369
rect 4965 14272 5207 14335
rect 4965 14238 4983 14272
rect 5017 14238 5155 14272
rect 5189 14238 5207 14272
rect 4965 14185 5207 14238
rect 5426 14274 6495 14335
rect 5426 14240 5443 14274
rect 5477 14240 6443 14274
rect 6477 14240 6495 14274
rect 5426 14226 6495 14240
rect 6530 14274 7599 14335
rect 6530 14240 6547 14274
rect 6581 14240 7547 14274
rect 7581 14240 7599 14274
rect 6530 14226 7599 14240
rect 7634 14274 8703 14335
rect 7634 14240 7651 14274
rect 7685 14240 8651 14274
rect 8685 14240 8703 14274
rect 7634 14226 8703 14240
rect 8738 14274 9807 14335
rect 8738 14240 8755 14274
rect 8789 14240 9755 14274
rect 9789 14240 9807 14274
rect 8738 14226 9807 14240
rect 9841 14241 9899 14335
rect 4965 14111 5069 14185
rect 4965 14077 5015 14111
rect 5049 14077 5069 14111
rect 5103 14117 5123 14151
rect 5157 14117 5207 14151
rect 5103 14043 5207 14117
rect 4965 13996 5207 14043
rect 4965 13962 4983 13996
rect 5017 13962 5155 13996
rect 5189 13962 5207 13996
rect 4965 13901 5207 13962
rect 5744 14147 5814 14162
rect 5744 14113 5763 14147
rect 5797 14113 5814 14147
rect 5744 13912 5814 14113
rect 6110 14111 6178 14226
rect 6110 14077 6127 14111
rect 6161 14077 6178 14111
rect 6110 14060 6178 14077
rect 6848 14147 6918 14162
rect 6848 14113 6867 14147
rect 6901 14113 6918 14147
rect 6848 13912 6918 14113
rect 7214 14111 7282 14226
rect 7214 14077 7231 14111
rect 7265 14077 7282 14111
rect 7214 14060 7282 14077
rect 7952 14147 8022 14162
rect 7952 14113 7971 14147
rect 8005 14113 8022 14147
rect 7952 13912 8022 14113
rect 8318 14111 8386 14226
rect 8318 14077 8335 14111
rect 8369 14077 8386 14111
rect 8318 14060 8386 14077
rect 9056 14147 9126 14162
rect 9056 14113 9075 14147
rect 9109 14113 9126 14147
rect 9056 13912 9126 14113
rect 9422 14111 9490 14226
rect 9841 14207 9853 14241
rect 9887 14207 9899 14241
rect 9841 14190 9899 14207
rect 10118 14243 10169 14299
rect 10203 14293 10264 14335
rect 10561 14297 10599 14335
rect 10203 14259 10219 14293
rect 10253 14259 10264 14293
rect 10203 14243 10264 14259
rect 10313 14277 10527 14293
rect 10313 14243 10343 14277
rect 10377 14259 10527 14277
rect 10118 14209 10135 14243
rect 10118 14193 10169 14209
rect 9422 14077 9439 14111
rect 9473 14077 9490 14111
rect 9422 14060 9490 14077
rect 10118 14063 10160 14193
rect 10313 14188 10377 14243
rect 10312 14153 10377 14188
rect 10194 14137 10377 14153
rect 10228 14103 10377 14137
rect 10194 14093 10377 14103
rect 10411 14199 10459 14225
rect 10411 14165 10425 14199
rect 10493 14213 10527 14259
rect 10595 14263 10599 14297
rect 10561 14247 10599 14263
rect 10633 14293 10823 14301
rect 10633 14259 10773 14293
rect 10807 14259 10823 14293
rect 10867 14263 10883 14297
rect 10917 14263 10937 14297
rect 10633 14245 10823 14259
rect 10493 14179 10599 14213
rect 10411 14145 10459 14165
rect 10555 14173 10599 14179
rect 10411 14111 10469 14145
rect 10503 14136 10519 14145
rect 10555 14139 10565 14173
rect 10555 14123 10599 14139
rect 10411 14102 10485 14111
rect 10194 14087 10342 14093
rect 9841 14023 9899 14058
rect 9841 13989 9853 14023
rect 9887 13989 9899 14023
rect 9841 13930 9899 13989
rect 4965 13867 4983 13901
rect 5017 13867 5155 13901
rect 5189 13867 5207 13901
rect 4965 13825 5207 13867
rect 5426 13901 6495 13912
rect 5426 13867 5443 13901
rect 5477 13867 6443 13901
rect 6477 13867 6495 13901
rect 5426 13825 6495 13867
rect 6530 13901 7599 13912
rect 6530 13867 6547 13901
rect 6581 13867 7547 13901
rect 7581 13867 7599 13901
rect 6530 13825 7599 13867
rect 7634 13901 8703 13912
rect 7634 13867 7651 13901
rect 7685 13867 8651 13901
rect 8685 13867 8703 13901
rect 7634 13825 8703 13867
rect 8738 13901 9807 13912
rect 8738 13867 8755 13901
rect 8789 13867 9755 13901
rect 9789 13867 9807 13901
rect 8738 13825 9807 13867
rect 9841 13896 9853 13930
rect 9887 13896 9899 13930
rect 9841 13825 9899 13896
rect 10118 14005 10169 14063
rect 10118 13971 10135 14005
rect 10118 13937 10169 13971
rect 10118 13927 10135 13937
rect 10118 13893 10129 13927
rect 10163 13893 10169 13903
rect 10118 13887 10169 13893
rect 10203 13969 10264 14053
rect 10203 13935 10219 13969
rect 10253 13935 10264 13969
rect 10308 13969 10342 14087
rect 10411 14071 10519 14102
rect 10633 14089 10667 14245
rect 10586 14055 10667 14089
rect 10701 14147 10771 14211
rect 10701 14131 10709 14147
rect 10743 14113 10771 14147
rect 10735 14097 10771 14113
rect 10701 14087 10771 14097
rect 10805 14195 10847 14211
rect 10839 14161 10847 14195
rect 10586 14037 10620 14055
rect 10805 14053 10847 14161
rect 10376 14003 10392 14037
rect 10426 14003 10620 14037
rect 10712 14021 10847 14053
rect 10308 13935 10468 13969
rect 10203 13901 10264 13935
rect 10434 13927 10468 13935
rect 10203 13867 10219 13901
rect 10253 13867 10264 13901
rect 10203 13825 10264 13867
rect 10332 13867 10348 13901
rect 10382 13867 10398 13901
rect 10586 13927 10620 14003
rect 10654 13987 10670 14021
rect 10704 14019 10847 14021
rect 10885 14185 10937 14263
rect 10979 14293 11045 14335
rect 10979 14259 10995 14293
rect 11029 14259 11045 14293
rect 11565 14297 11631 14335
rect 10979 14243 11045 14259
rect 11220 14257 11341 14291
rect 11375 14257 11391 14291
rect 11432 14257 11448 14291
rect 11482 14257 11531 14291
rect 11565 14263 11581 14297
rect 11615 14263 11631 14297
rect 11771 14293 11837 14335
rect 11703 14267 11737 14283
rect 10885 14047 10919 14185
rect 11021 14183 11073 14199
rect 10953 14135 10987 14151
rect 11021 14149 11049 14183
rect 11107 14165 11145 14199
rect 11083 14149 11179 14165
rect 11220 14115 11254 14257
rect 11288 14189 11359 14199
rect 11288 14155 11304 14189
rect 11338 14155 11359 14189
rect 10987 14101 11291 14115
rect 10953 14081 11291 14101
rect 10704 13995 10746 14019
rect 10654 13961 10701 13987
rect 10735 13961 10746 13995
rect 10885 14013 11135 14047
rect 11169 14013 11185 14047
rect 10885 13985 10919 14013
rect 10807 13951 10919 13985
rect 10434 13877 10468 13893
rect 10502 13901 10552 13917
rect 10332 13825 10398 13867
rect 10502 13867 10518 13901
rect 10502 13825 10552 13867
rect 10586 13902 10760 13927
rect 10586 13868 10710 13902
rect 10744 13868 10760 13902
rect 10586 13859 10760 13868
rect 10807 13909 10841 13951
rect 11008 13945 11223 13979
rect 11008 13927 11042 13945
rect 10807 13859 10841 13875
rect 10875 13901 10949 13917
rect 10875 13867 10895 13901
rect 10929 13867 10949 13901
rect 11189 13927 11223 13945
rect 11008 13877 11042 13893
rect 11076 13877 11092 13911
rect 11126 13877 11142 13911
rect 11189 13877 11223 13893
rect 11257 13925 11291 14081
rect 11325 14037 11359 14155
rect 11393 14183 11463 14199
rect 11393 14149 11406 14183
rect 11440 14149 11463 14183
rect 11393 14131 11463 14149
rect 11393 14097 11417 14131
rect 11451 14097 11463 14131
rect 11393 14075 11463 14097
rect 11325 14021 11418 14037
rect 11325 13995 11384 14021
rect 11359 13987 11384 13995
rect 11359 13961 11418 13987
rect 11497 13985 11531 14257
rect 11771 14259 11787 14293
rect 11821 14259 11837 14293
rect 11871 14267 11922 14283
rect 11565 14076 11657 14229
rect 11599 14063 11657 14076
rect 11599 14042 11601 14063
rect 11565 14029 11601 14042
rect 11635 14029 11657 14063
rect 11565 14019 11657 14029
rect 11325 13959 11418 13961
rect 11452 13951 11531 13985
rect 11452 13925 11486 13951
rect 11257 13903 11393 13925
rect 10875 13825 10949 13867
rect 11076 13825 11142 13877
rect 11257 13869 11343 13903
rect 11377 13869 11393 13903
rect 11257 13859 11393 13869
rect 11436 13909 11486 13925
rect 11470 13875 11486 13909
rect 11436 13859 11486 13875
rect 11520 13901 11570 13917
rect 11554 13867 11570 13901
rect 11520 13825 11570 13867
rect 11604 13862 11669 14019
rect 11703 13995 11737 14233
rect 11905 14233 11922 14267
rect 11871 14225 11922 14233
rect 11772 14191 11922 14225
rect 11957 14263 12009 14301
rect 11957 14229 11975 14263
rect 12045 14293 12111 14335
rect 12045 14259 12061 14293
rect 12095 14259 12111 14293
rect 12147 14280 12181 14301
rect 11957 14200 12009 14229
rect 12147 14225 12181 14246
rect 12251 14289 12311 14335
rect 12251 14255 12268 14289
rect 12302 14255 12311 14289
rect 12251 14239 12311 14255
rect 12345 14280 12397 14296
rect 12345 14246 12354 14280
rect 12388 14246 12397 14280
rect 11772 14131 11818 14191
rect 11772 14122 11784 14131
rect 11806 14088 11818 14097
rect 11772 13993 11818 14088
rect 11852 14137 11922 14157
rect 11852 14103 11874 14137
rect 11908 14103 11922 14137
rect 11852 14063 11922 14103
rect 11852 14029 11877 14063
rect 11911 14029 11922 14063
rect 11852 14027 11922 14029
rect 11957 14040 11991 14200
rect 12048 14191 12181 14225
rect 12345 14205 12397 14246
rect 12431 14289 12483 14335
rect 12431 14255 12440 14289
rect 12474 14255 12483 14289
rect 12431 14239 12483 14255
rect 12519 14280 12571 14296
rect 12519 14246 12526 14280
rect 12560 14246 12571 14280
rect 12519 14205 12571 14246
rect 12605 14289 12655 14335
rect 12605 14255 12612 14289
rect 12646 14255 12655 14289
rect 12605 14239 12655 14255
rect 12691 14280 12743 14296
rect 12691 14246 12698 14280
rect 12732 14246 12743 14280
rect 12691 14205 12743 14246
rect 12777 14289 12827 14335
rect 12777 14255 12784 14289
rect 12818 14255 12827 14289
rect 12777 14239 12827 14255
rect 12863 14280 12915 14296
rect 12863 14246 12870 14280
rect 12904 14246 12915 14280
rect 12863 14205 12915 14246
rect 12949 14289 12998 14335
rect 12949 14255 12955 14289
rect 12989 14255 12998 14289
rect 12949 14239 12998 14255
rect 13032 14280 13087 14296
rect 13032 14246 13041 14280
rect 13075 14246 13087 14280
rect 13032 14205 13087 14246
rect 13121 14289 13170 14335
rect 13121 14255 13127 14289
rect 13161 14255 13170 14289
rect 13121 14239 13170 14255
rect 13204 14280 13256 14296
rect 13204 14246 13213 14280
rect 13247 14246 13256 14280
rect 13204 14205 13256 14246
rect 13290 14289 13342 14335
rect 13290 14255 13299 14289
rect 13333 14255 13342 14289
rect 13290 14239 13342 14255
rect 13376 14280 13428 14296
rect 13376 14246 13385 14280
rect 13419 14246 13428 14280
rect 13376 14205 13428 14246
rect 13462 14289 13514 14335
rect 13462 14255 13471 14289
rect 13505 14255 13514 14289
rect 13462 14239 13514 14255
rect 13548 14280 13600 14296
rect 13548 14246 13557 14280
rect 13591 14246 13600 14280
rect 13548 14205 13600 14246
rect 13634 14280 13686 14335
rect 13634 14246 13643 14280
rect 13677 14246 13686 14280
rect 13634 14223 13686 14246
rect 13720 14280 13770 14299
rect 13720 14246 13729 14280
rect 13763 14246 13770 14280
rect 12048 14140 12082 14191
rect 12251 14171 13600 14205
rect 12025 14124 12082 14140
rect 12059 14090 12082 14124
rect 12025 14074 12082 14090
rect 12129 14137 12195 14155
rect 12129 14103 12145 14137
rect 12179 14131 12195 14137
rect 12129 14097 12153 14103
rect 12187 14097 12195 14131
rect 12129 14081 12195 14097
rect 12048 14045 12082 14074
rect 12251 14053 12484 14171
rect 13720 14137 13770 14246
rect 13806 14280 13858 14335
rect 13806 14246 13815 14280
rect 13849 14246 13858 14280
rect 13806 14230 13858 14246
rect 13892 14280 13942 14299
rect 13892 14246 13901 14280
rect 13935 14246 13942 14280
rect 13892 14137 13942 14246
rect 13978 14293 14039 14335
rect 13978 14259 13987 14293
rect 14021 14259 14039 14293
rect 13978 14233 14039 14259
rect 14280 14267 14337 14301
rect 14280 14233 14297 14267
rect 14331 14233 14337 14267
rect 14371 14293 14425 14335
rect 14371 14259 14381 14293
rect 14415 14259 14425 14293
rect 14371 14243 14425 14259
rect 14505 14267 14585 14301
rect 14280 14209 14337 14233
rect 14505 14233 14535 14267
rect 14569 14233 14585 14267
rect 12518 14103 12538 14137
rect 12572 14103 12606 14137
rect 12640 14103 12674 14137
rect 12708 14103 12742 14137
rect 12776 14103 12810 14137
rect 12844 14103 12878 14137
rect 12912 14103 12946 14137
rect 12980 14103 13014 14137
rect 13048 14103 13082 14137
rect 13116 14103 13150 14137
rect 13184 14103 13218 14137
rect 13252 14103 13286 14137
rect 13320 14103 13354 14137
rect 13388 14103 13422 14137
rect 13456 14103 13490 14137
rect 13524 14103 13558 14137
rect 13592 14103 13942 14137
rect 12518 14087 13942 14103
rect 13976 14165 13993 14199
rect 14027 14165 14039 14199
rect 14280 14175 14471 14209
rect 13976 14137 14039 14165
rect 13976 14103 13985 14137
rect 14019 14103 14039 14137
rect 13976 14087 14039 14103
rect 14257 14137 14395 14141
rect 14257 14103 14321 14137
rect 14355 14103 14395 14137
rect 11957 13995 12011 14040
rect 12048 14011 12181 14045
rect 11772 13977 11922 13993
rect 11772 13959 11871 13977
rect 11703 13909 11737 13943
rect 11905 13943 11922 13977
rect 11703 13859 11737 13875
rect 11771 13891 11787 13925
rect 11821 13891 11837 13925
rect 11771 13825 11837 13891
rect 11871 13909 11922 13943
rect 11905 13875 11922 13909
rect 11871 13859 11922 13875
rect 11957 13961 11969 13995
rect 12003 13990 12011 13995
rect 11957 13956 11975 13961
rect 12009 13956 12011 13990
rect 12147 13977 12181 14011
rect 12251 14031 13600 14053
rect 12251 14008 12354 14031
rect 11957 13909 12011 13956
rect 11957 13875 11975 13909
rect 12009 13875 12011 13909
rect 11957 13859 12011 13875
rect 12045 13943 12061 13977
rect 12095 13943 12111 13977
rect 12045 13909 12111 13943
rect 12045 13875 12061 13909
rect 12095 13875 12111 13909
rect 12045 13825 12111 13875
rect 12339 13997 12354 14008
rect 12388 14008 12526 14031
rect 12388 13997 12397 14008
rect 12147 13909 12181 13943
rect 12147 13859 12181 13875
rect 12251 13925 12305 13974
rect 12251 13891 12268 13925
rect 12302 13891 12305 13925
rect 12251 13825 12305 13891
rect 12339 13945 12397 13997
rect 12519 13997 12526 14008
rect 12560 14005 12698 14031
rect 12560 13997 12571 14005
rect 12339 13911 12354 13945
rect 12388 13911 12397 13945
rect 12339 13860 12397 13911
rect 12431 13925 12482 13971
rect 12431 13891 12440 13925
rect 12474 13891 12482 13925
rect 12431 13826 12482 13891
rect 12519 13945 12571 13997
rect 12691 13997 12698 14005
rect 12732 14005 12870 14031
rect 12732 13997 12743 14005
rect 12519 13911 12526 13945
rect 12560 13911 12571 13945
rect 12519 13860 12571 13911
rect 12605 13925 12654 13971
rect 12605 13891 12612 13925
rect 12646 13891 12654 13925
rect 12605 13826 12654 13891
rect 12691 13945 12743 13997
rect 12863 13997 12870 14005
rect 12904 14005 13041 14031
rect 12904 13997 12915 14005
rect 12691 13911 12698 13945
rect 12732 13927 12743 13945
rect 12691 13893 12705 13911
rect 12739 13893 12743 13927
rect 12691 13860 12743 13893
rect 12777 13925 12826 13971
rect 12777 13891 12784 13925
rect 12818 13891 12826 13925
rect 12777 13826 12826 13891
rect 12863 13945 12915 13997
rect 13032 13997 13041 14005
rect 13075 14005 13213 14031
rect 13075 13997 13084 14005
rect 12863 13911 12870 13945
rect 12904 13911 12915 13945
rect 12863 13860 12915 13911
rect 12949 13925 12998 13971
rect 12949 13891 12955 13925
rect 12989 13891 12998 13925
rect 12949 13826 12998 13891
rect 13032 13945 13084 13997
rect 13204 13997 13213 14005
rect 13247 14005 13385 14031
rect 13247 13997 13256 14005
rect 13032 13911 13041 13945
rect 13075 13911 13084 13945
rect 13032 13860 13084 13911
rect 13118 13925 13170 13971
rect 13118 13891 13127 13925
rect 13161 13891 13170 13925
rect 13118 13826 13170 13891
rect 13204 13945 13256 13997
rect 13376 13997 13385 14005
rect 13419 14005 13557 14031
rect 13419 13997 13428 14005
rect 13204 13911 13213 13945
rect 13247 13911 13256 13945
rect 13204 13860 13256 13911
rect 13290 13925 13342 13971
rect 13290 13891 13299 13925
rect 13333 13891 13342 13925
rect 13290 13826 13342 13891
rect 13376 13945 13428 13997
rect 13548 13997 13557 14005
rect 13591 13997 13600 14031
rect 13376 13911 13385 13945
rect 13419 13911 13428 13945
rect 13376 13860 13428 13911
rect 13462 13925 13514 13971
rect 13462 13891 13471 13925
rect 13505 13891 13514 13925
rect 13462 13826 13514 13891
rect 13548 13945 13600 13997
rect 13720 13985 13770 14087
rect 13548 13911 13557 13945
rect 13591 13911 13600 13945
rect 13548 13860 13600 13911
rect 13634 13969 13686 13985
rect 13634 13935 13643 13969
rect 13677 13935 13686 13969
rect 13634 13901 13686 13935
rect 13634 13867 13643 13901
rect 13677 13867 13686 13901
rect 13634 13826 13686 13867
rect 13720 13951 13729 13985
rect 13763 13951 13770 13985
rect 13720 13917 13770 13951
rect 13720 13883 13729 13917
rect 13763 13883 13770 13917
rect 13720 13860 13770 13883
rect 13806 13969 13858 13987
rect 13806 13935 13815 13969
rect 13849 13935 13858 13969
rect 13806 13901 13858 13935
rect 13806 13867 13815 13901
rect 13849 13867 13858 13901
rect 12431 13825 13686 13826
rect 13806 13825 13858 13867
rect 13893 13977 13942 14087
rect 14257 14063 14395 14103
rect 14257 14029 14269 14063
rect 14303 14029 14395 14063
rect 14429 14137 14471 14175
rect 14429 14103 14435 14137
rect 14469 14103 14471 14137
rect 14429 13995 14471 14103
rect 13893 13943 13901 13977
rect 13935 13943 13942 13977
rect 13893 13909 13942 13943
rect 13893 13875 13901 13909
rect 13935 13875 13942 13909
rect 13893 13859 13942 13875
rect 13978 13969 14037 13987
rect 13978 13935 13987 13969
rect 14021 13935 14037 13969
rect 13978 13901 14037 13935
rect 13978 13867 13987 13901
rect 14021 13867 14037 13901
rect 13978 13825 14037 13867
rect 14280 13951 14471 13995
rect 14505 14141 14585 14233
rect 14623 14267 14679 14301
rect 14623 14233 14639 14267
rect 14673 14233 14679 14267
rect 14783 14293 14848 14335
rect 14783 14259 14798 14293
rect 14832 14259 14848 14293
rect 14783 14243 14848 14259
rect 14882 14267 14959 14301
rect 14623 14209 14679 14233
rect 14882 14233 14888 14267
rect 14922 14233 14959 14267
rect 14623 14175 14848 14209
rect 14882 14187 14959 14233
rect 14993 14241 15051 14335
rect 14993 14207 15005 14241
rect 15039 14207 15051 14241
rect 14993 14190 15051 14207
rect 15178 14274 15229 14301
rect 15178 14267 15195 14274
rect 15178 14233 15189 14267
rect 15263 14293 15329 14335
rect 15263 14259 15279 14293
rect 15313 14259 15329 14293
rect 15263 14255 15329 14259
rect 15414 14278 15520 14301
rect 15223 14233 15229 14240
rect 14758 14153 14848 14175
rect 14505 14137 14724 14141
rect 14505 14103 14639 14137
rect 14673 14103 14724 14137
rect 14505 14029 14724 14103
rect 14758 14137 14869 14153
rect 14758 14103 14835 14137
rect 14758 14087 14869 14103
rect 14903 14131 14959 14187
rect 14903 14097 14913 14131
rect 14947 14097 14959 14131
rect 14280 13927 14337 13951
rect 14280 13893 14297 13927
rect 14331 13893 14337 13927
rect 14505 13927 14585 14029
rect 14758 13995 14848 14087
rect 14903 14053 14959 14097
rect 15178 14187 15229 14233
rect 15414 14244 15486 14278
rect 15414 14228 15520 14244
rect 15414 14221 15449 14228
rect 15263 14187 15449 14221
rect 14280 13859 14337 13893
rect 14371 13901 14425 13917
rect 14371 13867 14381 13901
rect 14415 13867 14425 13901
rect 14371 13825 14425 13867
rect 14505 13893 14535 13927
rect 14569 13893 14585 13927
rect 14505 13859 14585 13893
rect 14623 13951 14848 13995
rect 14623 13927 14679 13951
rect 14623 13893 14639 13927
rect 14673 13893 14679 13927
rect 14882 13927 14959 14053
rect 14623 13859 14679 13893
rect 14783 13901 14848 13917
rect 14783 13867 14798 13901
rect 14832 13867 14848 13901
rect 14783 13825 14848 13867
rect 14882 13893 14888 13927
rect 14922 13893 14959 13927
rect 14882 13859 14959 13893
rect 14993 14023 15051 14058
rect 14993 13989 15005 14023
rect 15039 13989 15051 14023
rect 14993 13930 15051 13989
rect 14993 13896 15005 13930
rect 15039 13896 15051 13930
rect 14993 13825 15051 13896
rect 15178 14053 15212 14187
rect 15263 14153 15297 14187
rect 15246 14137 15297 14153
rect 15280 14103 15297 14137
rect 15246 14087 15297 14103
rect 15342 14137 15381 14153
rect 15376 14103 15381 14137
rect 15342 14087 15381 14103
rect 15178 14037 15245 14053
rect 15178 14003 15195 14037
rect 15229 14003 15245 14037
rect 15178 13969 15245 14003
rect 15178 13935 15195 13969
rect 15229 13935 15245 13969
rect 15178 13901 15245 13935
rect 15178 13867 15195 13901
rect 15229 13867 15245 13901
rect 15178 13859 15245 13867
rect 15279 14037 15313 14053
rect 15279 13969 15313 14003
rect 15279 13901 15313 13935
rect 15279 13825 15313 13867
rect 15347 13893 15381 14087
rect 15415 13961 15449 14187
rect 15483 14173 15517 14189
rect 15483 14029 15517 14139
rect 15558 14173 15613 14301
rect 15558 14139 15579 14173
rect 15558 14131 15613 14139
rect 15591 14097 15613 14131
rect 15558 14069 15613 14097
rect 15647 14267 15685 14301
rect 15647 14233 15649 14267
rect 15683 14233 15685 14267
rect 15647 14060 15685 14233
rect 15721 14278 15823 14335
rect 15755 14244 15789 14278
rect 15721 14228 15823 14244
rect 15867 14278 15916 14294
rect 15867 14244 15873 14278
rect 15907 14244 15916 14278
rect 15867 14173 15916 14244
rect 16005 14267 16057 14301
rect 16005 14233 16017 14267
rect 16051 14263 16057 14267
rect 16093 14293 16159 14335
rect 16093 14259 16109 14293
rect 16143 14259 16159 14293
rect 16195 14280 16229 14301
rect 16005 14229 16023 14233
rect 16005 14200 16057 14229
rect 16195 14225 16229 14246
rect 15725 14139 15741 14173
rect 15775 14139 15971 14173
rect 15647 14029 15651 14060
rect 15483 14026 15651 14029
rect 15483 13995 15685 14026
rect 15719 14063 15869 14064
rect 15719 14060 15833 14063
rect 15719 14026 15819 14060
rect 15867 14029 15869 14063
rect 15853 14026 15869 14029
rect 15415 13927 15515 13961
rect 15549 13927 15590 13961
rect 15624 13927 15640 13961
rect 15719 13893 15753 14026
rect 15903 13977 15971 14139
rect 15347 13859 15753 13893
rect 15787 13961 15821 13977
rect 15787 13825 15821 13927
rect 15868 13961 15971 13977
rect 15868 13927 15873 13961
rect 15907 13927 15971 13961
rect 15868 13895 15971 13927
rect 16005 14040 16039 14200
rect 16096 14191 16229 14225
rect 16281 14263 16333 14301
rect 16281 14229 16299 14263
rect 16369 14293 16435 14335
rect 16369 14259 16385 14293
rect 16419 14259 16435 14293
rect 16471 14280 16505 14301
rect 16281 14200 16333 14229
rect 16471 14225 16505 14246
rect 16650 14274 17719 14335
rect 16650 14240 16667 14274
rect 16701 14240 17667 14274
rect 17701 14240 17719 14274
rect 16650 14226 17719 14240
rect 17754 14274 18823 14335
rect 17754 14240 17771 14274
rect 17805 14240 18771 14274
rect 18805 14240 18823 14274
rect 17754 14226 18823 14240
rect 18858 14274 19927 14335
rect 18858 14240 18875 14274
rect 18909 14240 19875 14274
rect 19909 14240 19927 14274
rect 18858 14226 19927 14240
rect 19961 14272 20203 14335
rect 19961 14238 19979 14272
rect 20013 14238 20151 14272
rect 20185 14238 20203 14272
rect 16096 14140 16130 14191
rect 16073 14124 16130 14140
rect 16107 14090 16130 14124
rect 16073 14074 16130 14090
rect 16177 14137 16243 14155
rect 16177 14103 16193 14137
rect 16227 14131 16243 14137
rect 16177 14097 16201 14103
rect 16235 14097 16243 14131
rect 16177 14081 16243 14097
rect 16096 14045 16130 14074
rect 16005 13990 16059 14040
rect 16096 14011 16229 14045
rect 16005 13956 16023 13990
rect 16057 13956 16059 13990
rect 16195 13977 16229 14011
rect 16005 13909 16059 13956
rect 16005 13875 16023 13909
rect 16057 13875 16059 13909
rect 16005 13859 16059 13875
rect 16093 13943 16109 13977
rect 16143 13943 16159 13977
rect 16093 13909 16159 13943
rect 16093 13875 16109 13909
rect 16143 13875 16159 13909
rect 16093 13825 16159 13875
rect 16195 13909 16229 13943
rect 16195 13859 16229 13875
rect 16281 14040 16315 14200
rect 16372 14191 16505 14225
rect 16372 14140 16406 14191
rect 16349 14124 16406 14140
rect 16383 14090 16406 14124
rect 16349 14074 16406 14090
rect 16453 14137 16519 14155
rect 16453 14103 16469 14137
rect 16503 14131 16519 14137
rect 16453 14097 16477 14103
rect 16511 14097 16519 14131
rect 16453 14081 16519 14097
rect 16968 14147 17038 14162
rect 16968 14113 16987 14147
rect 17021 14113 17038 14147
rect 16372 14045 16406 14074
rect 16281 13990 16335 14040
rect 16372 14011 16505 14045
rect 16281 13956 16299 13990
rect 16333 13956 16335 13990
rect 16471 13977 16505 14011
rect 16281 13927 16335 13956
rect 16281 13893 16293 13927
rect 16327 13909 16335 13927
rect 16281 13875 16299 13893
rect 16333 13875 16335 13909
rect 16281 13859 16335 13875
rect 16369 13943 16385 13977
rect 16419 13943 16435 13977
rect 16369 13909 16435 13943
rect 16369 13875 16385 13909
rect 16419 13875 16435 13909
rect 16369 13825 16435 13875
rect 16471 13909 16505 13943
rect 16968 13912 17038 14113
rect 17334 14111 17402 14226
rect 17334 14077 17351 14111
rect 17385 14077 17402 14111
rect 17334 14060 17402 14077
rect 18072 14147 18142 14162
rect 18072 14113 18091 14147
rect 18125 14113 18142 14147
rect 18072 13912 18142 14113
rect 18438 14111 18506 14226
rect 18438 14077 18455 14111
rect 18489 14077 18506 14111
rect 18438 14060 18506 14077
rect 19176 14147 19246 14162
rect 19176 14113 19195 14147
rect 19229 14113 19246 14147
rect 19176 13912 19246 14113
rect 19542 14111 19610 14226
rect 19961 14185 20203 14238
rect 19542 14077 19559 14111
rect 19593 14077 19610 14111
rect 19542 14060 19610 14077
rect 19961 14117 20011 14151
rect 20045 14117 20065 14151
rect 19961 14043 20065 14117
rect 20099 14111 20203 14185
rect 20099 14077 20119 14111
rect 20153 14077 20203 14111
rect 19961 13996 20203 14043
rect 19961 13962 19979 13996
rect 20013 13962 20151 13996
rect 20185 13962 20203 13996
rect 16471 13859 16505 13875
rect 16650 13901 17719 13912
rect 16650 13867 16667 13901
rect 16701 13867 17667 13901
rect 17701 13867 17719 13901
rect 16650 13825 17719 13867
rect 17754 13901 18823 13912
rect 17754 13867 17771 13901
rect 17805 13867 18771 13901
rect 18805 13867 18823 13901
rect 17754 13825 18823 13867
rect 18858 13901 19927 13912
rect 18858 13867 18875 13901
rect 18909 13867 19875 13901
rect 19909 13867 19927 13901
rect 18858 13825 19927 13867
rect 19961 13901 20203 13962
rect 19961 13867 19979 13901
rect 20013 13867 20151 13901
rect 20185 13867 20203 13901
rect 19961 13825 20203 13867
rect 4948 13791 4977 13825
rect 5011 13791 5069 13825
rect 5103 13791 5161 13825
rect 5195 13791 5253 13825
rect 5287 13791 5345 13825
rect 5379 13791 5437 13825
rect 5471 13791 5529 13825
rect 5563 13791 5621 13825
rect 5655 13791 5713 13825
rect 5747 13791 5805 13825
rect 5839 13791 5897 13825
rect 5931 13791 5989 13825
rect 6023 13791 6081 13825
rect 6115 13791 6173 13825
rect 6207 13791 6265 13825
rect 6299 13791 6357 13825
rect 6391 13791 6449 13825
rect 6483 13791 6541 13825
rect 6575 13791 6633 13825
rect 6667 13791 6725 13825
rect 6759 13791 6817 13825
rect 6851 13791 6909 13825
rect 6943 13791 7001 13825
rect 7035 13791 7093 13825
rect 7127 13791 7185 13825
rect 7219 13791 7277 13825
rect 7311 13791 7369 13825
rect 7403 13791 7461 13825
rect 7495 13791 7553 13825
rect 7587 13791 7645 13825
rect 7679 13791 7737 13825
rect 7771 13791 7829 13825
rect 7863 13791 7921 13825
rect 7955 13791 8013 13825
rect 8047 13791 8105 13825
rect 8139 13791 8197 13825
rect 8231 13791 8289 13825
rect 8323 13791 8381 13825
rect 8415 13791 8473 13825
rect 8507 13791 8565 13825
rect 8599 13791 8657 13825
rect 8691 13791 8749 13825
rect 8783 13791 8841 13825
rect 8875 13791 8933 13825
rect 8967 13791 9025 13825
rect 9059 13791 9117 13825
rect 9151 13791 9209 13825
rect 9243 13791 9301 13825
rect 9335 13791 9393 13825
rect 9427 13791 9485 13825
rect 9519 13791 9577 13825
rect 9611 13791 9669 13825
rect 9703 13791 9761 13825
rect 9795 13791 9853 13825
rect 9887 13791 9945 13825
rect 9979 13791 10037 13825
rect 10071 13791 10129 13825
rect 10163 13791 10221 13825
rect 10255 13791 10313 13825
rect 10347 13791 10405 13825
rect 10439 13791 10497 13825
rect 10531 13791 10589 13825
rect 10623 13791 10681 13825
rect 10715 13791 10773 13825
rect 10807 13791 10865 13825
rect 10899 13791 10957 13825
rect 10991 13791 11049 13825
rect 11083 13791 11141 13825
rect 11175 13791 11233 13825
rect 11267 13791 11325 13825
rect 11359 13791 11417 13825
rect 11451 13791 11509 13825
rect 11543 13791 11601 13825
rect 11635 13791 11693 13825
rect 11727 13791 11785 13825
rect 11819 13791 11877 13825
rect 11911 13791 11969 13825
rect 12003 13791 12061 13825
rect 12095 13791 12153 13825
rect 12187 13791 12245 13825
rect 12279 13791 12337 13825
rect 12371 13791 12429 13825
rect 12463 13791 12521 13825
rect 12555 13791 12613 13825
rect 12647 13791 12705 13825
rect 12739 13791 12797 13825
rect 12831 13791 12889 13825
rect 12923 13791 12981 13825
rect 13015 13791 13073 13825
rect 13107 13791 13165 13825
rect 13199 13791 13257 13825
rect 13291 13791 13349 13825
rect 13383 13791 13441 13825
rect 13475 13791 13533 13825
rect 13567 13791 13625 13825
rect 13659 13791 13717 13825
rect 13751 13791 13809 13825
rect 13843 13791 13901 13825
rect 13935 13791 13993 13825
rect 14027 13791 14085 13825
rect 14119 13791 14177 13825
rect 14211 13791 14269 13825
rect 14303 13791 14361 13825
rect 14395 13791 14453 13825
rect 14487 13791 14545 13825
rect 14579 13791 14637 13825
rect 14671 13791 14729 13825
rect 14763 13791 14821 13825
rect 14855 13791 14913 13825
rect 14947 13791 15005 13825
rect 15039 13791 15097 13825
rect 15131 13791 15189 13825
rect 15223 13791 15281 13825
rect 15315 13791 15373 13825
rect 15407 13791 15465 13825
rect 15499 13791 15557 13825
rect 15591 13791 15649 13825
rect 15683 13791 15741 13825
rect 15775 13791 15833 13825
rect 15867 13791 15925 13825
rect 15959 13791 16017 13825
rect 16051 13791 16109 13825
rect 16143 13791 16201 13825
rect 16235 13791 16293 13825
rect 16327 13791 16385 13825
rect 16419 13791 16477 13825
rect 16511 13791 16569 13825
rect 16603 13791 16661 13825
rect 16695 13791 16753 13825
rect 16787 13791 16845 13825
rect 16879 13791 16937 13825
rect 16971 13791 17029 13825
rect 17063 13791 17121 13825
rect 17155 13791 17213 13825
rect 17247 13791 17305 13825
rect 17339 13791 17397 13825
rect 17431 13791 17489 13825
rect 17523 13791 17581 13825
rect 17615 13791 17673 13825
rect 17707 13791 17765 13825
rect 17799 13791 17857 13825
rect 17891 13791 17949 13825
rect 17983 13791 18041 13825
rect 18075 13791 18133 13825
rect 18167 13791 18225 13825
rect 18259 13791 18317 13825
rect 18351 13791 18409 13825
rect 18443 13791 18501 13825
rect 18535 13791 18593 13825
rect 18627 13791 18685 13825
rect 18719 13791 18777 13825
rect 18811 13791 18869 13825
rect 18903 13791 18961 13825
rect 18995 13791 19053 13825
rect 19087 13791 19145 13825
rect 19179 13791 19237 13825
rect 19271 13791 19329 13825
rect 19363 13791 19421 13825
rect 19455 13791 19513 13825
rect 19547 13791 19605 13825
rect 19639 13791 19697 13825
rect 19731 13791 19789 13825
rect 19823 13791 19881 13825
rect 19915 13791 19973 13825
rect 20007 13791 20065 13825
rect 20099 13791 20157 13825
rect 20191 13791 20220 13825
rect 4965 13749 5207 13791
rect 4965 13715 4983 13749
rect 5017 13715 5155 13749
rect 5189 13715 5207 13749
rect 4965 13654 5207 13715
rect 4965 13620 4983 13654
rect 5017 13620 5155 13654
rect 5189 13620 5207 13654
rect 4965 13573 5207 13620
rect 4965 13505 5015 13539
rect 5049 13505 5069 13539
rect 4965 13431 5069 13505
rect 5103 13499 5207 13573
rect 5103 13465 5123 13499
rect 5157 13465 5207 13499
rect 5425 13749 6127 13791
rect 5425 13715 5443 13749
rect 5477 13715 6075 13749
rect 6109 13715 6127 13749
rect 5425 13647 6127 13715
rect 6162 13749 7231 13791
rect 6162 13715 6179 13749
rect 6213 13715 7179 13749
rect 7213 13715 7231 13749
rect 6162 13704 7231 13715
rect 7265 13720 7323 13791
rect 5425 13613 5443 13647
rect 5477 13613 6075 13647
rect 6109 13613 6127 13647
rect 5425 13573 6127 13613
rect 5425 13503 5763 13573
rect 5425 13469 5503 13503
rect 5537 13469 5606 13503
rect 5640 13469 5709 13503
rect 5743 13469 5763 13503
rect 5797 13505 5817 13539
rect 5851 13505 5916 13539
rect 5950 13505 6015 13539
rect 6049 13505 6127 13539
rect 5797 13435 6127 13505
rect 6480 13503 6550 13704
rect 7265 13686 7277 13720
rect 7311 13686 7323 13720
rect 7450 13749 8519 13791
rect 7450 13715 7467 13749
rect 7501 13715 8467 13749
rect 8501 13715 8519 13749
rect 7450 13704 8519 13715
rect 8554 13749 9623 13791
rect 8554 13715 8571 13749
rect 8605 13715 9571 13749
rect 9605 13715 9623 13749
rect 8554 13704 9623 13715
rect 9675 13741 9709 13757
rect 7265 13627 7323 13686
rect 7265 13593 7277 13627
rect 7311 13593 7323 13627
rect 7265 13558 7323 13593
rect 6480 13469 6499 13503
rect 6533 13469 6550 13503
rect 6480 13454 6550 13469
rect 6846 13539 6914 13556
rect 6846 13505 6863 13539
rect 6897 13505 6914 13539
rect 4965 13378 5207 13431
rect 4965 13344 4983 13378
rect 5017 13344 5155 13378
rect 5189 13344 5207 13378
rect 4965 13281 5207 13344
rect 5425 13376 6127 13435
rect 6846 13390 6914 13505
rect 7768 13503 7838 13704
rect 7768 13469 7787 13503
rect 7821 13469 7838 13503
rect 7768 13454 7838 13469
rect 8134 13539 8202 13556
rect 8134 13505 8151 13539
rect 8185 13505 8202 13539
rect 7265 13409 7323 13426
rect 5425 13342 5443 13376
rect 5477 13342 6075 13376
rect 6109 13342 6127 13376
rect 5425 13281 6127 13342
rect 6162 13376 7231 13390
rect 6162 13342 6179 13376
rect 6213 13342 7179 13376
rect 7213 13342 7231 13376
rect 6162 13281 7231 13342
rect 7265 13375 7277 13409
rect 7311 13375 7323 13409
rect 8134 13390 8202 13505
rect 8872 13503 8942 13704
rect 9675 13673 9709 13707
rect 9745 13741 9811 13791
rect 9745 13707 9761 13741
rect 9795 13707 9811 13741
rect 9745 13673 9811 13707
rect 9745 13639 9761 13673
rect 9795 13639 9811 13673
rect 9845 13741 9899 13757
rect 9845 13707 9847 13741
rect 9881 13707 9899 13741
rect 9845 13660 9899 13707
rect 9675 13605 9709 13639
rect 9845 13626 9847 13660
rect 9881 13626 9899 13660
rect 9951 13725 10005 13791
rect 10131 13790 11386 13791
rect 9951 13691 9968 13725
rect 10002 13691 10005 13725
rect 9951 13642 10005 13691
rect 10039 13705 10097 13756
rect 10039 13671 10054 13705
rect 10088 13671 10097 13705
rect 9675 13571 9808 13605
rect 9845 13576 9899 13626
rect 10039 13619 10097 13671
rect 10131 13725 10182 13790
rect 10131 13691 10140 13725
rect 10174 13691 10182 13725
rect 10131 13645 10182 13691
rect 10219 13705 10271 13756
rect 10219 13671 10226 13705
rect 10260 13671 10271 13705
rect 10039 13608 10054 13619
rect 8872 13469 8891 13503
rect 8925 13469 8942 13503
rect 8872 13454 8942 13469
rect 9238 13539 9306 13556
rect 9238 13505 9255 13539
rect 9289 13505 9306 13539
rect 9774 13542 9808 13571
rect 9238 13390 9306 13505
rect 9661 13519 9727 13535
rect 9661 13485 9669 13519
rect 9703 13513 9727 13519
rect 9661 13479 9677 13485
rect 9711 13479 9727 13513
rect 9661 13461 9727 13479
rect 9774 13526 9831 13542
rect 9774 13492 9797 13526
rect 9774 13476 9831 13492
rect 9774 13425 9808 13476
rect 9675 13391 9808 13425
rect 9865 13416 9899 13576
rect 7265 13281 7323 13375
rect 7450 13376 8519 13390
rect 7450 13342 7467 13376
rect 7501 13342 8467 13376
rect 8501 13342 8519 13376
rect 7450 13281 8519 13342
rect 8554 13376 9623 13390
rect 8554 13342 8571 13376
rect 8605 13342 9571 13376
rect 9605 13342 9623 13376
rect 8554 13281 9623 13342
rect 9675 13370 9709 13391
rect 9847 13387 9899 13416
rect 9951 13585 10054 13608
rect 10088 13608 10097 13619
rect 10219 13619 10271 13671
rect 10305 13725 10354 13790
rect 10305 13691 10312 13725
rect 10346 13691 10354 13725
rect 10305 13645 10354 13691
rect 10391 13723 10443 13756
rect 10391 13705 10405 13723
rect 10391 13671 10398 13705
rect 10439 13689 10443 13723
rect 10432 13671 10443 13689
rect 10219 13608 10226 13619
rect 10088 13585 10226 13608
rect 10260 13611 10271 13619
rect 10391 13619 10443 13671
rect 10477 13725 10526 13790
rect 10477 13691 10484 13725
rect 10518 13691 10526 13725
rect 10477 13645 10526 13691
rect 10563 13705 10615 13756
rect 10563 13671 10570 13705
rect 10604 13671 10615 13705
rect 10391 13611 10398 13619
rect 10260 13585 10398 13611
rect 10432 13611 10443 13619
rect 10563 13619 10615 13671
rect 10649 13725 10698 13790
rect 10649 13691 10655 13725
rect 10689 13691 10698 13725
rect 10649 13645 10698 13691
rect 10732 13705 10784 13756
rect 10732 13671 10741 13705
rect 10775 13671 10784 13705
rect 10563 13611 10570 13619
rect 10432 13585 10570 13611
rect 10604 13611 10615 13619
rect 10732 13619 10784 13671
rect 10818 13725 10870 13790
rect 10818 13691 10827 13725
rect 10861 13691 10870 13725
rect 10818 13645 10870 13691
rect 10904 13705 10956 13756
rect 10904 13671 10913 13705
rect 10947 13671 10956 13705
rect 10732 13611 10741 13619
rect 10604 13585 10741 13611
rect 10775 13611 10784 13619
rect 10904 13619 10956 13671
rect 10990 13725 11042 13790
rect 10990 13691 10999 13725
rect 11033 13691 11042 13725
rect 10990 13645 11042 13691
rect 11076 13705 11128 13756
rect 11076 13671 11085 13705
rect 11119 13671 11128 13705
rect 10904 13611 10913 13619
rect 10775 13585 10913 13611
rect 10947 13611 10956 13619
rect 11076 13619 11128 13671
rect 11162 13725 11214 13790
rect 11162 13691 11171 13725
rect 11205 13691 11214 13725
rect 11162 13645 11214 13691
rect 11248 13705 11300 13756
rect 11248 13671 11257 13705
rect 11291 13671 11300 13705
rect 11076 13611 11085 13619
rect 10947 13585 11085 13611
rect 11119 13611 11128 13619
rect 11248 13619 11300 13671
rect 11334 13749 11386 13790
rect 11334 13715 11343 13749
rect 11377 13715 11386 13749
rect 11334 13681 11386 13715
rect 11334 13647 11343 13681
rect 11377 13647 11386 13681
rect 11334 13631 11386 13647
rect 11420 13733 11470 13756
rect 11420 13699 11429 13733
rect 11463 13699 11470 13733
rect 11420 13665 11470 13699
rect 11420 13631 11429 13665
rect 11463 13631 11470 13665
rect 11248 13611 11257 13619
rect 11119 13585 11257 13611
rect 11291 13585 11300 13619
rect 9951 13563 11300 13585
rect 9951 13445 10184 13563
rect 11420 13529 11470 13631
rect 11506 13749 11558 13791
rect 11506 13715 11515 13749
rect 11549 13715 11558 13749
rect 11506 13681 11558 13715
rect 11506 13647 11515 13681
rect 11549 13647 11558 13681
rect 11506 13629 11558 13647
rect 11593 13741 11642 13757
rect 11593 13707 11601 13741
rect 11635 13707 11642 13741
rect 11593 13673 11642 13707
rect 11593 13639 11601 13673
rect 11635 13639 11642 13673
rect 11593 13529 11642 13639
rect 11678 13749 11737 13791
rect 11678 13715 11687 13749
rect 11721 13715 11737 13749
rect 11678 13681 11737 13715
rect 11678 13647 11687 13681
rect 11721 13647 11737 13681
rect 11678 13629 11737 13647
rect 11865 13749 12383 13791
rect 11865 13715 11883 13749
rect 11917 13715 12331 13749
rect 12365 13715 12383 13749
rect 11865 13647 12383 13715
rect 11865 13613 11883 13647
rect 11917 13613 12331 13647
rect 12365 13613 12383 13647
rect 11865 13573 12383 13613
rect 12417 13720 12475 13791
rect 12417 13686 12429 13720
rect 12463 13686 12475 13720
rect 12417 13627 12475 13686
rect 12417 13593 12429 13627
rect 12463 13593 12475 13627
rect 10218 13513 11642 13529
rect 10218 13479 10238 13513
rect 10272 13479 10306 13513
rect 10340 13479 10374 13513
rect 10408 13479 10442 13513
rect 10476 13479 10510 13513
rect 10544 13479 10578 13513
rect 10612 13479 10646 13513
rect 10680 13479 10714 13513
rect 10748 13479 10782 13513
rect 10816 13479 10850 13513
rect 10884 13479 10918 13513
rect 10952 13479 10986 13513
rect 11020 13479 11054 13513
rect 11088 13479 11122 13513
rect 11156 13479 11190 13513
rect 11224 13479 11258 13513
rect 11292 13479 11642 13513
rect 9951 13411 11300 13445
rect 9881 13383 9899 13387
rect 9675 13315 9709 13336
rect 9745 13323 9761 13357
rect 9795 13323 9811 13357
rect 9745 13281 9811 13323
rect 9847 13349 9853 13353
rect 9887 13349 9899 13383
rect 9847 13315 9899 13349
rect 9951 13361 10011 13377
rect 9951 13327 9968 13361
rect 10002 13327 10011 13361
rect 9951 13281 10011 13327
rect 10045 13370 10097 13411
rect 10045 13336 10054 13370
rect 10088 13336 10097 13370
rect 10045 13320 10097 13336
rect 10131 13361 10183 13377
rect 10131 13327 10140 13361
rect 10174 13327 10183 13361
rect 10131 13281 10183 13327
rect 10219 13370 10271 13411
rect 10219 13336 10226 13370
rect 10260 13336 10271 13370
rect 10219 13320 10271 13336
rect 10305 13361 10355 13377
rect 10305 13327 10312 13361
rect 10346 13327 10355 13361
rect 10305 13281 10355 13327
rect 10391 13370 10443 13411
rect 10391 13336 10398 13370
rect 10432 13336 10443 13370
rect 10391 13320 10443 13336
rect 10477 13361 10527 13377
rect 10477 13327 10484 13361
rect 10518 13327 10527 13361
rect 10477 13281 10527 13327
rect 10563 13370 10615 13411
rect 10563 13336 10570 13370
rect 10604 13336 10615 13370
rect 10563 13320 10615 13336
rect 10649 13361 10698 13377
rect 10649 13327 10655 13361
rect 10689 13327 10698 13361
rect 10649 13281 10698 13327
rect 10732 13370 10787 13411
rect 10732 13336 10741 13370
rect 10775 13336 10787 13370
rect 10732 13320 10787 13336
rect 10821 13361 10870 13377
rect 10821 13327 10827 13361
rect 10861 13327 10870 13361
rect 10821 13281 10870 13327
rect 10904 13370 10956 13411
rect 10904 13336 10913 13370
rect 10947 13336 10956 13370
rect 10904 13320 10956 13336
rect 10990 13361 11042 13377
rect 10990 13327 10999 13361
rect 11033 13327 11042 13361
rect 10990 13281 11042 13327
rect 11076 13370 11128 13411
rect 11076 13336 11085 13370
rect 11119 13336 11128 13370
rect 11076 13320 11128 13336
rect 11162 13361 11214 13377
rect 11162 13327 11171 13361
rect 11205 13327 11214 13361
rect 11162 13281 11214 13327
rect 11248 13370 11300 13411
rect 11248 13336 11257 13370
rect 11291 13336 11300 13370
rect 11248 13320 11300 13336
rect 11334 13370 11386 13393
rect 11334 13336 11343 13370
rect 11377 13336 11386 13370
rect 11334 13281 11386 13336
rect 11420 13370 11470 13479
rect 11420 13336 11429 13370
rect 11463 13336 11470 13370
rect 11420 13317 11470 13336
rect 11506 13370 11558 13386
rect 11506 13336 11515 13370
rect 11549 13336 11558 13370
rect 11506 13281 11558 13336
rect 11592 13370 11642 13479
rect 11676 13519 11739 13529
rect 11676 13513 11693 13519
rect 11676 13479 11685 13513
rect 11727 13485 11739 13519
rect 11719 13479 11739 13485
rect 11676 13417 11739 13479
rect 11865 13503 12107 13573
rect 12417 13558 12475 13593
rect 12509 13741 12563 13757
rect 12509 13707 12527 13741
rect 12561 13707 12563 13741
rect 12509 13660 12563 13707
rect 12509 13626 12527 13660
rect 12561 13626 12563 13660
rect 12597 13741 12663 13791
rect 12597 13707 12613 13741
rect 12647 13707 12663 13741
rect 12597 13673 12663 13707
rect 12597 13639 12613 13673
rect 12647 13639 12663 13673
rect 12699 13741 12733 13757
rect 12963 13749 13024 13791
rect 12699 13673 12733 13707
rect 12509 13576 12563 13626
rect 12699 13605 12733 13639
rect 11865 13469 11943 13503
rect 11977 13469 12053 13503
rect 12087 13469 12107 13503
rect 12141 13505 12161 13539
rect 12195 13505 12271 13539
rect 12305 13505 12383 13539
rect 12141 13435 12383 13505
rect 11592 13336 11601 13370
rect 11635 13336 11642 13370
rect 11592 13317 11642 13336
rect 11678 13357 11739 13383
rect 11678 13323 11687 13357
rect 11721 13323 11739 13357
rect 11678 13281 11739 13323
rect 11865 13376 12383 13435
rect 11865 13342 11883 13376
rect 11917 13342 12331 13376
rect 12365 13342 12383 13376
rect 11865 13281 12383 13342
rect 12417 13409 12475 13426
rect 12417 13375 12429 13409
rect 12463 13375 12475 13409
rect 12417 13281 12475 13375
rect 12509 13416 12543 13576
rect 12600 13571 12733 13605
rect 12878 13723 12929 13729
rect 12878 13689 12889 13723
rect 12923 13713 12929 13723
rect 12878 13679 12895 13689
rect 12878 13645 12929 13679
rect 12878 13611 12895 13645
rect 12600 13542 12634 13571
rect 12577 13526 12634 13542
rect 12878 13553 12929 13611
rect 12963 13715 12979 13749
rect 13013 13715 13024 13749
rect 13092 13749 13158 13791
rect 13092 13715 13108 13749
rect 13142 13715 13158 13749
rect 13262 13749 13312 13791
rect 13194 13723 13228 13739
rect 12963 13681 13024 13715
rect 13262 13715 13278 13749
rect 13262 13699 13312 13715
rect 13346 13748 13520 13757
rect 13346 13714 13470 13748
rect 13504 13714 13520 13748
rect 13194 13681 13228 13689
rect 12963 13647 12979 13681
rect 13013 13647 13024 13681
rect 12963 13563 13024 13647
rect 13068 13647 13228 13681
rect 13346 13689 13520 13714
rect 13567 13741 13601 13757
rect 12611 13492 12634 13526
rect 12577 13476 12634 13492
rect 12600 13425 12634 13476
rect 12681 13519 12747 13535
rect 12681 13513 12705 13519
rect 12681 13479 12697 13513
rect 12739 13485 12747 13519
rect 12731 13479 12747 13485
rect 12681 13461 12747 13479
rect 12509 13387 12561 13416
rect 12600 13391 12733 13425
rect 12509 13383 12527 13387
rect 12509 13349 12521 13383
rect 12699 13370 12733 13391
rect 12555 13349 12561 13353
rect 12509 13315 12561 13349
rect 12597 13323 12613 13357
rect 12647 13323 12663 13357
rect 12597 13281 12663 13323
rect 12699 13315 12733 13336
rect 12878 13423 12920 13553
rect 13068 13529 13102 13647
rect 13346 13613 13380 13689
rect 13567 13665 13601 13707
rect 13635 13749 13709 13791
rect 13635 13715 13655 13749
rect 13689 13715 13709 13749
rect 13836 13739 13902 13791
rect 14017 13747 14153 13757
rect 13635 13699 13709 13715
rect 13768 13723 13802 13739
rect 13836 13705 13852 13739
rect 13886 13705 13902 13739
rect 13949 13723 13983 13739
rect 13768 13671 13802 13689
rect 13949 13671 13983 13689
rect 13136 13579 13152 13613
rect 13186 13579 13380 13613
rect 13414 13629 13461 13655
rect 13414 13595 13430 13629
rect 13495 13621 13506 13655
rect 13567 13631 13679 13665
rect 13768 13637 13983 13671
rect 14017 13713 14103 13747
rect 14137 13713 14153 13747
rect 14017 13691 14153 13713
rect 14196 13741 14246 13757
rect 14230 13707 14246 13741
rect 14196 13691 14246 13707
rect 14280 13749 14330 13791
rect 14314 13715 14330 13749
rect 14280 13699 14330 13715
rect 13464 13597 13506 13621
rect 13645 13603 13679 13631
rect 13464 13595 13607 13597
rect 13346 13561 13380 13579
rect 13472 13563 13607 13595
rect 12954 13523 13102 13529
rect 12954 13513 13137 13523
rect 12988 13479 13137 13513
rect 12954 13463 13137 13479
rect 13072 13428 13137 13463
rect 12878 13407 12929 13423
rect 12878 13373 12895 13407
rect 13073 13373 13137 13428
rect 13171 13514 13279 13545
rect 13346 13527 13427 13561
rect 13171 13505 13245 13514
rect 13171 13471 13229 13505
rect 13263 13471 13279 13480
rect 13315 13477 13359 13493
rect 13171 13451 13219 13471
rect 13171 13417 13185 13451
rect 13315 13443 13325 13477
rect 13315 13437 13359 13443
rect 13171 13391 13219 13417
rect 13253 13403 13359 13437
rect 12878 13317 12929 13373
rect 12963 13357 13024 13373
rect 12963 13323 12979 13357
rect 13013 13323 13024 13357
rect 13073 13339 13103 13373
rect 13253 13357 13287 13403
rect 13393 13371 13427 13527
rect 13461 13519 13531 13529
rect 13495 13503 13531 13519
rect 13461 13469 13469 13485
rect 13503 13469 13531 13503
rect 13461 13405 13531 13469
rect 13565 13455 13607 13563
rect 13599 13421 13607 13455
rect 13565 13405 13607 13421
rect 13645 13569 13895 13603
rect 13929 13569 13945 13603
rect 13645 13431 13679 13569
rect 14017 13535 14051 13691
rect 14212 13665 14246 13691
rect 13713 13515 14051 13535
rect 13747 13501 14051 13515
rect 14085 13655 14178 13657
rect 14119 13629 14178 13655
rect 14212 13631 14291 13665
rect 14119 13621 14144 13629
rect 14085 13595 14144 13621
rect 14085 13579 14178 13595
rect 13713 13465 13747 13481
rect 13781 13433 13809 13467
rect 13843 13451 13939 13467
rect 13137 13339 13287 13357
rect 13073 13323 13287 13339
rect 13321 13353 13359 13369
rect 12963 13281 13024 13323
rect 13355 13319 13359 13353
rect 13321 13281 13359 13319
rect 13393 13357 13583 13371
rect 13393 13323 13533 13357
rect 13567 13323 13583 13357
rect 13645 13353 13697 13431
rect 13781 13417 13833 13433
rect 13867 13417 13905 13451
rect 13393 13315 13583 13323
rect 13627 13319 13643 13353
rect 13677 13319 13697 13353
rect 13739 13357 13805 13373
rect 13739 13323 13755 13357
rect 13789 13323 13805 13357
rect 13980 13359 14014 13501
rect 14085 13461 14119 13579
rect 14048 13427 14064 13461
rect 14098 13427 14119 13461
rect 14048 13417 14119 13427
rect 14153 13519 14223 13541
rect 14153 13485 14177 13519
rect 14211 13485 14223 13519
rect 14153 13467 14223 13485
rect 14153 13433 14166 13467
rect 14200 13433 14223 13467
rect 14153 13417 14223 13433
rect 14257 13359 14291 13631
rect 14364 13597 14429 13754
rect 14463 13741 14497 13757
rect 14463 13673 14497 13707
rect 14531 13725 14597 13791
rect 14531 13691 14547 13725
rect 14581 13691 14597 13725
rect 14631 13741 14682 13757
rect 14665 13707 14682 13741
rect 14631 13673 14682 13707
rect 14325 13574 14417 13597
rect 14359 13540 14417 13574
rect 14325 13451 14417 13540
rect 14325 13417 14361 13451
rect 14395 13417 14417 13451
rect 14325 13387 14417 13417
rect 13980 13325 14101 13359
rect 14135 13325 14151 13359
rect 14192 13325 14208 13359
rect 14242 13325 14291 13359
rect 14463 13383 14497 13621
rect 14532 13639 14631 13657
rect 14665 13639 14682 13673
rect 14532 13623 14682 13639
rect 14719 13749 14778 13791
rect 14719 13715 14735 13749
rect 14769 13715 14778 13749
rect 14719 13681 14778 13715
rect 14719 13647 14735 13681
rect 14769 13647 14778 13681
rect 14719 13629 14778 13647
rect 14814 13741 14863 13757
rect 14814 13707 14821 13741
rect 14855 13707 14863 13741
rect 14814 13673 14863 13707
rect 14814 13639 14821 13673
rect 14855 13639 14863 13673
rect 14532 13528 14578 13623
rect 14566 13519 14578 13528
rect 14532 13485 14544 13494
rect 14532 13425 14578 13485
rect 14612 13587 14682 13589
rect 14612 13553 14637 13587
rect 14671 13553 14682 13587
rect 14612 13513 14682 13553
rect 14814 13529 14863 13639
rect 14898 13749 14950 13791
rect 15070 13790 16325 13791
rect 14898 13715 14907 13749
rect 14941 13715 14950 13749
rect 14898 13681 14950 13715
rect 14898 13647 14907 13681
rect 14941 13647 14950 13681
rect 14898 13629 14950 13647
rect 14986 13733 15036 13756
rect 14986 13699 14993 13733
rect 15027 13699 15036 13733
rect 14986 13665 15036 13699
rect 14986 13631 14993 13665
rect 15027 13631 15036 13665
rect 15070 13749 15122 13790
rect 15070 13715 15079 13749
rect 15113 13715 15122 13749
rect 15070 13681 15122 13715
rect 15070 13647 15079 13681
rect 15113 13647 15122 13681
rect 15070 13631 15122 13647
rect 15156 13705 15208 13756
rect 15156 13671 15165 13705
rect 15199 13671 15208 13705
rect 14986 13529 15036 13631
rect 15156 13619 15208 13671
rect 15242 13725 15294 13790
rect 15242 13691 15251 13725
rect 15285 13691 15294 13725
rect 15242 13645 15294 13691
rect 15328 13705 15380 13756
rect 15328 13671 15337 13705
rect 15371 13671 15380 13705
rect 15156 13585 15165 13619
rect 15199 13611 15208 13619
rect 15328 13619 15380 13671
rect 15414 13725 15466 13790
rect 15414 13691 15423 13725
rect 15457 13691 15466 13725
rect 15414 13645 15466 13691
rect 15500 13705 15552 13756
rect 15500 13671 15509 13705
rect 15543 13671 15552 13705
rect 15328 13611 15337 13619
rect 15199 13585 15337 13611
rect 15371 13611 15380 13619
rect 15500 13619 15552 13671
rect 15586 13725 15638 13790
rect 15586 13691 15595 13725
rect 15629 13691 15638 13725
rect 15586 13645 15638 13691
rect 15672 13705 15724 13756
rect 15672 13671 15681 13705
rect 15715 13671 15724 13705
rect 15500 13611 15509 13619
rect 15371 13585 15509 13611
rect 15543 13611 15552 13619
rect 15672 13619 15724 13671
rect 15758 13725 15807 13790
rect 15758 13691 15767 13725
rect 15801 13691 15807 13725
rect 15758 13645 15807 13691
rect 15841 13705 15893 13756
rect 15841 13671 15852 13705
rect 15886 13671 15893 13705
rect 15672 13611 15681 13619
rect 15543 13585 15681 13611
rect 15715 13611 15724 13619
rect 15841 13619 15893 13671
rect 15930 13725 15979 13790
rect 15930 13691 15938 13725
rect 15972 13691 15979 13725
rect 15930 13645 15979 13691
rect 16013 13705 16065 13756
rect 16013 13671 16024 13705
rect 16058 13671 16065 13705
rect 15841 13611 15852 13619
rect 15715 13585 15852 13611
rect 15886 13611 15893 13619
rect 16013 13619 16065 13671
rect 16102 13725 16151 13790
rect 16102 13691 16110 13725
rect 16144 13691 16151 13725
rect 16102 13645 16151 13691
rect 16185 13723 16237 13756
rect 16185 13705 16201 13723
rect 16185 13671 16196 13705
rect 16235 13689 16237 13723
rect 16230 13671 16237 13689
rect 16013 13611 16024 13619
rect 15886 13585 16024 13611
rect 16058 13611 16065 13619
rect 16185 13619 16237 13671
rect 16274 13725 16325 13790
rect 16274 13691 16282 13725
rect 16316 13691 16325 13725
rect 16274 13645 16325 13691
rect 16359 13705 16417 13756
rect 16359 13671 16368 13705
rect 16402 13671 16417 13705
rect 16185 13611 16196 13619
rect 16058 13585 16196 13611
rect 16230 13608 16237 13619
rect 16359 13619 16417 13671
rect 16451 13725 16505 13791
rect 16451 13691 16454 13725
rect 16488 13691 16505 13725
rect 16451 13642 16505 13691
rect 16558 13749 16625 13757
rect 16558 13723 16575 13749
rect 16558 13689 16569 13723
rect 16609 13715 16625 13749
rect 16603 13689 16625 13715
rect 16558 13681 16625 13689
rect 16558 13647 16575 13681
rect 16609 13647 16625 13681
rect 16359 13608 16368 13619
rect 16230 13585 16368 13608
rect 16402 13608 16417 13619
rect 16558 13613 16625 13647
rect 16402 13585 16505 13608
rect 15156 13563 16505 13585
rect 14612 13479 14634 13513
rect 14668 13479 14682 13513
rect 14612 13459 14682 13479
rect 14717 13519 14780 13529
rect 14717 13485 14729 13519
rect 14763 13513 14780 13519
rect 14717 13479 14737 13485
rect 14771 13479 14780 13513
rect 14532 13391 14682 13425
rect 14717 13417 14780 13479
rect 14814 13513 16238 13529
rect 14814 13479 15164 13513
rect 15198 13479 15232 13513
rect 15266 13479 15300 13513
rect 15334 13479 15368 13513
rect 15402 13479 15436 13513
rect 15470 13479 15504 13513
rect 15538 13479 15572 13513
rect 15606 13479 15640 13513
rect 15674 13479 15708 13513
rect 15742 13479 15776 13513
rect 15810 13479 15844 13513
rect 15878 13479 15912 13513
rect 15946 13479 15980 13513
rect 16014 13479 16048 13513
rect 16082 13479 16116 13513
rect 16150 13479 16184 13513
rect 16218 13479 16238 13513
rect 13739 13281 13805 13323
rect 14325 13319 14341 13353
rect 14375 13319 14391 13353
rect 14631 13383 14682 13391
rect 14463 13333 14497 13349
rect 14325 13281 14391 13319
rect 14531 13323 14547 13357
rect 14581 13323 14597 13357
rect 14665 13349 14682 13383
rect 14631 13333 14682 13349
rect 14717 13357 14778 13383
rect 14531 13281 14597 13323
rect 14717 13323 14735 13357
rect 14769 13323 14778 13357
rect 14717 13281 14778 13323
rect 14814 13370 14864 13479
rect 14814 13336 14821 13370
rect 14855 13336 14864 13370
rect 14814 13317 14864 13336
rect 14898 13370 14950 13386
rect 14898 13336 14907 13370
rect 14941 13336 14950 13370
rect 14898 13281 14950 13336
rect 14986 13370 15036 13479
rect 16272 13445 16505 13563
rect 15156 13411 16505 13445
rect 16558 13579 16575 13613
rect 16609 13579 16625 13613
rect 16558 13563 16625 13579
rect 16659 13749 16693 13791
rect 16659 13681 16693 13715
rect 16659 13613 16693 13647
rect 16659 13563 16693 13579
rect 16727 13723 17133 13757
rect 16558 13429 16592 13563
rect 16727 13529 16761 13723
rect 16626 13513 16677 13529
rect 16660 13479 16677 13513
rect 16626 13463 16677 13479
rect 16722 13513 16761 13529
rect 16756 13479 16761 13513
rect 16722 13463 16761 13479
rect 16795 13655 16895 13689
rect 16929 13655 16970 13689
rect 17004 13655 17020 13689
rect 16643 13429 16677 13463
rect 16795 13429 16829 13655
rect 14986 13336 14993 13370
rect 15027 13336 15036 13370
rect 14986 13317 15036 13336
rect 15070 13370 15122 13393
rect 15070 13336 15079 13370
rect 15113 13336 15122 13370
rect 15070 13281 15122 13336
rect 15156 13370 15208 13411
rect 15156 13336 15165 13370
rect 15199 13336 15208 13370
rect 15156 13320 15208 13336
rect 15242 13361 15294 13377
rect 15242 13327 15251 13361
rect 15285 13327 15294 13361
rect 15242 13281 15294 13327
rect 15328 13370 15380 13411
rect 15328 13336 15337 13370
rect 15371 13336 15380 13370
rect 15328 13320 15380 13336
rect 15414 13361 15466 13377
rect 15414 13327 15423 13361
rect 15457 13327 15466 13361
rect 15414 13281 15466 13327
rect 15500 13370 15552 13411
rect 15500 13336 15509 13370
rect 15543 13336 15552 13370
rect 15500 13320 15552 13336
rect 15586 13361 15635 13377
rect 15586 13327 15595 13361
rect 15629 13327 15635 13361
rect 15586 13281 15635 13327
rect 15669 13370 15724 13411
rect 15669 13336 15681 13370
rect 15715 13336 15724 13370
rect 15669 13320 15724 13336
rect 15758 13361 15807 13377
rect 15758 13327 15767 13361
rect 15801 13327 15807 13361
rect 15758 13281 15807 13327
rect 15841 13370 15893 13411
rect 15841 13336 15852 13370
rect 15886 13336 15893 13370
rect 15841 13320 15893 13336
rect 15929 13361 15979 13377
rect 15929 13327 15938 13361
rect 15972 13327 15979 13361
rect 15929 13281 15979 13327
rect 16013 13370 16065 13411
rect 16013 13336 16024 13370
rect 16058 13336 16065 13370
rect 16013 13320 16065 13336
rect 16101 13361 16151 13377
rect 16101 13327 16110 13361
rect 16144 13327 16151 13361
rect 16101 13281 16151 13327
rect 16185 13370 16237 13411
rect 16185 13336 16196 13370
rect 16230 13336 16237 13370
rect 16185 13320 16237 13336
rect 16273 13361 16325 13377
rect 16273 13327 16282 13361
rect 16316 13327 16325 13361
rect 16273 13281 16325 13327
rect 16359 13370 16411 13411
rect 16359 13336 16368 13370
rect 16402 13336 16411 13370
rect 16359 13320 16411 13336
rect 16445 13361 16505 13377
rect 16445 13327 16454 13361
rect 16488 13327 16505 13361
rect 16445 13281 16505 13327
rect 16558 13376 16609 13429
rect 16643 13395 16829 13429
rect 16863 13590 17065 13621
rect 16863 13587 17031 13590
rect 16863 13477 16897 13587
rect 17027 13556 17031 13587
rect 16938 13519 16993 13547
rect 16971 13485 16993 13519
rect 16863 13427 16897 13443
rect 16938 13477 16993 13485
rect 16938 13443 16959 13477
rect 16558 13342 16575 13376
rect 16794 13388 16829 13395
rect 16794 13372 16900 13388
rect 16558 13315 16609 13342
rect 16643 13357 16709 13361
rect 16643 13323 16659 13357
rect 16693 13323 16709 13357
rect 16643 13281 16709 13323
rect 16794 13338 16866 13372
rect 16794 13315 16900 13338
rect 16938 13315 16993 13443
rect 17027 13383 17065 13556
rect 17099 13590 17133 13723
rect 17167 13689 17201 13791
rect 17167 13639 17201 13655
rect 17248 13689 17351 13721
rect 17248 13655 17253 13689
rect 17287 13655 17351 13689
rect 17248 13639 17351 13655
rect 17099 13587 17199 13590
rect 17099 13553 17121 13587
rect 17155 13556 17199 13587
rect 17233 13556 17249 13590
rect 17155 13553 17249 13556
rect 17099 13552 17249 13553
rect 17283 13477 17351 13639
rect 17569 13720 17627 13791
rect 17569 13686 17581 13720
rect 17615 13686 17627 13720
rect 17754 13749 18823 13791
rect 17754 13715 17771 13749
rect 17805 13715 18771 13749
rect 18805 13715 18823 13749
rect 17754 13704 18823 13715
rect 18858 13749 19927 13791
rect 18858 13715 18875 13749
rect 18909 13715 19875 13749
rect 19909 13715 19927 13749
rect 18858 13704 19927 13715
rect 19961 13749 20203 13791
rect 19961 13715 19979 13749
rect 20013 13715 20151 13749
rect 20185 13715 20203 13749
rect 17569 13627 17627 13686
rect 17569 13593 17581 13627
rect 17615 13593 17627 13627
rect 17569 13558 17627 13593
rect 17105 13443 17121 13477
rect 17155 13443 17351 13477
rect 18072 13503 18142 13704
rect 18072 13469 18091 13503
rect 18125 13469 18142 13503
rect 18072 13454 18142 13469
rect 18438 13539 18506 13556
rect 18438 13505 18455 13539
rect 18489 13505 18506 13539
rect 17027 13349 17029 13383
rect 17063 13349 17065 13383
rect 17027 13315 17065 13349
rect 17101 13372 17203 13388
rect 17135 13338 17169 13372
rect 17101 13281 17203 13338
rect 17247 13372 17296 13443
rect 17247 13338 17253 13372
rect 17287 13338 17296 13372
rect 17247 13322 17296 13338
rect 17569 13409 17627 13426
rect 17569 13375 17581 13409
rect 17615 13375 17627 13409
rect 18438 13390 18506 13505
rect 19176 13503 19246 13704
rect 19961 13654 20203 13715
rect 19961 13620 19979 13654
rect 20013 13620 20151 13654
rect 20185 13620 20203 13654
rect 19961 13573 20203 13620
rect 19176 13469 19195 13503
rect 19229 13469 19246 13503
rect 19176 13454 19246 13469
rect 19542 13539 19610 13556
rect 19542 13505 19559 13539
rect 19593 13505 19610 13539
rect 19542 13390 19610 13505
rect 19961 13499 20065 13573
rect 19961 13465 20011 13499
rect 20045 13465 20065 13499
rect 20099 13505 20119 13539
rect 20153 13505 20203 13539
rect 20099 13431 20203 13505
rect 17569 13281 17627 13375
rect 17754 13376 18823 13390
rect 17754 13342 17771 13376
rect 17805 13342 18771 13376
rect 18805 13342 18823 13376
rect 17754 13281 18823 13342
rect 18858 13376 19927 13390
rect 18858 13342 18875 13376
rect 18909 13342 19875 13376
rect 19909 13342 19927 13376
rect 18858 13281 19927 13342
rect 19961 13378 20203 13431
rect 19961 13344 19979 13378
rect 20013 13344 20151 13378
rect 20185 13344 20203 13378
rect 19961 13281 20203 13344
rect 4948 13247 4977 13281
rect 5011 13247 5069 13281
rect 5103 13247 5161 13281
rect 5195 13247 5253 13281
rect 5287 13247 5345 13281
rect 5379 13247 5437 13281
rect 5471 13247 5529 13281
rect 5563 13247 5621 13281
rect 5655 13247 5713 13281
rect 5747 13247 5805 13281
rect 5839 13247 5897 13281
rect 5931 13247 5989 13281
rect 6023 13247 6081 13281
rect 6115 13247 6173 13281
rect 6207 13247 6265 13281
rect 6299 13247 6357 13281
rect 6391 13247 6449 13281
rect 6483 13247 6541 13281
rect 6575 13247 6633 13281
rect 6667 13247 6725 13281
rect 6759 13247 6817 13281
rect 6851 13247 6909 13281
rect 6943 13247 7001 13281
rect 7035 13247 7093 13281
rect 7127 13247 7185 13281
rect 7219 13247 7277 13281
rect 7311 13247 7369 13281
rect 7403 13247 7461 13281
rect 7495 13247 7553 13281
rect 7587 13247 7645 13281
rect 7679 13247 7737 13281
rect 7771 13247 7829 13281
rect 7863 13247 7921 13281
rect 7955 13247 8013 13281
rect 8047 13247 8105 13281
rect 8139 13247 8197 13281
rect 8231 13247 8289 13281
rect 8323 13247 8381 13281
rect 8415 13247 8473 13281
rect 8507 13247 8565 13281
rect 8599 13247 8657 13281
rect 8691 13247 8749 13281
rect 8783 13247 8841 13281
rect 8875 13247 8933 13281
rect 8967 13247 9025 13281
rect 9059 13247 9117 13281
rect 9151 13247 9209 13281
rect 9243 13247 9301 13281
rect 9335 13247 9393 13281
rect 9427 13247 9485 13281
rect 9519 13247 9577 13281
rect 9611 13247 9669 13281
rect 9703 13247 9761 13281
rect 9795 13247 9853 13281
rect 9887 13247 9945 13281
rect 9979 13247 10037 13281
rect 10071 13247 10129 13281
rect 10163 13247 10221 13281
rect 10255 13247 10313 13281
rect 10347 13247 10405 13281
rect 10439 13247 10497 13281
rect 10531 13247 10589 13281
rect 10623 13247 10681 13281
rect 10715 13247 10773 13281
rect 10807 13247 10865 13281
rect 10899 13247 10957 13281
rect 10991 13247 11049 13281
rect 11083 13247 11141 13281
rect 11175 13247 11233 13281
rect 11267 13247 11325 13281
rect 11359 13247 11417 13281
rect 11451 13247 11509 13281
rect 11543 13247 11601 13281
rect 11635 13247 11693 13281
rect 11727 13247 11785 13281
rect 11819 13247 11877 13281
rect 11911 13247 11969 13281
rect 12003 13247 12061 13281
rect 12095 13247 12153 13281
rect 12187 13247 12245 13281
rect 12279 13247 12337 13281
rect 12371 13247 12429 13281
rect 12463 13247 12521 13281
rect 12555 13247 12613 13281
rect 12647 13247 12705 13281
rect 12739 13247 12797 13281
rect 12831 13247 12889 13281
rect 12923 13247 12981 13281
rect 13015 13247 13073 13281
rect 13107 13247 13165 13281
rect 13199 13247 13257 13281
rect 13291 13247 13349 13281
rect 13383 13247 13441 13281
rect 13475 13247 13533 13281
rect 13567 13247 13625 13281
rect 13659 13247 13717 13281
rect 13751 13247 13809 13281
rect 13843 13247 13901 13281
rect 13935 13247 13993 13281
rect 14027 13247 14085 13281
rect 14119 13247 14177 13281
rect 14211 13247 14269 13281
rect 14303 13247 14361 13281
rect 14395 13247 14453 13281
rect 14487 13247 14545 13281
rect 14579 13247 14637 13281
rect 14671 13247 14729 13281
rect 14763 13247 14821 13281
rect 14855 13247 14913 13281
rect 14947 13247 15005 13281
rect 15039 13247 15097 13281
rect 15131 13247 15189 13281
rect 15223 13247 15281 13281
rect 15315 13247 15373 13281
rect 15407 13247 15465 13281
rect 15499 13247 15557 13281
rect 15591 13247 15649 13281
rect 15683 13247 15741 13281
rect 15775 13247 15833 13281
rect 15867 13247 15925 13281
rect 15959 13247 16017 13281
rect 16051 13247 16109 13281
rect 16143 13247 16201 13281
rect 16235 13247 16293 13281
rect 16327 13247 16385 13281
rect 16419 13247 16477 13281
rect 16511 13247 16569 13281
rect 16603 13247 16661 13281
rect 16695 13247 16753 13281
rect 16787 13247 16845 13281
rect 16879 13247 16937 13281
rect 16971 13247 17029 13281
rect 17063 13247 17121 13281
rect 17155 13247 17213 13281
rect 17247 13247 17305 13281
rect 17339 13247 17397 13281
rect 17431 13247 17489 13281
rect 17523 13247 17581 13281
rect 17615 13247 17673 13281
rect 17707 13247 17765 13281
rect 17799 13247 17857 13281
rect 17891 13247 17949 13281
rect 17983 13247 18041 13281
rect 18075 13247 18133 13281
rect 18167 13247 18225 13281
rect 18259 13247 18317 13281
rect 18351 13247 18409 13281
rect 18443 13247 18501 13281
rect 18535 13247 18593 13281
rect 18627 13247 18685 13281
rect 18719 13247 18777 13281
rect 18811 13247 18869 13281
rect 18903 13247 18961 13281
rect 18995 13247 19053 13281
rect 19087 13247 19145 13281
rect 19179 13247 19237 13281
rect 19271 13247 19329 13281
rect 19363 13247 19421 13281
rect 19455 13247 19513 13281
rect 19547 13247 19605 13281
rect 19639 13247 19697 13281
rect 19731 13247 19789 13281
rect 19823 13247 19881 13281
rect 19915 13247 19973 13281
rect 20007 13247 20065 13281
rect 20099 13247 20157 13281
rect 20191 13247 20220 13281
rect 4965 13184 5207 13247
rect 4965 13150 4983 13184
rect 5017 13150 5155 13184
rect 5189 13150 5207 13184
rect 4965 13097 5207 13150
rect 5241 13186 5759 13247
rect 5241 13152 5259 13186
rect 5293 13152 5707 13186
rect 5741 13152 5759 13186
rect 4965 13023 5069 13097
rect 5241 13093 5759 13152
rect 5794 13186 6863 13247
rect 5794 13152 5811 13186
rect 5845 13152 6811 13186
rect 6845 13152 6863 13186
rect 5794 13138 6863 13152
rect 6898 13186 7967 13247
rect 6898 13152 6915 13186
rect 6949 13152 7915 13186
rect 7949 13152 7967 13186
rect 6898 13138 7967 13152
rect 8002 13186 9071 13247
rect 8002 13152 8019 13186
rect 8053 13152 9019 13186
rect 9053 13152 9071 13186
rect 8002 13138 9071 13152
rect 9128 13179 9185 13213
rect 9128 13145 9145 13179
rect 9179 13145 9185 13179
rect 9219 13205 9273 13247
rect 9219 13171 9229 13205
rect 9263 13171 9273 13205
rect 9219 13155 9273 13171
rect 9353 13179 9433 13213
rect 4965 12989 5015 13023
rect 5049 12989 5069 13023
rect 5103 13029 5123 13063
rect 5157 13029 5207 13063
rect 5103 12955 5207 13029
rect 4965 12908 5207 12955
rect 4965 12874 4983 12908
rect 5017 12874 5155 12908
rect 5189 12874 5207 12908
rect 4965 12813 5207 12874
rect 4965 12779 4983 12813
rect 5017 12779 5155 12813
rect 5189 12779 5207 12813
rect 4965 12737 5207 12779
rect 5241 13025 5319 13059
rect 5353 13025 5429 13059
rect 5463 13025 5483 13059
rect 5241 12955 5483 13025
rect 5517 13023 5759 13093
rect 5517 12989 5537 13023
rect 5571 12989 5647 13023
rect 5681 12989 5759 13023
rect 6112 13059 6182 13074
rect 6112 13025 6131 13059
rect 6165 13025 6182 13059
rect 5241 12915 5759 12955
rect 5241 12881 5259 12915
rect 5293 12881 5707 12915
rect 5741 12881 5759 12915
rect 5241 12813 5759 12881
rect 6112 12824 6182 13025
rect 6478 13023 6546 13138
rect 6478 12989 6495 13023
rect 6529 12989 6546 13023
rect 6478 12972 6546 12989
rect 7216 13059 7286 13074
rect 7216 13025 7235 13059
rect 7269 13025 7286 13059
rect 7216 12824 7286 13025
rect 7582 13023 7650 13138
rect 7582 12989 7599 13023
rect 7633 12989 7650 13023
rect 7582 12972 7650 12989
rect 8320 13059 8390 13074
rect 8320 13025 8339 13059
rect 8373 13025 8390 13059
rect 8320 12824 8390 13025
rect 8686 13023 8754 13138
rect 9128 13121 9185 13145
rect 9353 13145 9383 13179
rect 9417 13145 9433 13179
rect 9128 13087 9319 13121
rect 8686 12989 8703 13023
rect 8737 12989 8754 13023
rect 8686 12972 8754 12989
rect 9105 13049 9243 13053
rect 9105 13015 9169 13049
rect 9203 13015 9243 13049
rect 9105 12975 9243 13015
rect 9105 12941 9209 12975
rect 9277 13049 9319 13087
rect 9277 13015 9283 13049
rect 9317 13015 9319 13049
rect 9277 12907 9319 13015
rect 9128 12863 9319 12907
rect 9353 13053 9433 13145
rect 9471 13179 9527 13213
rect 9471 13145 9487 13179
rect 9521 13145 9527 13179
rect 9631 13205 9696 13247
rect 9631 13171 9646 13205
rect 9680 13171 9696 13205
rect 9631 13155 9696 13171
rect 9730 13179 9807 13213
rect 9471 13121 9527 13145
rect 9730 13145 9736 13179
rect 9770 13145 9807 13179
rect 9471 13087 9696 13121
rect 9730 13099 9807 13145
rect 9841 13153 9899 13247
rect 9841 13119 9853 13153
rect 9887 13119 9899 13153
rect 9841 13102 9899 13119
rect 10025 13179 10359 13247
rect 10025 13145 10043 13179
rect 10077 13145 10307 13179
rect 10341 13145 10359 13179
rect 9606 13065 9696 13087
rect 9353 13049 9572 13053
rect 9353 13015 9487 13049
rect 9521 13015 9572 13049
rect 9353 12941 9572 13015
rect 9606 13049 9717 13065
rect 9606 13015 9683 13049
rect 9606 12999 9717 13015
rect 9128 12839 9185 12863
rect 5241 12779 5259 12813
rect 5293 12779 5707 12813
rect 5741 12779 5759 12813
rect 5241 12737 5759 12779
rect 5794 12813 6863 12824
rect 5794 12779 5811 12813
rect 5845 12779 6811 12813
rect 6845 12779 6863 12813
rect 5794 12737 6863 12779
rect 6898 12813 7967 12824
rect 6898 12779 6915 12813
rect 6949 12779 7915 12813
rect 7949 12779 7967 12813
rect 6898 12737 7967 12779
rect 8002 12813 9071 12824
rect 8002 12779 8019 12813
rect 8053 12779 9019 12813
rect 9053 12779 9071 12813
rect 8002 12737 9071 12779
rect 9128 12805 9145 12839
rect 9179 12805 9185 12839
rect 9353 12839 9433 12941
rect 9606 12907 9696 12999
rect 9751 12965 9807 13099
rect 10025 13093 10359 13145
rect 10025 13025 10045 13059
rect 10079 13025 10175 13059
rect 9128 12771 9185 12805
rect 9219 12813 9273 12829
rect 9219 12779 9229 12813
rect 9263 12779 9273 12813
rect 9219 12737 9273 12779
rect 9353 12805 9383 12839
rect 9417 12805 9433 12839
rect 9353 12771 9433 12805
rect 9471 12863 9696 12907
rect 9471 12839 9527 12863
rect 9471 12805 9487 12839
rect 9521 12805 9527 12839
rect 9730 12839 9807 12965
rect 9471 12771 9527 12805
rect 9631 12813 9696 12829
rect 9631 12779 9646 12813
rect 9680 12779 9696 12813
rect 9631 12737 9696 12779
rect 9730 12805 9736 12839
rect 9795 12805 9807 12839
rect 9730 12771 9807 12805
rect 9841 12935 9899 12970
rect 9841 12901 9853 12935
rect 9887 12901 9899 12935
rect 9841 12842 9899 12901
rect 9841 12808 9853 12842
rect 9887 12808 9899 12842
rect 9841 12737 9899 12808
rect 10025 12955 10175 13025
rect 10209 13023 10359 13093
rect 10209 12989 10305 13023
rect 10339 12989 10359 13023
rect 10394 13155 10445 13211
rect 10479 13205 10540 13247
rect 10837 13209 10875 13247
rect 10479 13171 10495 13205
rect 10529 13171 10540 13205
rect 10479 13155 10540 13171
rect 10589 13189 10803 13205
rect 10589 13155 10619 13189
rect 10653 13171 10803 13189
rect 10394 13121 10411 13155
rect 10394 13105 10445 13121
rect 10394 12975 10436 13105
rect 10589 13100 10653 13155
rect 10588 13065 10653 13100
rect 10470 13049 10653 13065
rect 10504 13015 10653 13049
rect 10470 13005 10653 13015
rect 10687 13111 10735 13137
rect 10687 13077 10701 13111
rect 10769 13125 10803 13171
rect 10871 13175 10875 13209
rect 10837 13159 10875 13175
rect 10909 13205 11099 13213
rect 10909 13171 11049 13205
rect 11083 13171 11099 13205
rect 11143 13175 11159 13209
rect 11193 13175 11213 13209
rect 10909 13157 11099 13171
rect 10769 13091 10875 13125
rect 10687 13057 10735 13077
rect 10831 13085 10875 13091
rect 10687 13023 10745 13057
rect 10779 13048 10795 13057
rect 10831 13051 10841 13085
rect 10831 13035 10875 13051
rect 10687 13014 10761 13023
rect 10470 12999 10618 13005
rect 10025 12915 10359 12955
rect 10025 12881 10043 12915
rect 10077 12881 10307 12915
rect 10341 12881 10359 12915
rect 10025 12813 10359 12881
rect 10025 12779 10043 12813
rect 10077 12779 10307 12813
rect 10341 12779 10359 12813
rect 10394 12941 10405 12975
rect 10439 12941 10445 12975
rect 10394 12917 10445 12941
rect 10394 12883 10411 12917
rect 10394 12849 10445 12883
rect 10394 12815 10411 12849
rect 10394 12799 10445 12815
rect 10479 12881 10540 12965
rect 10479 12847 10495 12881
rect 10529 12847 10540 12881
rect 10584 12881 10618 12999
rect 10687 12983 10795 13014
rect 10909 13001 10943 13157
rect 10862 12967 10943 13001
rect 10977 13059 11047 13123
rect 10977 13043 10985 13059
rect 11019 13025 11047 13059
rect 11011 13009 11047 13025
rect 10977 12999 11047 13009
rect 11081 13107 11123 13123
rect 11115 13073 11123 13107
rect 10862 12949 10896 12967
rect 11081 12965 11123 13073
rect 10652 12915 10668 12949
rect 10702 12915 10896 12949
rect 10988 12933 11123 12965
rect 10584 12847 10744 12881
rect 10479 12813 10540 12847
rect 10710 12839 10744 12847
rect 10025 12737 10359 12779
rect 10479 12779 10495 12813
rect 10529 12779 10540 12813
rect 10479 12737 10540 12779
rect 10608 12779 10624 12813
rect 10658 12779 10674 12813
rect 10862 12839 10896 12915
rect 10930 12899 10946 12933
rect 10980 12931 11123 12933
rect 11161 13097 11213 13175
rect 11255 13205 11321 13247
rect 11255 13171 11271 13205
rect 11305 13171 11321 13205
rect 11841 13209 11907 13247
rect 11255 13155 11321 13171
rect 11496 13169 11617 13203
rect 11651 13169 11667 13203
rect 11708 13169 11724 13203
rect 11758 13169 11807 13203
rect 11841 13175 11857 13209
rect 11891 13175 11907 13209
rect 12047 13205 12113 13247
rect 11979 13179 12013 13195
rect 11161 12959 11195 13097
rect 11297 13095 11349 13111
rect 11229 13047 11263 13063
rect 11297 13061 11325 13095
rect 11383 13077 11421 13111
rect 11359 13061 11455 13077
rect 11496 13027 11530 13169
rect 11564 13101 11635 13111
rect 11564 13067 11580 13101
rect 11614 13067 11635 13101
rect 11263 13013 11567 13027
rect 11229 12993 11567 13013
rect 10980 12907 11022 12931
rect 10930 12873 10977 12899
rect 11011 12873 11022 12907
rect 11161 12925 11411 12959
rect 11445 12925 11461 12959
rect 11161 12897 11195 12925
rect 11083 12863 11195 12897
rect 10710 12789 10744 12805
rect 10778 12813 10828 12829
rect 10608 12737 10674 12779
rect 10778 12779 10794 12813
rect 10778 12737 10828 12779
rect 10862 12814 11036 12839
rect 10862 12780 10986 12814
rect 11020 12780 11036 12814
rect 10862 12771 11036 12780
rect 11083 12821 11117 12863
rect 11284 12857 11499 12891
rect 11284 12839 11318 12857
rect 11083 12771 11117 12787
rect 11151 12813 11225 12829
rect 11151 12779 11171 12813
rect 11205 12779 11225 12813
rect 11465 12839 11499 12857
rect 11284 12789 11318 12805
rect 11352 12789 11368 12823
rect 11402 12789 11418 12823
rect 11465 12789 11499 12805
rect 11533 12837 11567 12993
rect 11601 12949 11635 13067
rect 11669 13095 11739 13111
rect 11669 13061 11682 13095
rect 11716 13061 11739 13095
rect 11669 13043 11739 13061
rect 11669 13009 11693 13043
rect 11727 13009 11739 13043
rect 11669 12987 11739 13009
rect 11601 12933 11694 12949
rect 11601 12907 11660 12933
rect 11635 12899 11660 12907
rect 11635 12873 11694 12899
rect 11773 12897 11807 13169
rect 12047 13171 12063 13205
rect 12097 13171 12113 13205
rect 12319 13205 12385 13247
rect 12147 13179 12198 13195
rect 11841 12988 11933 13141
rect 11875 12975 11933 12988
rect 11875 12954 11877 12975
rect 11841 12941 11877 12954
rect 11911 12941 11933 12975
rect 11841 12931 11933 12941
rect 11601 12871 11694 12873
rect 11728 12863 11807 12897
rect 11728 12837 11762 12863
rect 11533 12815 11669 12837
rect 11151 12737 11225 12779
rect 11352 12737 11418 12789
rect 11533 12781 11619 12815
rect 11653 12781 11669 12815
rect 11533 12771 11669 12781
rect 11712 12821 11762 12837
rect 11746 12787 11762 12821
rect 11712 12771 11762 12787
rect 11796 12813 11846 12829
rect 11830 12779 11846 12813
rect 11796 12737 11846 12779
rect 11880 12774 11945 12931
rect 11979 12907 12013 13145
rect 12181 13145 12198 13179
rect 12147 13137 12198 13145
rect 12048 13103 12198 13137
rect 12234 13179 12285 13195
rect 12234 13145 12251 13179
rect 12319 13171 12335 13205
rect 12369 13171 12385 13205
rect 12525 13209 12591 13247
rect 12419 13179 12453 13195
rect 12234 13137 12285 13145
rect 12525 13175 12541 13209
rect 12575 13175 12591 13209
rect 13111 13205 13177 13247
rect 12234 13103 12384 13137
rect 12048 13043 12094 13103
rect 12048 13034 12060 13043
rect 12082 13000 12094 13009
rect 12048 12905 12094 13000
rect 12128 13049 12198 13069
rect 12128 13015 12150 13049
rect 12184 13043 12198 13049
rect 12128 13009 12153 13015
rect 12187 13009 12198 13043
rect 12128 12939 12198 13009
rect 12234 13049 12304 13069
rect 12234 13043 12248 13049
rect 12234 13009 12245 13043
rect 12282 13015 12304 13049
rect 12279 13009 12304 13015
rect 12234 12939 12304 13009
rect 12338 13043 12384 13103
rect 12372 13034 12384 13043
rect 12338 13000 12350 13009
rect 12338 12905 12384 13000
rect 12048 12889 12198 12905
rect 12048 12871 12147 12889
rect 11979 12821 12013 12855
rect 12181 12855 12198 12889
rect 11979 12771 12013 12787
rect 12047 12803 12063 12837
rect 12097 12803 12113 12837
rect 12047 12737 12113 12803
rect 12147 12821 12198 12855
rect 12181 12787 12198 12821
rect 12147 12771 12198 12787
rect 12234 12889 12384 12905
rect 12234 12855 12251 12889
rect 12285 12871 12384 12889
rect 12419 12907 12453 13145
rect 12625 13169 12674 13203
rect 12708 13169 12724 13203
rect 12765 13169 12781 13203
rect 12815 13169 12936 13203
rect 12499 12988 12591 13141
rect 12499 12975 12557 12988
rect 12499 12941 12521 12975
rect 12555 12954 12557 12975
rect 12555 12941 12591 12954
rect 12499 12931 12591 12941
rect 12234 12821 12285 12855
rect 12234 12787 12251 12821
rect 12234 12771 12285 12787
rect 12319 12803 12335 12837
rect 12369 12803 12385 12837
rect 12319 12737 12385 12803
rect 12419 12821 12453 12855
rect 12419 12771 12453 12787
rect 12487 12774 12552 12931
rect 12625 12897 12659 13169
rect 12693 13095 12763 13111
rect 12693 13061 12716 13095
rect 12750 13061 12763 13095
rect 12693 13043 12763 13061
rect 12693 13009 12705 13043
rect 12739 13009 12763 13043
rect 12693 12987 12763 13009
rect 12797 13101 12868 13111
rect 12797 13067 12818 13101
rect 12852 13067 12868 13101
rect 12797 12949 12831 13067
rect 12902 13027 12936 13169
rect 13111 13171 13127 13205
rect 13161 13171 13177 13205
rect 13111 13155 13177 13171
rect 13219 13175 13239 13209
rect 13273 13175 13289 13209
rect 13333 13205 13523 13213
rect 13011 13077 13049 13111
rect 13083 13095 13135 13111
rect 13219 13097 13271 13175
rect 13333 13171 13349 13205
rect 13383 13171 13523 13205
rect 13333 13157 13523 13171
rect 13557 13209 13595 13247
rect 13557 13175 13561 13209
rect 13892 13205 13953 13247
rect 13557 13159 13595 13175
rect 13629 13189 13843 13205
rect 13629 13171 13779 13189
rect 12977 13061 13073 13077
rect 13107 13061 13135 13095
rect 13169 13047 13203 13063
rect 12738 12933 12831 12949
rect 12772 12907 12831 12933
rect 12772 12899 12797 12907
rect 12625 12863 12704 12897
rect 12738 12873 12797 12899
rect 12738 12871 12831 12873
rect 12865 13013 13169 13027
rect 12865 12993 13203 13013
rect 12670 12837 12704 12863
rect 12865 12837 12899 12993
rect 13237 12959 13271 13097
rect 12971 12925 12987 12959
rect 13021 12925 13271 12959
rect 13309 13107 13351 13123
rect 13309 13073 13317 13107
rect 13309 12965 13351 13073
rect 13385 13059 13455 13123
rect 13385 13025 13413 13059
rect 13447 13043 13455 13059
rect 13385 13009 13421 13025
rect 13385 12999 13455 13009
rect 13489 13001 13523 13157
rect 13629 13125 13663 13171
rect 13813 13155 13843 13189
rect 13892 13171 13903 13205
rect 13937 13171 13953 13205
rect 13892 13155 13953 13171
rect 13987 13155 14038 13211
rect 13557 13091 13663 13125
rect 13697 13111 13745 13137
rect 13557 13085 13601 13091
rect 13591 13051 13601 13085
rect 13731 13077 13745 13111
rect 13697 13057 13745 13077
rect 13557 13035 13601 13051
rect 13637 13048 13653 13057
rect 13687 13023 13745 13057
rect 13671 13014 13745 13023
rect 13489 12967 13570 13001
rect 13637 12983 13745 13014
rect 13779 13100 13843 13155
rect 14021 13121 14038 13155
rect 13987 13105 14038 13121
rect 13779 13065 13844 13100
rect 13779 13049 13962 13065
rect 13779 13015 13928 13049
rect 13779 13005 13962 13015
rect 13814 12999 13962 13005
rect 13309 12933 13444 12965
rect 13536 12949 13570 12967
rect 13309 12931 13452 12933
rect 13237 12897 13271 12925
rect 13410 12907 13452 12931
rect 12586 12813 12636 12829
rect 12586 12779 12602 12813
rect 12586 12737 12636 12779
rect 12670 12821 12720 12837
rect 12670 12787 12686 12821
rect 12670 12771 12720 12787
rect 12763 12815 12899 12837
rect 12763 12781 12779 12815
rect 12813 12781 12899 12815
rect 12933 12857 13148 12891
rect 13237 12863 13349 12897
rect 13410 12873 13421 12907
rect 13486 12899 13502 12933
rect 13455 12873 13502 12899
rect 13536 12915 13730 12949
rect 13764 12915 13780 12949
rect 12933 12839 12967 12857
rect 13114 12839 13148 12857
rect 12933 12789 12967 12805
rect 13014 12789 13030 12823
rect 13064 12789 13080 12823
rect 13114 12789 13148 12805
rect 13207 12813 13281 12829
rect 12763 12771 12899 12781
rect 13014 12737 13080 12789
rect 13207 12779 13227 12813
rect 13261 12779 13281 12813
rect 13207 12737 13281 12779
rect 13315 12821 13349 12863
rect 13536 12839 13570 12915
rect 13814 12881 13848 12999
rect 13996 12975 14038 13105
rect 13315 12771 13349 12787
rect 13396 12814 13570 12839
rect 13688 12847 13848 12881
rect 13892 12881 13953 12965
rect 13892 12847 13903 12881
rect 13937 12847 13953 12881
rect 13688 12839 13722 12847
rect 13396 12780 13412 12814
rect 13446 12780 13570 12814
rect 13396 12771 13570 12780
rect 13604 12813 13654 12829
rect 13638 12779 13654 12813
rect 13892 12813 13953 12847
rect 13688 12789 13722 12805
rect 13604 12737 13654 12779
rect 13758 12779 13774 12813
rect 13808 12779 13824 12813
rect 13758 12737 13824 12779
rect 13892 12779 13903 12813
rect 13937 12779 13953 12813
rect 13987 12917 14038 12975
rect 14021 12883 14038 12917
rect 13987 12849 14038 12883
rect 14021 12839 14038 12849
rect 13987 12805 13993 12815
rect 14027 12805 14038 12839
rect 13987 12799 14038 12805
rect 14074 13186 14125 13213
rect 14074 13152 14091 13186
rect 14159 13205 14225 13247
rect 14159 13171 14175 13205
rect 14209 13171 14225 13205
rect 14159 13167 14225 13171
rect 14310 13190 14416 13213
rect 14074 13099 14125 13152
rect 14310 13156 14382 13190
rect 14310 13140 14416 13156
rect 14310 13133 14345 13140
rect 14159 13099 14345 13133
rect 14074 12965 14108 13099
rect 14159 13065 14193 13099
rect 14142 13049 14193 13065
rect 14176 13015 14193 13049
rect 14142 12999 14193 13015
rect 14238 13049 14277 13065
rect 14272 13015 14277 13049
rect 14238 12999 14277 13015
rect 14074 12949 14141 12965
rect 14074 12915 14091 12949
rect 14125 12915 14141 12949
rect 14074 12907 14141 12915
rect 14074 12873 14085 12907
rect 14119 12881 14141 12907
rect 14074 12847 14091 12873
rect 14125 12847 14141 12881
rect 14074 12813 14141 12847
rect 13892 12737 13953 12779
rect 14074 12779 14091 12813
rect 14125 12779 14141 12813
rect 14074 12771 14141 12779
rect 14175 12949 14209 12965
rect 14175 12881 14209 12915
rect 14175 12813 14209 12847
rect 14175 12737 14209 12779
rect 14243 12805 14277 12999
rect 14311 12873 14345 13099
rect 14379 13085 14413 13101
rect 14379 12941 14413 13051
rect 14454 13085 14509 13213
rect 14454 13051 14475 13085
rect 14454 13043 14509 13051
rect 14487 13009 14509 13043
rect 14454 12981 14509 13009
rect 14543 13111 14581 13213
rect 14617 13190 14719 13247
rect 14651 13156 14685 13190
rect 14617 13140 14719 13156
rect 14763 13190 14812 13206
rect 14763 13156 14769 13190
rect 14803 13156 14812 13190
rect 14543 13077 14545 13111
rect 14579 13077 14581 13111
rect 14763 13085 14812 13156
rect 14993 13153 15051 13247
rect 14993 13119 15005 13153
rect 15039 13119 15051 13153
rect 14993 13102 15051 13119
rect 15086 13155 15137 13211
rect 15171 13205 15232 13247
rect 15529 13209 15567 13247
rect 15171 13171 15187 13205
rect 15221 13171 15232 13205
rect 15171 13155 15232 13171
rect 15281 13189 15495 13205
rect 15281 13155 15311 13189
rect 15345 13171 15495 13189
rect 15086 13121 15103 13155
rect 15086 13105 15137 13121
rect 14543 12972 14581 13077
rect 14621 13051 14637 13085
rect 14671 13051 14867 13085
rect 14543 12941 14547 12972
rect 14379 12938 14547 12941
rect 14379 12907 14581 12938
rect 14615 12975 14765 12976
rect 14615 12972 14729 12975
rect 14615 12938 14715 12972
rect 14763 12941 14765 12975
rect 14749 12938 14765 12941
rect 14311 12839 14411 12873
rect 14445 12839 14486 12873
rect 14520 12839 14536 12873
rect 14615 12805 14649 12938
rect 14799 12889 14867 13051
rect 15086 12975 15128 13105
rect 15281 13100 15345 13155
rect 15280 13065 15345 13100
rect 15162 13049 15345 13065
rect 15196 13015 15345 13049
rect 15162 13005 15345 13015
rect 15379 13111 15427 13137
rect 15379 13077 15393 13111
rect 15461 13125 15495 13171
rect 15563 13175 15567 13209
rect 15529 13159 15567 13175
rect 15601 13205 15791 13213
rect 15601 13171 15741 13205
rect 15775 13171 15791 13205
rect 15835 13175 15851 13209
rect 15885 13175 15905 13209
rect 15601 13157 15791 13171
rect 15461 13091 15567 13125
rect 15379 13057 15427 13077
rect 15523 13085 15567 13091
rect 15379 13023 15437 13057
rect 15471 13048 15487 13057
rect 15523 13051 15533 13085
rect 15523 13035 15567 13051
rect 15379 13014 15453 13023
rect 15162 12999 15310 13005
rect 14243 12771 14649 12805
rect 14683 12873 14717 12889
rect 14683 12737 14717 12839
rect 14764 12873 14867 12889
rect 14764 12839 14769 12873
rect 14803 12839 14867 12873
rect 14764 12807 14867 12839
rect 14993 12935 15051 12970
rect 14993 12901 15005 12935
rect 15039 12901 15051 12935
rect 14993 12842 15051 12901
rect 14993 12808 15005 12842
rect 15039 12808 15051 12842
rect 14993 12737 15051 12808
rect 15086 12917 15137 12975
rect 15086 12883 15103 12917
rect 15086 12849 15137 12883
rect 15086 12839 15103 12849
rect 15086 12805 15097 12839
rect 15131 12805 15137 12815
rect 15086 12799 15137 12805
rect 15171 12881 15232 12965
rect 15171 12847 15187 12881
rect 15221 12847 15232 12881
rect 15276 12881 15310 12999
rect 15379 12983 15487 13014
rect 15601 13001 15635 13157
rect 15554 12967 15635 13001
rect 15669 13059 15739 13123
rect 15669 13043 15677 13059
rect 15711 13025 15739 13059
rect 15703 13009 15739 13025
rect 15669 12999 15739 13009
rect 15773 13107 15815 13123
rect 15807 13073 15815 13107
rect 15554 12949 15588 12967
rect 15773 12965 15815 13073
rect 15344 12915 15360 12949
rect 15394 12915 15588 12949
rect 15680 12933 15815 12965
rect 15276 12847 15436 12881
rect 15171 12813 15232 12847
rect 15402 12839 15436 12847
rect 15171 12779 15187 12813
rect 15221 12779 15232 12813
rect 15171 12737 15232 12779
rect 15300 12779 15316 12813
rect 15350 12779 15366 12813
rect 15554 12839 15588 12915
rect 15622 12899 15638 12933
rect 15672 12931 15815 12933
rect 15853 13097 15905 13175
rect 15947 13205 16013 13247
rect 15947 13171 15963 13205
rect 15997 13171 16013 13205
rect 16533 13209 16599 13247
rect 15947 13155 16013 13171
rect 16188 13169 16309 13203
rect 16343 13169 16359 13203
rect 16400 13169 16416 13203
rect 16450 13169 16499 13203
rect 16533 13175 16549 13209
rect 16583 13175 16599 13209
rect 16739 13205 16805 13247
rect 16671 13179 16705 13195
rect 15853 12959 15887 13097
rect 15989 13095 16041 13111
rect 15921 13047 15955 13063
rect 15989 13061 16017 13095
rect 16075 13077 16113 13111
rect 16051 13061 16147 13077
rect 16188 13027 16222 13169
rect 16256 13101 16327 13111
rect 16256 13067 16272 13101
rect 16306 13067 16327 13101
rect 15955 13013 16259 13027
rect 15921 12993 16259 13013
rect 15672 12907 15714 12931
rect 15622 12873 15669 12899
rect 15703 12873 15714 12907
rect 15853 12925 16103 12959
rect 16137 12925 16153 12959
rect 15853 12897 15887 12925
rect 15775 12863 15887 12897
rect 15402 12789 15436 12805
rect 15470 12813 15520 12829
rect 15300 12737 15366 12779
rect 15470 12779 15486 12813
rect 15470 12737 15520 12779
rect 15554 12814 15728 12839
rect 15554 12780 15678 12814
rect 15712 12780 15728 12814
rect 15554 12771 15728 12780
rect 15775 12821 15809 12863
rect 15976 12857 16191 12891
rect 15976 12839 16010 12857
rect 15775 12771 15809 12787
rect 15843 12813 15917 12829
rect 15843 12779 15863 12813
rect 15897 12779 15917 12813
rect 16157 12839 16191 12857
rect 15976 12789 16010 12805
rect 16044 12789 16060 12823
rect 16094 12789 16110 12823
rect 16157 12789 16191 12805
rect 16225 12837 16259 12993
rect 16293 12949 16327 13067
rect 16361 13095 16431 13111
rect 16361 13061 16374 13095
rect 16408 13061 16431 13095
rect 16361 13043 16431 13061
rect 16361 13009 16385 13043
rect 16419 13009 16431 13043
rect 16361 12987 16431 13009
rect 16293 12933 16386 12949
rect 16293 12907 16352 12933
rect 16327 12899 16352 12907
rect 16327 12873 16386 12899
rect 16465 12897 16499 13169
rect 16739 13171 16755 13205
rect 16789 13171 16805 13205
rect 16839 13179 16890 13195
rect 16533 12988 16625 13141
rect 16567 12975 16625 12988
rect 16567 12954 16569 12975
rect 16533 12941 16569 12954
rect 16603 12941 16625 12975
rect 16533 12931 16625 12941
rect 16293 12871 16386 12873
rect 16420 12863 16499 12897
rect 16420 12837 16454 12863
rect 16225 12815 16361 12837
rect 15843 12737 15917 12779
rect 16044 12737 16110 12789
rect 16225 12781 16311 12815
rect 16345 12781 16361 12815
rect 16225 12771 16361 12781
rect 16404 12821 16454 12837
rect 16438 12787 16454 12821
rect 16404 12771 16454 12787
rect 16488 12813 16538 12829
rect 16522 12779 16538 12813
rect 16488 12737 16538 12779
rect 16572 12774 16637 12931
rect 16671 12907 16705 13145
rect 16873 13145 16890 13179
rect 16839 13137 16890 13145
rect 16740 13103 16890 13137
rect 16925 13179 17002 13213
rect 16925 13145 16937 13179
rect 16996 13145 17002 13179
rect 17036 13205 17101 13247
rect 17036 13171 17052 13205
rect 17086 13171 17101 13205
rect 17036 13155 17101 13171
rect 17205 13179 17261 13213
rect 16740 13043 16786 13103
rect 16925 13099 17002 13145
rect 17205 13145 17211 13179
rect 17245 13145 17261 13179
rect 17205 13121 17261 13145
rect 16740 13034 16752 13043
rect 16774 13000 16786 13009
rect 16740 12905 16786 13000
rect 16820 13049 16890 13069
rect 16820 13015 16842 13049
rect 16876 13043 16890 13049
rect 16820 13009 16845 13015
rect 16879 13009 16890 13043
rect 16820 12939 16890 13009
rect 16925 12965 16981 13099
rect 17036 13087 17261 13121
rect 17299 13179 17379 13213
rect 17299 13145 17315 13179
rect 17349 13145 17379 13179
rect 17459 13205 17513 13247
rect 17459 13171 17469 13205
rect 17503 13171 17513 13205
rect 17459 13155 17513 13171
rect 17547 13179 17604 13213
rect 17036 13065 17126 13087
rect 17015 13049 17126 13065
rect 17299 13053 17379 13145
rect 17547 13145 17553 13179
rect 17587 13145 17604 13179
rect 17547 13121 17604 13145
rect 17754 13186 18823 13247
rect 17754 13152 17771 13186
rect 17805 13152 18771 13186
rect 18805 13152 18823 13186
rect 17754 13138 18823 13152
rect 18858 13186 19927 13247
rect 18858 13152 18875 13186
rect 18909 13152 19875 13186
rect 19909 13152 19927 13186
rect 18858 13138 19927 13152
rect 19961 13184 20203 13247
rect 19961 13150 19979 13184
rect 20013 13150 20151 13184
rect 20185 13150 20203 13184
rect 17049 13015 17126 13049
rect 17015 12999 17126 13015
rect 16740 12889 16890 12905
rect 16740 12871 16839 12889
rect 16671 12821 16705 12855
rect 16873 12855 16890 12889
rect 16671 12771 16705 12787
rect 16739 12803 16755 12837
rect 16789 12803 16805 12837
rect 16739 12737 16805 12803
rect 16839 12821 16890 12855
rect 16873 12787 16890 12821
rect 16839 12771 16890 12787
rect 16925 12839 17002 12965
rect 17036 12907 17126 12999
rect 17160 13049 17379 13053
rect 17160 13015 17211 13049
rect 17245 13015 17379 13049
rect 17160 12941 17379 13015
rect 17036 12863 17261 12907
rect 16925 12805 16962 12839
rect 16996 12805 17002 12839
rect 17205 12839 17261 12863
rect 16925 12771 17002 12805
rect 17036 12813 17101 12829
rect 17036 12779 17052 12813
rect 17086 12779 17101 12813
rect 17036 12737 17101 12779
rect 17205 12805 17211 12839
rect 17245 12805 17261 12839
rect 17205 12771 17261 12805
rect 17299 12839 17379 12941
rect 17413 13087 17604 13121
rect 17413 13049 17455 13087
rect 18072 13059 18142 13074
rect 17413 13015 17415 13049
rect 17449 13015 17455 13049
rect 17413 12907 17455 13015
rect 17489 13049 17627 13053
rect 17489 13015 17529 13049
rect 17563 13015 17627 13049
rect 17489 12975 17627 13015
rect 17489 12941 17581 12975
rect 17615 12941 17627 12975
rect 18072 13025 18091 13059
rect 18125 13025 18142 13059
rect 17413 12863 17604 12907
rect 17299 12805 17315 12839
rect 17349 12805 17379 12839
rect 17547 12839 17604 12863
rect 17299 12771 17379 12805
rect 17459 12813 17513 12829
rect 17459 12779 17469 12813
rect 17503 12779 17513 12813
rect 17459 12737 17513 12779
rect 17547 12805 17553 12839
rect 17587 12805 17604 12839
rect 18072 12824 18142 13025
rect 18438 13023 18506 13138
rect 18438 12989 18455 13023
rect 18489 12989 18506 13023
rect 18438 12972 18506 12989
rect 19176 13059 19246 13074
rect 19176 13025 19195 13059
rect 19229 13025 19246 13059
rect 19176 12824 19246 13025
rect 19542 13023 19610 13138
rect 19961 13097 20203 13150
rect 19542 12989 19559 13023
rect 19593 12989 19610 13023
rect 19542 12972 19610 12989
rect 19961 13029 20011 13063
rect 20045 13029 20065 13063
rect 19961 12955 20065 13029
rect 20099 13023 20203 13097
rect 20099 12989 20119 13023
rect 20153 12989 20203 13023
rect 19961 12908 20203 12955
rect 19961 12874 19979 12908
rect 20013 12874 20151 12908
rect 20185 12874 20203 12908
rect 17547 12771 17604 12805
rect 17754 12813 18823 12824
rect 17754 12779 17771 12813
rect 17805 12779 18771 12813
rect 18805 12779 18823 12813
rect 17754 12737 18823 12779
rect 18858 12813 19927 12824
rect 18858 12779 18875 12813
rect 18909 12779 19875 12813
rect 19909 12779 19927 12813
rect 18858 12737 19927 12779
rect 19961 12813 20203 12874
rect 19961 12779 19979 12813
rect 20013 12779 20151 12813
rect 20185 12779 20203 12813
rect 19961 12737 20203 12779
rect 4948 12703 4977 12737
rect 5011 12703 5069 12737
rect 5103 12703 5161 12737
rect 5195 12703 5253 12737
rect 5287 12703 5345 12737
rect 5379 12703 5437 12737
rect 5471 12703 5529 12737
rect 5563 12703 5621 12737
rect 5655 12703 5713 12737
rect 5747 12703 5805 12737
rect 5839 12703 5897 12737
rect 5931 12703 5989 12737
rect 6023 12703 6081 12737
rect 6115 12703 6173 12737
rect 6207 12703 6265 12737
rect 6299 12703 6357 12737
rect 6391 12703 6449 12737
rect 6483 12703 6541 12737
rect 6575 12703 6633 12737
rect 6667 12703 6725 12737
rect 6759 12703 6817 12737
rect 6851 12703 6909 12737
rect 6943 12703 7001 12737
rect 7035 12703 7093 12737
rect 7127 12703 7185 12737
rect 7219 12703 7277 12737
rect 7311 12703 7369 12737
rect 7403 12703 7461 12737
rect 7495 12703 7553 12737
rect 7587 12703 7645 12737
rect 7679 12703 7737 12737
rect 7771 12703 7829 12737
rect 7863 12703 7921 12737
rect 7955 12703 8013 12737
rect 8047 12703 8105 12737
rect 8139 12703 8197 12737
rect 8231 12703 8289 12737
rect 8323 12703 8381 12737
rect 8415 12703 8473 12737
rect 8507 12703 8565 12737
rect 8599 12703 8657 12737
rect 8691 12703 8749 12737
rect 8783 12703 8841 12737
rect 8875 12703 8933 12737
rect 8967 12703 9025 12737
rect 9059 12703 9117 12737
rect 9151 12703 9209 12737
rect 9243 12703 9301 12737
rect 9335 12703 9393 12737
rect 9427 12703 9485 12737
rect 9519 12703 9577 12737
rect 9611 12703 9669 12737
rect 9703 12703 9761 12737
rect 9795 12703 9853 12737
rect 9887 12703 9945 12737
rect 9979 12703 10037 12737
rect 10071 12703 10129 12737
rect 10163 12703 10221 12737
rect 10255 12703 10313 12737
rect 10347 12703 10405 12737
rect 10439 12703 10497 12737
rect 10531 12703 10589 12737
rect 10623 12703 10681 12737
rect 10715 12703 10773 12737
rect 10807 12703 10865 12737
rect 10899 12703 10957 12737
rect 10991 12703 11049 12737
rect 11083 12703 11141 12737
rect 11175 12703 11233 12737
rect 11267 12703 11325 12737
rect 11359 12703 11417 12737
rect 11451 12703 11509 12737
rect 11543 12703 11601 12737
rect 11635 12703 11693 12737
rect 11727 12703 11785 12737
rect 11819 12703 11877 12737
rect 11911 12703 11969 12737
rect 12003 12703 12061 12737
rect 12095 12703 12153 12737
rect 12187 12703 12245 12737
rect 12279 12703 12337 12737
rect 12371 12703 12429 12737
rect 12463 12703 12521 12737
rect 12555 12703 12613 12737
rect 12647 12703 12705 12737
rect 12739 12703 12797 12737
rect 12831 12703 12889 12737
rect 12923 12703 12981 12737
rect 13015 12703 13073 12737
rect 13107 12703 13165 12737
rect 13199 12703 13257 12737
rect 13291 12703 13349 12737
rect 13383 12703 13441 12737
rect 13475 12703 13533 12737
rect 13567 12703 13625 12737
rect 13659 12703 13717 12737
rect 13751 12703 13809 12737
rect 13843 12703 13901 12737
rect 13935 12703 13993 12737
rect 14027 12703 14085 12737
rect 14119 12703 14177 12737
rect 14211 12703 14269 12737
rect 14303 12703 14361 12737
rect 14395 12703 14453 12737
rect 14487 12703 14545 12737
rect 14579 12703 14637 12737
rect 14671 12703 14729 12737
rect 14763 12703 14821 12737
rect 14855 12703 14913 12737
rect 14947 12703 15005 12737
rect 15039 12703 15097 12737
rect 15131 12703 15189 12737
rect 15223 12703 15281 12737
rect 15315 12703 15373 12737
rect 15407 12703 15465 12737
rect 15499 12703 15557 12737
rect 15591 12703 15649 12737
rect 15683 12703 15741 12737
rect 15775 12703 15833 12737
rect 15867 12703 15925 12737
rect 15959 12703 16017 12737
rect 16051 12703 16109 12737
rect 16143 12703 16201 12737
rect 16235 12703 16293 12737
rect 16327 12703 16385 12737
rect 16419 12703 16477 12737
rect 16511 12703 16569 12737
rect 16603 12703 16661 12737
rect 16695 12703 16753 12737
rect 16787 12703 16845 12737
rect 16879 12703 16937 12737
rect 16971 12703 17029 12737
rect 17063 12703 17121 12737
rect 17155 12703 17213 12737
rect 17247 12703 17305 12737
rect 17339 12703 17397 12737
rect 17431 12703 17489 12737
rect 17523 12703 17581 12737
rect 17615 12703 17673 12737
rect 17707 12703 17765 12737
rect 17799 12703 17857 12737
rect 17891 12703 17949 12737
rect 17983 12703 18041 12737
rect 18075 12703 18133 12737
rect 18167 12703 18225 12737
rect 18259 12703 18317 12737
rect 18351 12703 18409 12737
rect 18443 12703 18501 12737
rect 18535 12703 18593 12737
rect 18627 12703 18685 12737
rect 18719 12703 18777 12737
rect 18811 12703 18869 12737
rect 18903 12703 18961 12737
rect 18995 12703 19053 12737
rect 19087 12703 19145 12737
rect 19179 12703 19237 12737
rect 19271 12703 19329 12737
rect 19363 12703 19421 12737
rect 19455 12703 19513 12737
rect 19547 12703 19605 12737
rect 19639 12703 19697 12737
rect 19731 12703 19789 12737
rect 19823 12703 19881 12737
rect 19915 12703 19973 12737
rect 20007 12703 20065 12737
rect 20099 12703 20157 12737
rect 20191 12703 20220 12737
rect 4965 12661 5207 12703
rect 4965 12627 4983 12661
rect 5017 12627 5155 12661
rect 5189 12627 5207 12661
rect 4965 12566 5207 12627
rect 4965 12532 4983 12566
rect 5017 12532 5155 12566
rect 5189 12532 5207 12566
rect 4965 12485 5207 12532
rect 4965 12417 5015 12451
rect 5049 12417 5069 12451
rect 4965 12343 5069 12417
rect 5103 12411 5207 12485
rect 5103 12377 5123 12411
rect 5157 12377 5207 12411
rect 5241 12660 5345 12669
rect 5241 12626 5295 12660
rect 5329 12626 5345 12660
rect 5241 12592 5345 12626
rect 5241 12558 5295 12592
rect 5329 12558 5345 12592
rect 5379 12660 5445 12703
rect 5379 12626 5395 12660
rect 5429 12626 5445 12660
rect 5379 12592 5445 12626
rect 5610 12661 6679 12703
rect 5610 12627 5627 12661
rect 5661 12627 6627 12661
rect 6661 12627 6679 12661
rect 5610 12616 6679 12627
rect 6724 12647 6781 12703
rect 5379 12558 5395 12592
rect 5429 12558 5445 12592
rect 5241 12431 5345 12558
rect 5241 12397 5253 12431
rect 5287 12397 5345 12431
rect 5241 12359 5345 12397
rect 4965 12290 5207 12343
rect 5379 12329 5483 12524
rect 5928 12415 5998 12616
rect 6724 12613 6739 12647
rect 6773 12613 6781 12647
rect 6724 12579 6781 12613
rect 6724 12545 6739 12579
rect 6773 12545 6781 12579
rect 6724 12529 6781 12545
rect 6815 12653 6867 12669
rect 6815 12619 6825 12653
rect 6859 12619 6867 12653
rect 6815 12585 6867 12619
rect 6902 12661 6953 12703
rect 6902 12627 6911 12661
rect 6945 12627 6953 12661
rect 6902 12611 6953 12627
rect 6987 12626 7039 12669
rect 6815 12551 6825 12585
rect 6859 12577 6867 12585
rect 6987 12592 6997 12626
rect 7031 12592 7039 12626
rect 6987 12577 7039 12592
rect 6859 12551 7039 12577
rect 6815 12543 7039 12551
rect 7073 12661 7135 12703
rect 7073 12627 7093 12661
rect 7127 12627 7135 12661
rect 7073 12593 7135 12627
rect 7073 12559 7093 12593
rect 7127 12559 7135 12593
rect 7073 12543 7135 12559
rect 7169 12653 7231 12669
rect 7169 12619 7179 12653
rect 7213 12619 7231 12653
rect 6815 12517 6867 12543
rect 6815 12493 6825 12517
rect 6716 12483 6825 12493
rect 6859 12483 6867 12517
rect 7169 12531 7231 12619
rect 7169 12509 7179 12531
rect 5928 12381 5947 12415
rect 5981 12381 5998 12415
rect 5928 12366 5998 12381
rect 6294 12451 6362 12468
rect 6294 12417 6311 12451
rect 6345 12417 6362 12451
rect 4965 12256 4983 12290
rect 5017 12256 5155 12290
rect 5189 12256 5207 12290
rect 4965 12193 5207 12256
rect 5277 12291 5295 12325
rect 5329 12291 5345 12325
rect 5277 12257 5345 12291
rect 5277 12223 5295 12257
rect 5329 12223 5345 12257
rect 5379 12295 5395 12329
rect 5429 12295 5483 12329
rect 6294 12302 6362 12417
rect 6716 12459 6867 12483
rect 7025 12497 7179 12509
rect 7213 12497 7231 12531
rect 7025 12475 7231 12497
rect 6716 12357 6797 12459
rect 7025 12425 7059 12475
rect 6831 12391 6847 12425
rect 6881 12391 6915 12425
rect 6949 12391 6983 12425
rect 7017 12391 7059 12425
rect 7093 12425 7163 12441
rect 7093 12391 7129 12425
rect 7093 12363 7163 12391
rect 6716 12323 7046 12357
rect 7127 12329 7163 12363
rect 7093 12327 7163 12329
rect 5379 12261 5483 12295
rect 5379 12227 5395 12261
rect 5429 12227 5483 12261
rect 5610 12288 6679 12302
rect 6815 12295 6867 12323
rect 5610 12254 5627 12288
rect 5661 12254 6627 12288
rect 6661 12254 6679 12288
rect 5277 12193 5345 12223
rect 5610 12193 6679 12254
rect 6725 12273 6781 12289
rect 6725 12239 6738 12273
rect 6772 12239 6781 12273
rect 6815 12261 6824 12295
rect 6858 12261 6867 12295
rect 6987 12295 7046 12323
rect 6815 12245 6867 12261
rect 6902 12273 6953 12289
rect 6725 12193 6781 12239
rect 6902 12239 6910 12273
rect 6944 12239 6953 12273
rect 6987 12261 6996 12295
rect 7035 12261 7046 12295
rect 7197 12293 7231 12475
rect 7265 12632 7323 12703
rect 7265 12598 7277 12632
rect 7311 12598 7323 12632
rect 7265 12539 7323 12598
rect 7265 12505 7277 12539
rect 7311 12505 7323 12539
rect 7265 12470 7323 12505
rect 7357 12661 7691 12703
rect 7357 12627 7375 12661
rect 7409 12627 7639 12661
rect 7673 12627 7691 12661
rect 7357 12559 7691 12627
rect 7726 12661 8795 12703
rect 7726 12627 7743 12661
rect 7777 12627 8743 12661
rect 8777 12627 8795 12661
rect 7726 12616 8795 12627
rect 8840 12647 8897 12703
rect 7357 12525 7375 12559
rect 7409 12525 7639 12559
rect 7673 12525 7691 12559
rect 7357 12485 7691 12525
rect 7357 12415 7507 12485
rect 7357 12381 7377 12415
rect 7411 12381 7507 12415
rect 7541 12417 7637 12451
rect 7671 12417 7691 12451
rect 7541 12347 7691 12417
rect 8044 12415 8114 12616
rect 8840 12613 8855 12647
rect 8889 12613 8897 12647
rect 8840 12579 8897 12613
rect 8840 12545 8855 12579
rect 8889 12545 8897 12579
rect 8840 12529 8897 12545
rect 8931 12653 8983 12669
rect 8931 12619 8941 12653
rect 8975 12619 8983 12653
rect 8931 12585 8983 12619
rect 9018 12661 9069 12703
rect 9018 12627 9027 12661
rect 9061 12627 9069 12661
rect 9018 12611 9069 12627
rect 9103 12626 9155 12669
rect 8931 12551 8941 12585
rect 8975 12577 8983 12585
rect 9103 12592 9113 12626
rect 9147 12592 9155 12626
rect 9103 12577 9155 12592
rect 8975 12551 9155 12577
rect 8931 12543 9155 12551
rect 9189 12661 9251 12703
rect 9189 12627 9209 12661
rect 9243 12627 9251 12661
rect 9189 12593 9251 12627
rect 9189 12559 9209 12593
rect 9243 12559 9251 12593
rect 9189 12543 9251 12559
rect 9285 12653 9347 12669
rect 9285 12619 9295 12653
rect 9329 12619 9347 12653
rect 8931 12517 8983 12543
rect 8931 12493 8941 12517
rect 8832 12483 8941 12493
rect 8975 12483 8983 12517
rect 9285 12531 9347 12619
rect 9285 12509 9295 12531
rect 8044 12381 8063 12415
rect 8097 12381 8114 12415
rect 8044 12366 8114 12381
rect 8410 12451 8478 12468
rect 8410 12417 8427 12451
rect 8461 12417 8478 12451
rect 6987 12245 7046 12261
rect 7082 12273 7137 12289
rect 6902 12193 6953 12239
rect 7082 12239 7093 12273
rect 7127 12239 7137 12273
rect 7082 12193 7137 12239
rect 7171 12277 7231 12293
rect 7171 12243 7179 12277
rect 7213 12243 7231 12277
rect 7171 12227 7231 12243
rect 7265 12321 7323 12338
rect 7265 12287 7277 12321
rect 7311 12287 7323 12321
rect 7265 12193 7323 12287
rect 7357 12295 7691 12347
rect 8410 12302 8478 12417
rect 8832 12459 8983 12483
rect 9141 12497 9295 12509
rect 9329 12497 9347 12531
rect 9141 12475 9347 12497
rect 8832 12357 8913 12459
rect 9141 12425 9175 12475
rect 8947 12391 8963 12425
rect 8997 12391 9031 12425
rect 9065 12391 9099 12425
rect 9133 12391 9175 12425
rect 9209 12431 9279 12441
rect 9243 12425 9279 12431
rect 9243 12397 9245 12425
rect 9209 12391 9245 12397
rect 8832 12323 9162 12357
rect 9209 12327 9279 12391
rect 7357 12261 7375 12295
rect 7409 12261 7639 12295
rect 7673 12261 7691 12295
rect 7357 12193 7691 12261
rect 7726 12288 8795 12302
rect 8931 12295 8983 12323
rect 7726 12254 7743 12288
rect 7777 12254 8743 12288
rect 8777 12254 8795 12288
rect 7726 12193 8795 12254
rect 8841 12273 8897 12289
rect 8841 12239 8854 12273
rect 8888 12239 8897 12273
rect 8931 12261 8940 12295
rect 8974 12261 8983 12295
rect 9103 12295 9162 12323
rect 8931 12245 8983 12261
rect 9018 12273 9069 12289
rect 8841 12193 8897 12239
rect 9018 12239 9026 12273
rect 9060 12239 9069 12273
rect 9103 12261 9112 12295
rect 9151 12261 9162 12295
rect 9313 12293 9347 12475
rect 9473 12661 9807 12703
rect 9473 12627 9491 12661
rect 9525 12627 9755 12661
rect 9789 12627 9807 12661
rect 9473 12559 9807 12627
rect 9473 12525 9491 12559
rect 9525 12525 9755 12559
rect 9789 12525 9807 12559
rect 9473 12485 9807 12525
rect 9841 12632 9899 12703
rect 9841 12598 9853 12632
rect 9887 12598 9899 12632
rect 9841 12539 9899 12598
rect 9841 12505 9853 12539
rect 9887 12505 9899 12539
rect 9944 12647 10001 12703
rect 9944 12613 9959 12647
rect 9993 12613 10001 12647
rect 9944 12579 10001 12613
rect 9944 12545 9959 12579
rect 9993 12545 10001 12579
rect 9944 12529 10001 12545
rect 10035 12653 10087 12669
rect 10035 12619 10045 12653
rect 10079 12619 10087 12653
rect 10035 12585 10087 12619
rect 10122 12661 10173 12703
rect 10122 12627 10131 12661
rect 10165 12627 10173 12661
rect 10122 12611 10173 12627
rect 10207 12635 10259 12669
rect 10207 12626 10221 12635
rect 10035 12551 10045 12585
rect 10079 12577 10087 12585
rect 10207 12592 10217 12626
rect 10255 12601 10259 12635
rect 10251 12592 10259 12601
rect 10207 12577 10259 12592
rect 10079 12551 10259 12577
rect 10035 12543 10259 12551
rect 10293 12661 10355 12703
rect 10293 12627 10313 12661
rect 10347 12627 10355 12661
rect 10293 12593 10355 12627
rect 10293 12559 10313 12593
rect 10347 12559 10355 12593
rect 10293 12543 10355 12559
rect 10389 12653 10451 12669
rect 10389 12619 10399 12653
rect 10433 12619 10451 12653
rect 9473 12415 9623 12485
rect 9841 12470 9899 12505
rect 10035 12517 10087 12543
rect 10035 12493 10045 12517
rect 9936 12483 10045 12493
rect 10079 12483 10087 12517
rect 10389 12531 10451 12619
rect 10389 12509 10399 12531
rect 9936 12459 10087 12483
rect 10245 12497 10399 12509
rect 10433 12497 10451 12531
rect 10245 12475 10451 12497
rect 9473 12381 9493 12415
rect 9527 12381 9623 12415
rect 9657 12417 9753 12451
rect 9787 12417 9807 12451
rect 9657 12347 9807 12417
rect 9103 12245 9162 12261
rect 9198 12273 9253 12289
rect 9018 12193 9069 12239
rect 9198 12239 9209 12273
rect 9243 12239 9253 12273
rect 9198 12193 9253 12239
rect 9287 12277 9347 12293
rect 9287 12243 9295 12277
rect 9329 12243 9347 12277
rect 9287 12227 9347 12243
rect 9473 12295 9807 12347
rect 9936 12357 10017 12459
rect 10245 12425 10279 12475
rect 10051 12391 10067 12425
rect 10101 12391 10135 12425
rect 10169 12391 10203 12425
rect 10237 12391 10279 12425
rect 10313 12425 10383 12441
rect 10313 12391 10349 12425
rect 10313 12363 10383 12391
rect 9473 12261 9491 12295
rect 9525 12261 9755 12295
rect 9789 12261 9807 12295
rect 9473 12193 9807 12261
rect 9841 12321 9899 12338
rect 9936 12323 10266 12357
rect 10347 12329 10383 12363
rect 10313 12327 10383 12329
rect 9841 12287 9853 12321
rect 9887 12287 9899 12321
rect 10035 12295 10087 12323
rect 9841 12193 9899 12287
rect 9945 12273 10001 12289
rect 9945 12239 9958 12273
rect 9992 12239 10001 12273
rect 10035 12261 10044 12295
rect 10078 12261 10087 12295
rect 10207 12295 10266 12323
rect 10035 12245 10087 12261
rect 10122 12273 10173 12289
rect 9945 12193 10001 12239
rect 10122 12239 10130 12273
rect 10164 12239 10173 12273
rect 10207 12261 10216 12295
rect 10250 12261 10266 12295
rect 10417 12293 10451 12475
rect 10207 12245 10266 12261
rect 10302 12273 10357 12289
rect 10122 12193 10173 12239
rect 10302 12239 10313 12273
rect 10347 12239 10357 12273
rect 10302 12193 10357 12239
rect 10391 12277 10451 12293
rect 10391 12243 10399 12277
rect 10433 12243 10451 12277
rect 10391 12227 10451 12243
rect 10486 12661 10553 12669
rect 10486 12627 10503 12661
rect 10537 12627 10553 12661
rect 10486 12593 10553 12627
rect 10486 12567 10503 12593
rect 10486 12533 10497 12567
rect 10537 12559 10553 12593
rect 10531 12533 10553 12559
rect 10486 12525 10553 12533
rect 10486 12491 10503 12525
rect 10537 12491 10553 12525
rect 10486 12475 10553 12491
rect 10587 12661 10621 12703
rect 10587 12593 10621 12627
rect 10587 12525 10621 12559
rect 10587 12475 10621 12491
rect 10655 12635 11061 12669
rect 10486 12341 10520 12475
rect 10655 12441 10689 12635
rect 10554 12425 10605 12441
rect 10588 12391 10605 12425
rect 10554 12375 10605 12391
rect 10650 12425 10689 12441
rect 10684 12391 10689 12425
rect 10650 12375 10689 12391
rect 10723 12567 10823 12601
rect 10857 12567 10898 12601
rect 10932 12567 10948 12601
rect 10571 12341 10605 12375
rect 10723 12341 10757 12567
rect 10486 12288 10537 12341
rect 10571 12307 10757 12341
rect 10791 12502 10993 12533
rect 10791 12499 10959 12502
rect 10791 12389 10825 12499
rect 10955 12465 10957 12499
rect 10991 12465 10993 12468
rect 10866 12431 10921 12459
rect 10899 12397 10921 12431
rect 10791 12339 10825 12355
rect 10866 12389 10921 12397
rect 10866 12355 10887 12389
rect 10486 12254 10503 12288
rect 10722 12300 10757 12307
rect 10722 12284 10828 12300
rect 10486 12227 10537 12254
rect 10571 12269 10637 12273
rect 10571 12235 10587 12269
rect 10621 12235 10637 12269
rect 10571 12193 10637 12235
rect 10722 12250 10794 12284
rect 10722 12227 10828 12250
rect 10866 12227 10921 12355
rect 10955 12227 10993 12465
rect 11027 12502 11061 12635
rect 11095 12601 11129 12703
rect 11095 12551 11129 12567
rect 11176 12601 11279 12633
rect 11176 12567 11181 12601
rect 11215 12567 11279 12601
rect 11176 12551 11279 12567
rect 11027 12468 11127 12502
rect 11161 12499 11177 12502
rect 11027 12465 11141 12468
rect 11175 12465 11177 12499
rect 11027 12464 11177 12465
rect 11211 12389 11279 12551
rect 11033 12355 11049 12389
rect 11083 12355 11279 12389
rect 11405 12601 11508 12633
rect 11405 12567 11469 12601
rect 11503 12567 11508 12601
rect 11405 12551 11508 12567
rect 11555 12601 11589 12703
rect 11555 12551 11589 12567
rect 11623 12635 12029 12669
rect 11405 12389 11473 12551
rect 11623 12502 11657 12635
rect 11736 12567 11752 12601
rect 11786 12567 11827 12601
rect 11861 12567 11961 12601
rect 11507 12468 11523 12502
rect 11557 12499 11657 12502
rect 11557 12468 11601 12499
rect 11507 12465 11601 12468
rect 11635 12465 11657 12499
rect 11507 12464 11657 12465
rect 11691 12502 11893 12533
rect 11725 12499 11893 12502
rect 11725 12468 11729 12499
rect 11405 12355 11601 12389
rect 11635 12355 11651 12389
rect 11029 12284 11131 12300
rect 11063 12250 11097 12284
rect 11029 12193 11131 12250
rect 11175 12284 11224 12355
rect 11175 12250 11181 12284
rect 11215 12250 11224 12284
rect 11175 12234 11224 12250
rect 11460 12284 11509 12355
rect 11460 12250 11469 12284
rect 11503 12250 11509 12284
rect 11460 12234 11509 12250
rect 11553 12284 11655 12300
rect 11587 12250 11621 12284
rect 11553 12193 11655 12250
rect 11691 12295 11729 12468
rect 11691 12261 11693 12295
rect 11727 12261 11729 12295
rect 11691 12227 11729 12261
rect 11763 12431 11818 12459
rect 11763 12397 11785 12431
rect 11763 12389 11818 12397
rect 11797 12355 11818 12389
rect 11763 12227 11818 12355
rect 11859 12389 11893 12499
rect 11859 12339 11893 12355
rect 11927 12341 11961 12567
rect 11995 12441 12029 12635
rect 12063 12661 12097 12703
rect 12063 12593 12097 12627
rect 12063 12525 12097 12559
rect 12063 12475 12097 12491
rect 12131 12661 12198 12669
rect 12131 12627 12147 12661
rect 12181 12635 12198 12661
rect 12131 12601 12153 12627
rect 12187 12601 12198 12635
rect 12131 12593 12198 12601
rect 12131 12559 12147 12593
rect 12181 12559 12198 12593
rect 12131 12525 12198 12559
rect 12131 12491 12147 12525
rect 12181 12491 12198 12525
rect 12131 12475 12198 12491
rect 11995 12425 12034 12441
rect 11995 12391 12000 12425
rect 11995 12375 12034 12391
rect 12079 12425 12130 12441
rect 12079 12391 12096 12425
rect 12079 12375 12130 12391
rect 12079 12341 12113 12375
rect 12164 12341 12198 12475
rect 12417 12632 12475 12703
rect 12417 12598 12429 12632
rect 12463 12598 12475 12632
rect 12417 12539 12475 12598
rect 12417 12505 12429 12539
rect 12463 12505 12475 12539
rect 12704 12647 12761 12703
rect 12704 12613 12719 12647
rect 12753 12613 12761 12647
rect 12704 12579 12761 12613
rect 12704 12545 12719 12579
rect 12753 12545 12761 12579
rect 12704 12529 12761 12545
rect 12795 12653 12847 12669
rect 12795 12619 12805 12653
rect 12839 12619 12847 12653
rect 12795 12585 12847 12619
rect 12882 12661 12933 12703
rect 12882 12627 12891 12661
rect 12925 12627 12933 12661
rect 12882 12611 12933 12627
rect 12967 12626 13019 12669
rect 12795 12551 12805 12585
rect 12839 12577 12847 12585
rect 12967 12592 12977 12626
rect 13011 12592 13019 12626
rect 12967 12577 13019 12592
rect 12839 12551 13019 12577
rect 12795 12543 13019 12551
rect 13053 12661 13115 12703
rect 13053 12627 13073 12661
rect 13107 12627 13115 12661
rect 13053 12593 13115 12627
rect 13053 12559 13073 12593
rect 13107 12559 13115 12593
rect 13053 12543 13115 12559
rect 13149 12653 13211 12669
rect 13149 12619 13159 12653
rect 13193 12619 13211 12653
rect 12417 12470 12475 12505
rect 12795 12517 12847 12543
rect 12795 12493 12805 12517
rect 12696 12483 12805 12493
rect 12839 12483 12847 12517
rect 13149 12531 13211 12619
rect 13149 12509 13159 12531
rect 11927 12307 12113 12341
rect 11927 12300 11962 12307
rect 11856 12284 11962 12300
rect 11890 12250 11962 12284
rect 12147 12288 12198 12341
rect 12696 12459 12847 12483
rect 13005 12497 13159 12509
rect 13193 12497 13211 12531
rect 13005 12475 13211 12497
rect 12696 12357 12777 12459
rect 13005 12425 13039 12475
rect 12811 12391 12827 12425
rect 12861 12391 12895 12425
rect 12929 12391 12963 12425
rect 12997 12391 13039 12425
rect 13073 12431 13143 12441
rect 13107 12425 13143 12431
rect 13107 12397 13109 12425
rect 13073 12391 13109 12397
rect 11856 12227 11962 12250
rect 12047 12269 12113 12273
rect 12047 12235 12063 12269
rect 12097 12235 12113 12269
rect 12047 12193 12113 12235
rect 12181 12254 12198 12288
rect 12147 12227 12198 12254
rect 12417 12321 12475 12338
rect 12696 12323 13026 12357
rect 13073 12327 13143 12391
rect 12417 12287 12429 12321
rect 12463 12287 12475 12321
rect 12795 12295 12847 12323
rect 12417 12193 12475 12287
rect 12705 12273 12761 12289
rect 12705 12239 12718 12273
rect 12752 12239 12761 12273
rect 12795 12261 12804 12295
rect 12838 12261 12847 12295
rect 12967 12295 13026 12323
rect 12795 12245 12847 12261
rect 12882 12273 12933 12289
rect 12705 12193 12761 12239
rect 12882 12239 12890 12273
rect 12924 12239 12933 12273
rect 12967 12261 12976 12295
rect 13015 12261 13026 12295
rect 13177 12293 13211 12475
rect 12967 12245 13026 12261
rect 13062 12273 13117 12289
rect 12882 12193 12933 12239
rect 13062 12239 13073 12273
rect 13107 12239 13117 12273
rect 13062 12193 13117 12239
rect 13151 12277 13211 12293
rect 13151 12243 13159 12277
rect 13193 12243 13211 12277
rect 13151 12227 13211 12243
rect 13245 12653 13307 12669
rect 13245 12619 13263 12653
rect 13297 12619 13307 12653
rect 13245 12531 13307 12619
rect 13341 12661 13403 12703
rect 13341 12627 13349 12661
rect 13383 12627 13403 12661
rect 13341 12593 13403 12627
rect 13341 12559 13349 12593
rect 13383 12559 13403 12593
rect 13341 12543 13403 12559
rect 13437 12626 13489 12669
rect 13437 12592 13445 12626
rect 13479 12592 13489 12626
rect 13523 12661 13574 12703
rect 13523 12627 13531 12661
rect 13565 12627 13574 12661
rect 13523 12611 13574 12627
rect 13609 12653 13661 12669
rect 13609 12619 13617 12653
rect 13651 12619 13661 12653
rect 13437 12577 13489 12592
rect 13609 12585 13661 12619
rect 13609 12577 13617 12585
rect 13437 12551 13617 12577
rect 13651 12551 13661 12585
rect 13437 12543 13661 12551
rect 13245 12497 13263 12531
rect 13297 12509 13307 12531
rect 13609 12517 13661 12543
rect 13695 12647 13752 12703
rect 13695 12613 13703 12647
rect 13737 12613 13752 12647
rect 13695 12579 13752 12613
rect 13695 12545 13703 12579
rect 13737 12545 13752 12579
rect 13695 12529 13752 12545
rect 13815 12653 13849 12669
rect 13815 12585 13849 12619
rect 13885 12653 13951 12703
rect 13885 12619 13901 12653
rect 13935 12619 13951 12653
rect 13885 12585 13951 12619
rect 13885 12551 13901 12585
rect 13935 12551 13951 12585
rect 13985 12653 14039 12669
rect 13985 12619 13987 12653
rect 14021 12635 14039 12653
rect 13985 12601 13993 12619
rect 14027 12601 14039 12635
rect 13985 12572 14039 12601
rect 13297 12497 13451 12509
rect 13245 12475 13451 12497
rect 13245 12293 13279 12475
rect 13313 12431 13383 12441
rect 13313 12425 13349 12431
rect 13347 12397 13349 12425
rect 13347 12391 13383 12397
rect 13417 12425 13451 12475
rect 13609 12483 13617 12517
rect 13651 12493 13661 12517
rect 13815 12517 13849 12551
rect 13985 12538 13987 12572
rect 14021 12538 14039 12572
rect 13651 12483 13760 12493
rect 13815 12483 13948 12517
rect 13985 12488 14039 12538
rect 14096 12635 14153 12669
rect 14096 12601 14113 12635
rect 14147 12601 14153 12635
rect 14187 12661 14241 12703
rect 14187 12627 14197 12661
rect 14231 12627 14241 12661
rect 14187 12611 14241 12627
rect 14321 12635 14401 12669
rect 14096 12577 14153 12601
rect 14321 12601 14351 12635
rect 14385 12601 14401 12635
rect 14096 12533 14287 12577
rect 13609 12459 13760 12483
rect 13417 12391 13459 12425
rect 13493 12391 13527 12425
rect 13561 12391 13595 12425
rect 13629 12391 13645 12425
rect 13313 12327 13383 12391
rect 13679 12357 13760 12459
rect 13914 12454 13948 12483
rect 13801 12431 13867 12447
rect 13801 12397 13809 12431
rect 13843 12425 13867 12431
rect 13801 12391 13817 12397
rect 13851 12391 13867 12425
rect 13801 12373 13867 12391
rect 13914 12438 13971 12454
rect 13914 12404 13937 12438
rect 13914 12388 13971 12404
rect 13430 12323 13760 12357
rect 13914 12337 13948 12388
rect 13430 12295 13489 12323
rect 13245 12277 13305 12293
rect 13245 12243 13263 12277
rect 13297 12243 13305 12277
rect 13245 12227 13305 12243
rect 13339 12273 13394 12289
rect 13339 12239 13349 12273
rect 13383 12239 13394 12273
rect 13430 12261 13446 12295
rect 13480 12261 13489 12295
rect 13609 12295 13661 12323
rect 13430 12245 13489 12261
rect 13523 12273 13574 12289
rect 13339 12193 13394 12239
rect 13523 12239 13532 12273
rect 13566 12239 13574 12273
rect 13609 12261 13618 12295
rect 13659 12261 13661 12295
rect 13815 12303 13948 12337
rect 14005 12328 14039 12488
rect 14073 12465 14177 12499
rect 14073 12425 14211 12465
rect 14073 12391 14137 12425
rect 14171 12391 14211 12425
rect 14073 12387 14211 12391
rect 14245 12425 14287 12533
rect 14245 12391 14251 12425
rect 14285 12391 14287 12425
rect 14245 12353 14287 12391
rect 13609 12245 13661 12261
rect 13695 12273 13751 12289
rect 13523 12193 13574 12239
rect 13695 12239 13704 12273
rect 13738 12239 13751 12273
rect 13695 12193 13751 12239
rect 13815 12282 13849 12303
rect 13987 12299 14039 12328
rect 13815 12227 13849 12248
rect 13885 12235 13901 12269
rect 13935 12235 13951 12269
rect 13885 12193 13951 12235
rect 14021 12265 14039 12299
rect 13987 12227 14039 12265
rect 14096 12319 14287 12353
rect 14321 12499 14401 12601
rect 14439 12635 14495 12669
rect 14439 12601 14455 12635
rect 14489 12601 14495 12635
rect 14599 12661 14664 12703
rect 14599 12627 14614 12661
rect 14648 12627 14664 12661
rect 14599 12611 14664 12627
rect 14698 12635 14775 12669
rect 14439 12577 14495 12601
rect 14698 12601 14704 12635
rect 14763 12601 14775 12635
rect 14439 12533 14664 12577
rect 14321 12425 14540 12499
rect 14321 12391 14455 12425
rect 14489 12391 14540 12425
rect 14321 12387 14540 12391
rect 14574 12441 14664 12533
rect 14698 12475 14775 12601
rect 14574 12425 14685 12441
rect 14574 12391 14651 12425
rect 14096 12295 14153 12319
rect 14096 12261 14113 12295
rect 14147 12261 14153 12295
rect 14321 12295 14401 12387
rect 14574 12375 14685 12391
rect 14574 12353 14664 12375
rect 14096 12227 14153 12261
rect 14187 12269 14241 12285
rect 14187 12235 14197 12269
rect 14231 12235 14241 12269
rect 14187 12193 14241 12235
rect 14321 12261 14351 12295
rect 14385 12261 14401 12295
rect 14321 12227 14401 12261
rect 14439 12319 14664 12353
rect 14719 12341 14775 12475
rect 14993 12632 15051 12703
rect 14993 12598 15005 12632
rect 15039 12598 15051 12632
rect 14993 12539 15051 12598
rect 14993 12505 15005 12539
rect 15039 12505 15051 12539
rect 15086 12653 15137 12669
rect 15086 12619 15103 12653
rect 15086 12585 15137 12619
rect 15171 12637 15237 12703
rect 15171 12603 15187 12637
rect 15221 12603 15237 12637
rect 15271 12653 15305 12669
rect 15086 12551 15103 12585
rect 15271 12585 15305 12619
rect 15137 12551 15236 12569
rect 15086 12535 15236 12551
rect 14993 12470 15051 12505
rect 15086 12499 15156 12501
rect 15086 12465 15097 12499
rect 15131 12465 15156 12499
rect 15086 12425 15156 12465
rect 15086 12391 15100 12425
rect 15134 12391 15156 12425
rect 15086 12371 15156 12391
rect 15190 12440 15236 12535
rect 15190 12431 15202 12440
rect 15224 12397 15236 12406
rect 14439 12295 14495 12319
rect 14439 12261 14455 12295
rect 14489 12261 14495 12295
rect 14698 12295 14775 12341
rect 14439 12227 14495 12261
rect 14599 12269 14664 12285
rect 14599 12235 14614 12269
rect 14648 12235 14664 12269
rect 14599 12193 14664 12235
rect 14698 12261 14704 12295
rect 14738 12261 14775 12295
rect 14698 12227 14775 12261
rect 14993 12321 15051 12338
rect 15190 12337 15236 12397
rect 14993 12287 15005 12321
rect 15039 12287 15051 12321
rect 14993 12193 15051 12287
rect 15086 12303 15236 12337
rect 15086 12295 15137 12303
rect 15086 12261 15103 12295
rect 15271 12295 15305 12533
rect 15339 12509 15404 12666
rect 15438 12661 15488 12703
rect 15438 12627 15454 12661
rect 15438 12611 15488 12627
rect 15522 12653 15572 12669
rect 15522 12619 15538 12653
rect 15522 12603 15572 12619
rect 15615 12659 15751 12669
rect 15615 12625 15631 12659
rect 15665 12625 15751 12659
rect 15866 12651 15932 12703
rect 16059 12661 16133 12703
rect 15615 12603 15751 12625
rect 15522 12577 15556 12603
rect 15477 12543 15556 12577
rect 15590 12567 15683 12569
rect 15351 12499 15443 12509
rect 15351 12465 15373 12499
rect 15407 12486 15443 12499
rect 15407 12465 15409 12486
rect 15351 12452 15409 12465
rect 15351 12299 15443 12452
rect 15086 12245 15137 12261
rect 15171 12235 15187 12269
rect 15221 12235 15237 12269
rect 15477 12271 15511 12543
rect 15590 12541 15649 12567
rect 15624 12533 15649 12541
rect 15624 12507 15683 12533
rect 15590 12491 15683 12507
rect 15545 12431 15615 12453
rect 15545 12397 15557 12431
rect 15591 12397 15615 12431
rect 15545 12379 15615 12397
rect 15545 12345 15568 12379
rect 15602 12345 15615 12379
rect 15545 12329 15615 12345
rect 15649 12373 15683 12491
rect 15717 12447 15751 12603
rect 15785 12635 15819 12651
rect 15866 12617 15882 12651
rect 15916 12617 15932 12651
rect 15966 12635 16000 12651
rect 15785 12583 15819 12601
rect 16059 12627 16079 12661
rect 16113 12627 16133 12661
rect 16059 12611 16133 12627
rect 16167 12653 16201 12669
rect 15966 12583 16000 12601
rect 15785 12549 16000 12583
rect 16167 12577 16201 12619
rect 16248 12660 16422 12669
rect 16248 12626 16264 12660
rect 16298 12626 16422 12660
rect 16248 12601 16422 12626
rect 16456 12661 16506 12703
rect 16490 12627 16506 12661
rect 16610 12661 16676 12703
rect 16456 12611 16506 12627
rect 16540 12635 16574 12651
rect 16089 12543 16201 12577
rect 16089 12515 16123 12543
rect 15823 12481 15839 12515
rect 15873 12481 16123 12515
rect 16262 12533 16273 12567
rect 16307 12541 16354 12567
rect 16262 12509 16304 12533
rect 15717 12427 16055 12447
rect 15717 12413 16021 12427
rect 15649 12339 15670 12373
rect 15704 12339 15720 12373
rect 15649 12329 15720 12339
rect 15754 12271 15788 12413
rect 15829 12363 15925 12379
rect 15863 12329 15901 12363
rect 15959 12345 15987 12379
rect 16021 12377 16055 12393
rect 15935 12329 15987 12345
rect 16089 12343 16123 12481
rect 15271 12245 15305 12261
rect 15171 12193 15237 12235
rect 15377 12231 15393 12265
rect 15427 12231 15443 12265
rect 15477 12237 15526 12271
rect 15560 12237 15576 12271
rect 15617 12237 15633 12271
rect 15667 12237 15788 12271
rect 15963 12269 16029 12285
rect 15377 12193 15443 12231
rect 15963 12235 15979 12269
rect 16013 12235 16029 12269
rect 15963 12193 16029 12235
rect 16071 12265 16123 12343
rect 16161 12507 16304 12509
rect 16338 12507 16354 12541
rect 16388 12525 16422 12601
rect 16610 12627 16626 12661
rect 16660 12627 16676 12661
rect 16744 12661 16805 12703
rect 16744 12627 16755 12661
rect 16789 12627 16805 12661
rect 17017 12653 17079 12669
rect 16540 12593 16574 12601
rect 16744 12593 16805 12627
rect 16540 12559 16700 12593
rect 16161 12475 16296 12507
rect 16388 12491 16582 12525
rect 16616 12491 16632 12525
rect 16161 12367 16203 12475
rect 16388 12473 16422 12491
rect 16161 12333 16169 12367
rect 16161 12317 16203 12333
rect 16237 12431 16307 12441
rect 16237 12415 16273 12431
rect 16237 12381 16265 12415
rect 16299 12381 16307 12397
rect 16237 12317 16307 12381
rect 16341 12439 16422 12473
rect 16341 12283 16375 12439
rect 16489 12426 16597 12457
rect 16666 12441 16700 12559
rect 16744 12559 16755 12593
rect 16789 12559 16805 12593
rect 16744 12475 16805 12559
rect 16839 12625 16890 12641
rect 16873 12591 16890 12625
rect 16839 12557 16890 12591
rect 16873 12523 16890 12557
rect 16839 12499 16890 12523
rect 16839 12465 16845 12499
rect 16879 12465 16890 12499
rect 16666 12435 16814 12441
rect 16523 12417 16597 12426
rect 16409 12389 16453 12405
rect 16443 12355 16453 12389
rect 16489 12383 16505 12392
rect 16539 12383 16597 12417
rect 16409 12349 16453 12355
rect 16549 12363 16597 12383
rect 16409 12315 16515 12349
rect 16185 12269 16375 12283
rect 16071 12231 16091 12265
rect 16125 12231 16141 12265
rect 16185 12235 16201 12269
rect 16235 12235 16375 12269
rect 16185 12227 16375 12235
rect 16409 12265 16447 12281
rect 16409 12231 16413 12265
rect 16481 12269 16515 12315
rect 16583 12329 16597 12363
rect 16549 12303 16597 12329
rect 16631 12425 16814 12435
rect 16631 12391 16780 12425
rect 16631 12375 16814 12391
rect 16631 12340 16696 12375
rect 16631 12285 16695 12340
rect 16848 12335 16890 12465
rect 16839 12319 16890 12335
rect 16873 12285 16890 12319
rect 16481 12251 16631 12269
rect 16665 12251 16695 12285
rect 16481 12235 16695 12251
rect 16744 12269 16805 12285
rect 16744 12235 16755 12269
rect 16789 12235 16805 12269
rect 16409 12193 16447 12231
rect 16744 12193 16805 12235
rect 16839 12229 16890 12285
rect 17017 12619 17035 12653
rect 17069 12619 17079 12653
rect 17017 12531 17079 12619
rect 17113 12661 17175 12703
rect 17113 12627 17121 12661
rect 17155 12627 17175 12661
rect 17113 12593 17175 12627
rect 17113 12559 17121 12593
rect 17155 12559 17175 12593
rect 17113 12543 17175 12559
rect 17209 12626 17261 12669
rect 17209 12592 17217 12626
rect 17251 12592 17261 12626
rect 17295 12661 17346 12703
rect 17295 12627 17303 12661
rect 17337 12627 17346 12661
rect 17295 12611 17346 12627
rect 17381 12653 17433 12669
rect 17381 12619 17389 12653
rect 17423 12619 17433 12653
rect 17209 12577 17261 12592
rect 17381 12585 17433 12619
rect 17381 12577 17389 12585
rect 17209 12551 17389 12577
rect 17423 12551 17433 12585
rect 17209 12543 17433 12551
rect 17017 12497 17035 12531
rect 17069 12509 17079 12531
rect 17381 12517 17433 12543
rect 17467 12647 17524 12703
rect 17467 12613 17475 12647
rect 17509 12613 17524 12647
rect 17467 12579 17524 12613
rect 17467 12545 17475 12579
rect 17509 12545 17524 12579
rect 17467 12529 17524 12545
rect 17569 12632 17627 12703
rect 17569 12598 17581 12632
rect 17615 12598 17627 12632
rect 17569 12539 17627 12598
rect 17069 12497 17223 12509
rect 17017 12475 17223 12497
rect 17017 12293 17051 12475
rect 17085 12431 17155 12441
rect 17085 12425 17121 12431
rect 17119 12397 17121 12425
rect 17119 12391 17155 12397
rect 17189 12425 17223 12475
rect 17381 12483 17389 12517
rect 17423 12493 17433 12517
rect 17569 12505 17581 12539
rect 17615 12505 17627 12539
rect 17423 12483 17532 12493
rect 17381 12459 17532 12483
rect 17569 12470 17627 12505
rect 17753 12661 18271 12703
rect 17753 12627 17771 12661
rect 17805 12627 18219 12661
rect 18253 12627 18271 12661
rect 17753 12559 18271 12627
rect 18306 12661 19375 12703
rect 18306 12627 18323 12661
rect 18357 12627 19323 12661
rect 19357 12627 19375 12661
rect 18306 12616 19375 12627
rect 19409 12653 19471 12669
rect 19409 12619 19427 12653
rect 19461 12619 19471 12653
rect 17753 12525 17771 12559
rect 17805 12525 18219 12559
rect 18253 12525 18271 12559
rect 17753 12485 18271 12525
rect 17189 12391 17231 12425
rect 17265 12391 17299 12425
rect 17333 12391 17367 12425
rect 17401 12391 17417 12425
rect 17085 12327 17155 12391
rect 17451 12363 17532 12459
rect 17753 12415 17995 12485
rect 17753 12381 17831 12415
rect 17865 12381 17941 12415
rect 17975 12381 17995 12415
rect 18029 12417 18049 12451
rect 18083 12417 18159 12451
rect 18193 12417 18271 12451
rect 17451 12357 17489 12363
rect 17202 12329 17489 12357
rect 17523 12329 17532 12363
rect 18029 12347 18271 12417
rect 18624 12415 18694 12616
rect 19409 12531 19471 12619
rect 19505 12661 19567 12703
rect 19505 12627 19513 12661
rect 19547 12627 19567 12661
rect 19505 12593 19567 12627
rect 19505 12559 19513 12593
rect 19547 12559 19567 12593
rect 19505 12543 19567 12559
rect 19601 12626 19653 12669
rect 19601 12592 19609 12626
rect 19643 12592 19653 12626
rect 19687 12661 19738 12703
rect 19687 12627 19695 12661
rect 19729 12627 19738 12661
rect 19687 12611 19738 12627
rect 19773 12653 19825 12669
rect 19773 12619 19781 12653
rect 19815 12619 19825 12653
rect 19601 12577 19653 12592
rect 19773 12585 19825 12619
rect 19773 12577 19781 12585
rect 19601 12551 19781 12577
rect 19815 12551 19825 12585
rect 19601 12543 19825 12551
rect 19409 12497 19427 12531
rect 19461 12509 19471 12531
rect 19773 12517 19825 12543
rect 19859 12647 19916 12703
rect 19859 12613 19867 12647
rect 19901 12613 19916 12647
rect 19859 12579 19916 12613
rect 19859 12545 19867 12579
rect 19901 12545 19916 12579
rect 19859 12529 19916 12545
rect 19961 12661 20203 12703
rect 19961 12627 19979 12661
rect 20013 12627 20151 12661
rect 20185 12627 20203 12661
rect 19961 12566 20203 12627
rect 19961 12532 19979 12566
rect 20013 12532 20151 12566
rect 20185 12532 20203 12566
rect 19461 12497 19615 12509
rect 19409 12475 19615 12497
rect 18624 12381 18643 12415
rect 18677 12381 18694 12415
rect 18624 12366 18694 12381
rect 18990 12451 19058 12468
rect 18990 12417 19007 12451
rect 19041 12417 19058 12451
rect 17202 12323 17532 12329
rect 17202 12295 17261 12323
rect 17017 12277 17077 12293
rect 17017 12243 17035 12277
rect 17069 12243 17077 12277
rect 17017 12227 17077 12243
rect 17111 12273 17166 12289
rect 17111 12239 17121 12273
rect 17155 12239 17166 12273
rect 17202 12261 17218 12295
rect 17252 12261 17261 12295
rect 17381 12295 17433 12323
rect 17202 12245 17261 12261
rect 17295 12273 17346 12289
rect 17111 12193 17166 12239
rect 17295 12239 17304 12273
rect 17338 12239 17346 12273
rect 17381 12261 17390 12295
rect 17424 12261 17433 12295
rect 17569 12321 17627 12338
rect 17381 12245 17433 12261
rect 17467 12273 17523 12289
rect 17295 12193 17346 12239
rect 17467 12239 17476 12273
rect 17510 12239 17523 12273
rect 17467 12193 17523 12239
rect 17569 12287 17581 12321
rect 17615 12287 17627 12321
rect 17569 12193 17627 12287
rect 17753 12288 18271 12347
rect 18990 12302 19058 12417
rect 17753 12254 17771 12288
rect 17805 12254 18219 12288
rect 18253 12254 18271 12288
rect 17753 12193 18271 12254
rect 18306 12288 19375 12302
rect 18306 12254 18323 12288
rect 18357 12254 19323 12288
rect 19357 12254 19375 12288
rect 18306 12193 19375 12254
rect 19409 12293 19443 12475
rect 19477 12431 19547 12441
rect 19477 12425 19513 12431
rect 19511 12397 19513 12425
rect 19511 12391 19547 12397
rect 19581 12425 19615 12475
rect 19773 12483 19781 12517
rect 19815 12493 19825 12517
rect 19815 12483 19924 12493
rect 19773 12459 19924 12483
rect 19581 12391 19623 12425
rect 19657 12391 19691 12425
rect 19725 12391 19759 12425
rect 19793 12391 19809 12425
rect 19477 12327 19547 12391
rect 19843 12363 19924 12459
rect 19961 12485 20203 12532
rect 19961 12411 20065 12485
rect 19961 12377 20011 12411
rect 20045 12377 20065 12411
rect 20099 12417 20119 12451
rect 20153 12417 20203 12451
rect 19843 12357 19881 12363
rect 19594 12329 19881 12357
rect 19915 12329 19924 12363
rect 20099 12343 20203 12417
rect 19594 12323 19924 12329
rect 19594 12295 19653 12323
rect 19409 12277 19469 12293
rect 19409 12243 19427 12277
rect 19461 12243 19469 12277
rect 19409 12227 19469 12243
rect 19503 12273 19558 12289
rect 19503 12239 19513 12273
rect 19547 12239 19558 12273
rect 19594 12261 19610 12295
rect 19644 12261 19653 12295
rect 19773 12295 19825 12323
rect 19594 12245 19653 12261
rect 19687 12273 19738 12289
rect 19503 12193 19558 12239
rect 19687 12239 19696 12273
rect 19730 12239 19738 12273
rect 19773 12261 19782 12295
rect 19816 12261 19825 12295
rect 19961 12290 20203 12343
rect 19773 12245 19825 12261
rect 19859 12273 19915 12289
rect 19687 12193 19738 12239
rect 19859 12239 19868 12273
rect 19902 12239 19915 12273
rect 19859 12193 19915 12239
rect 19961 12256 19979 12290
rect 20013 12256 20151 12290
rect 20185 12256 20203 12290
rect 19961 12193 20203 12256
rect 4948 12159 4977 12193
rect 5011 12159 5069 12193
rect 5103 12159 5161 12193
rect 5195 12159 5253 12193
rect 5287 12159 5345 12193
rect 5379 12159 5437 12193
rect 5471 12159 5529 12193
rect 5563 12159 5621 12193
rect 5655 12159 5713 12193
rect 5747 12159 5805 12193
rect 5839 12159 5897 12193
rect 5931 12159 5989 12193
rect 6023 12159 6081 12193
rect 6115 12159 6173 12193
rect 6207 12159 6265 12193
rect 6299 12159 6357 12193
rect 6391 12159 6449 12193
rect 6483 12159 6541 12193
rect 6575 12159 6633 12193
rect 6667 12159 6725 12193
rect 6759 12159 6817 12193
rect 6851 12159 6909 12193
rect 6943 12159 7001 12193
rect 7035 12159 7093 12193
rect 7127 12159 7185 12193
rect 7219 12159 7277 12193
rect 7311 12159 7369 12193
rect 7403 12159 7461 12193
rect 7495 12159 7553 12193
rect 7587 12159 7645 12193
rect 7679 12159 7737 12193
rect 7771 12159 7829 12193
rect 7863 12159 7921 12193
rect 7955 12159 8013 12193
rect 8047 12159 8105 12193
rect 8139 12159 8197 12193
rect 8231 12159 8289 12193
rect 8323 12159 8381 12193
rect 8415 12159 8473 12193
rect 8507 12159 8565 12193
rect 8599 12159 8657 12193
rect 8691 12159 8749 12193
rect 8783 12159 8841 12193
rect 8875 12159 8933 12193
rect 8967 12159 9025 12193
rect 9059 12159 9117 12193
rect 9151 12159 9209 12193
rect 9243 12159 9301 12193
rect 9335 12159 9393 12193
rect 9427 12159 9485 12193
rect 9519 12159 9577 12193
rect 9611 12159 9669 12193
rect 9703 12159 9761 12193
rect 9795 12159 9853 12193
rect 9887 12159 9945 12193
rect 9979 12159 10037 12193
rect 10071 12159 10129 12193
rect 10163 12159 10221 12193
rect 10255 12159 10313 12193
rect 10347 12159 10405 12193
rect 10439 12159 10497 12193
rect 10531 12159 10589 12193
rect 10623 12159 10681 12193
rect 10715 12159 10773 12193
rect 10807 12159 10865 12193
rect 10899 12159 10957 12193
rect 10991 12159 11049 12193
rect 11083 12159 11141 12193
rect 11175 12159 11233 12193
rect 11267 12159 11325 12193
rect 11359 12159 11417 12193
rect 11451 12159 11509 12193
rect 11543 12159 11601 12193
rect 11635 12159 11693 12193
rect 11727 12159 11785 12193
rect 11819 12159 11877 12193
rect 11911 12159 11969 12193
rect 12003 12159 12061 12193
rect 12095 12159 12153 12193
rect 12187 12159 12245 12193
rect 12279 12159 12337 12193
rect 12371 12159 12429 12193
rect 12463 12159 12521 12193
rect 12555 12159 12613 12193
rect 12647 12159 12705 12193
rect 12739 12159 12797 12193
rect 12831 12159 12889 12193
rect 12923 12159 12981 12193
rect 13015 12159 13073 12193
rect 13107 12159 13165 12193
rect 13199 12159 13257 12193
rect 13291 12159 13349 12193
rect 13383 12159 13441 12193
rect 13475 12159 13533 12193
rect 13567 12159 13625 12193
rect 13659 12159 13717 12193
rect 13751 12159 13809 12193
rect 13843 12159 13901 12193
rect 13935 12159 13993 12193
rect 14027 12159 14085 12193
rect 14119 12159 14177 12193
rect 14211 12159 14269 12193
rect 14303 12159 14361 12193
rect 14395 12159 14453 12193
rect 14487 12159 14545 12193
rect 14579 12159 14637 12193
rect 14671 12159 14729 12193
rect 14763 12159 14821 12193
rect 14855 12159 14913 12193
rect 14947 12159 15005 12193
rect 15039 12159 15097 12193
rect 15131 12159 15189 12193
rect 15223 12159 15281 12193
rect 15315 12159 15373 12193
rect 15407 12159 15465 12193
rect 15499 12159 15557 12193
rect 15591 12159 15649 12193
rect 15683 12159 15741 12193
rect 15775 12159 15833 12193
rect 15867 12159 15925 12193
rect 15959 12159 16017 12193
rect 16051 12159 16109 12193
rect 16143 12159 16201 12193
rect 16235 12159 16293 12193
rect 16327 12159 16385 12193
rect 16419 12159 16477 12193
rect 16511 12159 16569 12193
rect 16603 12159 16661 12193
rect 16695 12159 16753 12193
rect 16787 12159 16845 12193
rect 16879 12159 16937 12193
rect 16971 12159 17029 12193
rect 17063 12159 17121 12193
rect 17155 12159 17213 12193
rect 17247 12159 17305 12193
rect 17339 12159 17397 12193
rect 17431 12159 17489 12193
rect 17523 12159 17581 12193
rect 17615 12159 17673 12193
rect 17707 12159 17765 12193
rect 17799 12159 17857 12193
rect 17891 12159 17949 12193
rect 17983 12159 18041 12193
rect 18075 12159 18133 12193
rect 18167 12159 18225 12193
rect 18259 12159 18317 12193
rect 18351 12159 18409 12193
rect 18443 12159 18501 12193
rect 18535 12159 18593 12193
rect 18627 12159 18685 12193
rect 18719 12159 18777 12193
rect 18811 12159 18869 12193
rect 18903 12159 18961 12193
rect 18995 12159 19053 12193
rect 19087 12159 19145 12193
rect 19179 12159 19237 12193
rect 19271 12159 19329 12193
rect 19363 12159 19421 12193
rect 19455 12159 19513 12193
rect 19547 12159 19605 12193
rect 19639 12159 19697 12193
rect 19731 12159 19789 12193
rect 19823 12159 19881 12193
rect 19915 12159 19973 12193
rect 20007 12159 20065 12193
rect 20099 12159 20157 12193
rect 20191 12159 20220 12193
rect 25716 9190 25812 9224
rect 28176 9190 28272 9224
rect 25716 9128 25750 9190
rect 28238 9128 28272 9190
rect 25716 7050 25750 7112
rect 28238 7050 28272 7112
rect 25716 7016 25812 7050
rect 28176 7016 28272 7050
rect 29580 7050 34840 7070
rect 29580 7010 29680 7050
rect 34760 7010 34840 7050
rect 29580 6990 34840 7010
rect 16886 6850 16982 6884
rect 17120 6850 17216 6884
rect 16886 6788 16920 6850
rect 13286 6290 13382 6324
rect 13520 6290 13616 6324
rect 13286 6228 13320 6290
rect 9986 6010 10082 6044
rect 10220 6010 10316 6044
rect 3386 5966 3482 6000
rect 3620 5966 3716 6000
rect 3386 5904 3420 5966
rect 3682 5904 3716 5966
rect 9986 5948 10020 6010
rect 3386 4710 3420 4772
rect 3682 4710 3716 4772
rect 3386 4676 3482 4710
rect 3620 4676 3716 4710
rect 6686 5870 6782 5904
rect 6920 5870 7016 5904
rect 6686 5808 6720 5870
rect 6982 5808 7016 5870
rect 6686 4710 6720 4772
rect 6982 4710 7016 4772
rect 6686 4676 6782 4710
rect 6920 4676 7016 4710
rect 10282 5948 10316 6010
rect 9986 4710 10020 4772
rect 10282 4710 10316 4772
rect 9986 4676 10082 4710
rect 10220 4676 10316 4710
rect 13582 6228 13616 6290
rect 13286 4710 13320 4772
rect 13582 4710 13616 4772
rect 13286 4676 13382 4710
rect 13520 4676 13616 4710
rect 17182 6788 17216 6850
rect 16886 4710 16920 4772
rect 17182 4710 17216 4772
rect 16886 4676 16982 4710
rect 17120 4676 17216 4710
rect 20086 6850 20182 6884
rect 20638 6850 20734 6884
rect 20086 6788 20120 6850
rect 20700 6788 20734 6850
rect 20086 4710 20120 4772
rect 20700 4710 20734 4772
rect 20086 4676 20182 4710
rect 20638 4676 20734 4710
rect 23186 6850 23282 6884
rect 24374 6850 24470 6884
rect 23186 6788 23220 6850
rect 24436 6788 24470 6850
rect 23186 4710 23220 4772
rect 24436 4710 24470 4772
rect 23186 4676 23282 4710
rect 24374 4676 24470 4710
rect 25686 6850 25782 6884
rect 28146 6850 28242 6884
rect 25686 6788 25720 6850
rect 28208 6788 28242 6850
rect 25686 4710 25720 4772
rect 29580 4970 29600 6990
rect 29640 4990 29660 6990
rect 34760 6970 34840 6990
rect 29814 6797 29830 6831
rect 29998 6797 30014 6831
rect 30194 6797 30210 6831
rect 30378 6797 30394 6831
rect 30452 6797 30468 6831
rect 30636 6797 30652 6831
rect 30834 6797 30850 6831
rect 31018 6797 31034 6831
rect 31092 6797 31108 6831
rect 31276 6797 31292 6831
rect 31350 6797 31366 6831
rect 31534 6797 31550 6831
rect 31734 6797 31750 6831
rect 31918 6797 31934 6831
rect 31992 6797 32008 6831
rect 32176 6797 32192 6831
rect 32250 6797 32266 6831
rect 32434 6797 32450 6831
rect 32508 6797 32524 6831
rect 32692 6797 32708 6831
rect 32766 6797 32782 6831
rect 32950 6797 32966 6831
rect 33024 6797 33040 6831
rect 33208 6797 33224 6831
rect 33282 6797 33298 6831
rect 33466 6797 33482 6831
rect 33540 6797 33556 6831
rect 33724 6797 33740 6831
rect 33798 6797 33814 6831
rect 33982 6797 33998 6831
rect 34056 6797 34072 6831
rect 34240 6797 34256 6831
rect 34434 6797 34450 6831
rect 34618 6797 34634 6831
rect 29768 6738 29802 6754
rect 29768 6146 29802 6162
rect 30026 6738 30060 6754
rect 30026 6146 30060 6162
rect 30148 6738 30182 6754
rect 30148 6146 30182 6162
rect 30406 6738 30440 6754
rect 30406 6146 30440 6162
rect 30664 6738 30698 6754
rect 30664 6146 30698 6162
rect 30788 6738 30822 6754
rect 30788 6146 30822 6162
rect 31046 6738 31080 6754
rect 31046 6146 31080 6162
rect 31304 6738 31338 6754
rect 31304 6146 31338 6162
rect 31562 6738 31596 6754
rect 31562 6146 31596 6162
rect 31688 6738 31722 6754
rect 31688 6146 31722 6162
rect 31946 6738 31980 6754
rect 31946 6146 31980 6162
rect 32204 6738 32238 6754
rect 32204 6146 32238 6162
rect 32462 6738 32496 6754
rect 32462 6146 32496 6162
rect 32720 6738 32754 6754
rect 32720 6146 32754 6162
rect 32978 6738 33012 6754
rect 32978 6146 33012 6162
rect 33236 6738 33270 6754
rect 33236 6146 33270 6162
rect 33494 6738 33528 6754
rect 33494 6146 33528 6162
rect 33752 6738 33786 6754
rect 33752 6146 33786 6162
rect 34010 6738 34044 6754
rect 34010 6146 34044 6162
rect 34268 6738 34302 6754
rect 34268 6146 34302 6162
rect 34388 6738 34422 6754
rect 34388 6146 34422 6162
rect 34646 6738 34680 6754
rect 34646 6146 34680 6162
rect 29814 6069 29830 6103
rect 29998 6069 30014 6103
rect 30194 6069 30210 6103
rect 30378 6069 30394 6103
rect 30452 6069 30468 6103
rect 30636 6069 30652 6103
rect 30834 6069 30850 6103
rect 31018 6069 31034 6103
rect 31092 6069 31108 6103
rect 31276 6069 31292 6103
rect 31350 6069 31366 6103
rect 31534 6069 31550 6103
rect 31734 6069 31750 6103
rect 31918 6069 31934 6103
rect 31992 6069 32008 6103
rect 32176 6069 32192 6103
rect 32250 6069 32266 6103
rect 32434 6069 32450 6103
rect 32508 6069 32524 6103
rect 32692 6069 32708 6103
rect 32766 6069 32782 6103
rect 32950 6069 32966 6103
rect 33024 6069 33040 6103
rect 33208 6069 33224 6103
rect 33282 6069 33298 6103
rect 33466 6069 33482 6103
rect 33540 6069 33556 6103
rect 33724 6069 33740 6103
rect 33798 6069 33814 6103
rect 33982 6069 33998 6103
rect 34056 6069 34072 6103
rect 34240 6069 34256 6103
rect 34434 6069 34450 6103
rect 34618 6069 34634 6103
rect 30056 5777 30072 5811
rect 30106 5777 30122 5811
rect 30376 5777 30392 5811
rect 30426 5777 30442 5811
rect 30776 5777 30792 5811
rect 30826 5777 30842 5811
rect 31076 5777 31092 5811
rect 31126 5777 31142 5811
rect 30028 5718 30062 5734
rect 30028 5126 30062 5142
rect 30116 5718 30150 5734
rect 30116 5126 30150 5142
rect 30248 5718 30282 5734
rect 30248 5126 30282 5142
rect 30344 5718 30378 5734
rect 30344 5126 30378 5142
rect 30440 5718 30474 5734
rect 30440 5126 30474 5142
rect 30536 5718 30570 5734
rect 30536 5126 30570 5142
rect 30648 5718 30682 5734
rect 30648 5126 30682 5142
rect 30744 5718 30778 5734
rect 30744 5126 30778 5142
rect 30840 5718 30874 5734
rect 30840 5126 30874 5142
rect 30936 5718 30970 5734
rect 30936 5126 30970 5142
rect 31048 5718 31082 5734
rect 31048 5126 31082 5142
rect 31136 5718 31170 5734
rect 31136 5126 31170 5142
rect 30056 5049 30072 5083
rect 30106 5049 30122 5083
rect 30280 5049 30296 5083
rect 30330 5049 30346 5083
rect 30472 5049 30488 5083
rect 30522 5049 30538 5083
rect 30680 5049 30696 5083
rect 30730 5049 30746 5083
rect 30872 5049 30888 5083
rect 30922 5049 30938 5083
rect 31076 5049 31092 5083
rect 31126 5049 31142 5083
rect 34760 5030 34780 6970
rect 34820 5030 34840 6970
rect 34760 4990 34840 5030
rect 29640 4970 34840 4990
rect 29580 4930 29680 4970
rect 34780 4930 34840 4970
rect 29580 4910 34840 4930
rect 28208 4710 28242 4772
rect 25686 4676 25782 4710
rect 28146 4676 28242 4710
rect 29560 4810 34800 4830
rect 29560 4770 29660 4810
rect 34700 4790 34800 4810
rect 34700 4770 34740 4790
rect 29560 4750 34740 4770
rect 1290 4460 3410 4480
rect 1290 4440 1390 4460
rect 1290 3040 1310 4440
rect 1350 4420 1390 4440
rect 3310 4440 3410 4460
rect 3310 4420 3350 4440
rect 1350 4400 3350 4420
rect 1350 3580 1370 4400
rect 1466 4277 1482 4311
rect 1516 4277 1532 4311
rect 1979 4270 1995 4304
rect 2029 4270 2045 4304
rect 2171 4270 2187 4304
rect 2221 4270 2237 4304
rect 2363 4270 2379 4304
rect 2413 4270 2429 4304
rect 2555 4270 2571 4304
rect 2605 4270 2621 4304
rect 2747 4270 2763 4304
rect 2797 4270 2813 4304
rect 2939 4270 2955 4304
rect 2989 4270 3005 4304
rect 3166 4277 3182 4311
rect 3216 4277 3232 4311
rect 1360 3490 1370 3580
rect 1350 3100 1370 3490
rect 1438 4218 1472 4234
rect 1438 3226 1472 3242
rect 1526 4218 1560 4234
rect 1851 4211 1885 4227
rect 1666 3877 1682 3911
rect 1716 3877 1732 3911
rect 1526 3226 1560 3242
rect 1638 3818 1672 3834
rect 1638 3226 1672 3242
rect 1726 3818 1760 3834
rect 1726 3226 1760 3242
rect 1851 3219 1885 3235
rect 1947 4211 1981 4227
rect 1947 3219 1981 3235
rect 2043 4211 2077 4227
rect 2043 3219 2077 3235
rect 2139 4211 2173 4227
rect 2139 3219 2173 3235
rect 2235 4211 2269 4227
rect 2235 3219 2269 3235
rect 2331 4211 2365 4227
rect 2331 3219 2365 3235
rect 2427 4211 2461 4227
rect 2427 3219 2461 3235
rect 2523 4211 2557 4227
rect 2523 3219 2557 3235
rect 2619 4211 2653 4227
rect 2619 3219 2653 3235
rect 2715 4211 2749 4227
rect 2715 3219 2749 3235
rect 2811 4211 2845 4227
rect 2811 3219 2845 3235
rect 2907 4211 2941 4227
rect 2907 3219 2941 3235
rect 3003 4211 3037 4227
rect 3003 3219 3037 3235
rect 3138 4218 3172 4234
rect 3138 3226 3172 3242
rect 3226 4218 3260 4234
rect 3226 3226 3260 3242
rect 1466 3149 1482 3183
rect 1516 3149 1532 3183
rect 1666 3149 1682 3183
rect 1716 3149 1732 3183
rect 1883 3142 1899 3176
rect 1933 3142 1949 3176
rect 2075 3142 2091 3176
rect 2125 3142 2141 3176
rect 2267 3142 2283 3176
rect 2317 3142 2333 3176
rect 2459 3142 2475 3176
rect 2509 3142 2525 3176
rect 2651 3142 2667 3176
rect 2701 3142 2717 3176
rect 2843 3142 2859 3176
rect 2893 3142 2909 3176
rect 3166 3149 3182 3183
rect 3216 3149 3232 3183
rect 1350 3080 1390 3100
rect 3330 3080 3350 4400
rect 1350 3060 3350 3080
rect 1350 3040 1390 3060
rect 1290 3020 1390 3040
rect 3310 3040 3350 3060
rect 3390 3040 3410 4440
rect 3310 3020 3410 3040
rect 1290 3000 3410 3020
rect 4590 4460 6710 4480
rect 4590 4440 4690 4460
rect 4590 3040 4610 4440
rect 4650 4420 4690 4440
rect 6610 4440 6710 4460
rect 6610 4420 6650 4440
rect 4650 4400 6650 4420
rect 4650 3580 4670 4400
rect 4766 4277 4782 4311
rect 4816 4277 4832 4311
rect 5279 4270 5295 4304
rect 5329 4270 5345 4304
rect 5471 4270 5487 4304
rect 5521 4270 5537 4304
rect 5663 4270 5679 4304
rect 5713 4270 5729 4304
rect 5855 4270 5871 4304
rect 5905 4270 5921 4304
rect 6047 4270 6063 4304
rect 6097 4270 6113 4304
rect 6239 4270 6255 4304
rect 6289 4270 6305 4304
rect 6466 4277 6482 4311
rect 6516 4277 6532 4311
rect 4660 3490 4670 3580
rect 4650 3100 4670 3490
rect 4738 4218 4772 4234
rect 4738 3226 4772 3242
rect 4826 4218 4860 4234
rect 5151 4211 5185 4227
rect 4966 3877 4982 3911
rect 5016 3877 5032 3911
rect 4826 3226 4860 3242
rect 4938 3818 4972 3834
rect 4938 3226 4972 3242
rect 5026 3818 5060 3834
rect 5026 3226 5060 3242
rect 5151 3219 5185 3235
rect 5247 4211 5281 4227
rect 5247 3219 5281 3235
rect 5343 4211 5377 4227
rect 5343 3219 5377 3235
rect 5439 4211 5473 4227
rect 5439 3219 5473 3235
rect 5535 4211 5569 4227
rect 5535 3219 5569 3235
rect 5631 4211 5665 4227
rect 5631 3219 5665 3235
rect 5727 4211 5761 4227
rect 5727 3219 5761 3235
rect 5823 4211 5857 4227
rect 5823 3219 5857 3235
rect 5919 4211 5953 4227
rect 5919 3219 5953 3235
rect 6015 4211 6049 4227
rect 6015 3219 6049 3235
rect 6111 4211 6145 4227
rect 6111 3219 6145 3235
rect 6207 4211 6241 4227
rect 6207 3219 6241 3235
rect 6303 4211 6337 4227
rect 6303 3219 6337 3235
rect 6438 4218 6472 4234
rect 6438 3226 6472 3242
rect 6526 4218 6560 4234
rect 6526 3226 6560 3242
rect 4766 3149 4782 3183
rect 4816 3149 4832 3183
rect 4966 3149 4982 3183
rect 5016 3149 5032 3183
rect 5183 3142 5199 3176
rect 5233 3142 5249 3176
rect 5375 3142 5391 3176
rect 5425 3142 5441 3176
rect 5567 3142 5583 3176
rect 5617 3142 5633 3176
rect 5759 3142 5775 3176
rect 5809 3142 5825 3176
rect 5951 3142 5967 3176
rect 6001 3142 6017 3176
rect 6143 3142 6159 3176
rect 6193 3142 6209 3176
rect 6466 3149 6482 3183
rect 6516 3149 6532 3183
rect 4650 3080 4690 3100
rect 6630 3080 6650 4400
rect 4650 3060 6650 3080
rect 4650 3040 4690 3060
rect 4590 3020 4690 3040
rect 6610 3040 6650 3060
rect 6690 3040 6710 4440
rect 6610 3020 6710 3040
rect 4590 3000 6710 3020
rect 7890 4460 10010 4480
rect 7890 4440 7990 4460
rect 7890 3040 7910 4440
rect 7950 4420 7990 4440
rect 9910 4440 10010 4460
rect 9910 4420 9950 4440
rect 7950 4400 9950 4420
rect 7950 3580 7970 4400
rect 8066 4277 8082 4311
rect 8116 4277 8132 4311
rect 8579 4270 8595 4304
rect 8629 4270 8645 4304
rect 8771 4270 8787 4304
rect 8821 4270 8837 4304
rect 8963 4270 8979 4304
rect 9013 4270 9029 4304
rect 9155 4270 9171 4304
rect 9205 4270 9221 4304
rect 9347 4270 9363 4304
rect 9397 4270 9413 4304
rect 9539 4270 9555 4304
rect 9589 4270 9605 4304
rect 9766 4277 9782 4311
rect 9816 4277 9832 4311
rect 7960 3490 7970 3580
rect 7950 3100 7970 3490
rect 8038 4218 8072 4234
rect 8038 3226 8072 3242
rect 8126 4218 8160 4234
rect 8451 4211 8485 4227
rect 8266 3877 8282 3911
rect 8316 3877 8332 3911
rect 8126 3226 8160 3242
rect 8238 3818 8272 3834
rect 8238 3226 8272 3242
rect 8326 3818 8360 3834
rect 8326 3226 8360 3242
rect 8451 3219 8485 3235
rect 8547 4211 8581 4227
rect 8547 3219 8581 3235
rect 8643 4211 8677 4227
rect 8643 3219 8677 3235
rect 8739 4211 8773 4227
rect 8739 3219 8773 3235
rect 8835 4211 8869 4227
rect 8835 3219 8869 3235
rect 8931 4211 8965 4227
rect 8931 3219 8965 3235
rect 9027 4211 9061 4227
rect 9027 3219 9061 3235
rect 9123 4211 9157 4227
rect 9123 3219 9157 3235
rect 9219 4211 9253 4227
rect 9219 3219 9253 3235
rect 9315 4211 9349 4227
rect 9315 3219 9349 3235
rect 9411 4211 9445 4227
rect 9411 3219 9445 3235
rect 9507 4211 9541 4227
rect 9507 3219 9541 3235
rect 9603 4211 9637 4227
rect 9603 3219 9637 3235
rect 9738 4218 9772 4234
rect 9738 3226 9772 3242
rect 9826 4218 9860 4234
rect 9826 3226 9860 3242
rect 8066 3149 8082 3183
rect 8116 3149 8132 3183
rect 8266 3149 8282 3183
rect 8316 3149 8332 3183
rect 8483 3142 8499 3176
rect 8533 3142 8549 3176
rect 8675 3142 8691 3176
rect 8725 3142 8741 3176
rect 8867 3142 8883 3176
rect 8917 3142 8933 3176
rect 9059 3142 9075 3176
rect 9109 3142 9125 3176
rect 9251 3142 9267 3176
rect 9301 3142 9317 3176
rect 9443 3142 9459 3176
rect 9493 3142 9509 3176
rect 9766 3149 9782 3183
rect 9816 3149 9832 3183
rect 7950 3080 7990 3100
rect 9930 3080 9950 4400
rect 7950 3060 9950 3080
rect 7950 3040 7990 3060
rect 7890 3020 7990 3040
rect 9910 3040 9950 3060
rect 9990 3040 10010 4440
rect 9910 3020 10010 3040
rect 7890 3000 10010 3020
rect 11190 4460 13310 4480
rect 11190 4440 11290 4460
rect 11190 3040 11210 4440
rect 11250 4420 11290 4440
rect 13210 4440 13310 4460
rect 13210 4420 13250 4440
rect 11250 4400 13250 4420
rect 11250 3580 11270 4400
rect 11366 4277 11382 4311
rect 11416 4277 11432 4311
rect 11879 4270 11895 4304
rect 11929 4270 11945 4304
rect 12071 4270 12087 4304
rect 12121 4270 12137 4304
rect 12263 4270 12279 4304
rect 12313 4270 12329 4304
rect 12455 4270 12471 4304
rect 12505 4270 12521 4304
rect 12647 4270 12663 4304
rect 12697 4270 12713 4304
rect 12839 4270 12855 4304
rect 12889 4270 12905 4304
rect 13066 4277 13082 4311
rect 13116 4277 13132 4311
rect 11260 3490 11270 3580
rect 11250 3100 11270 3490
rect 11338 4218 11372 4234
rect 11338 3226 11372 3242
rect 11426 4218 11460 4234
rect 11751 4211 11785 4227
rect 11566 3877 11582 3911
rect 11616 3877 11632 3911
rect 11426 3226 11460 3242
rect 11538 3818 11572 3834
rect 11538 3226 11572 3242
rect 11626 3818 11660 3834
rect 11626 3226 11660 3242
rect 11751 3219 11785 3235
rect 11847 4211 11881 4227
rect 11847 3219 11881 3235
rect 11943 4211 11977 4227
rect 11943 3219 11977 3235
rect 12039 4211 12073 4227
rect 12039 3219 12073 3235
rect 12135 4211 12169 4227
rect 12135 3219 12169 3235
rect 12231 4211 12265 4227
rect 12231 3219 12265 3235
rect 12327 4211 12361 4227
rect 12327 3219 12361 3235
rect 12423 4211 12457 4227
rect 12423 3219 12457 3235
rect 12519 4211 12553 4227
rect 12519 3219 12553 3235
rect 12615 4211 12649 4227
rect 12615 3219 12649 3235
rect 12711 4211 12745 4227
rect 12711 3219 12745 3235
rect 12807 4211 12841 4227
rect 12807 3219 12841 3235
rect 12903 4211 12937 4227
rect 12903 3219 12937 3235
rect 13038 4218 13072 4234
rect 13038 3226 13072 3242
rect 13126 4218 13160 4234
rect 13126 3226 13160 3242
rect 11366 3149 11382 3183
rect 11416 3149 11432 3183
rect 11566 3149 11582 3183
rect 11616 3149 11632 3183
rect 11783 3142 11799 3176
rect 11833 3142 11849 3176
rect 11975 3142 11991 3176
rect 12025 3142 12041 3176
rect 12167 3142 12183 3176
rect 12217 3142 12233 3176
rect 12359 3142 12375 3176
rect 12409 3142 12425 3176
rect 12551 3142 12567 3176
rect 12601 3142 12617 3176
rect 12743 3142 12759 3176
rect 12793 3142 12809 3176
rect 13066 3149 13082 3183
rect 13116 3149 13132 3183
rect 11250 3080 11290 3100
rect 13230 3080 13250 4400
rect 11250 3060 13250 3080
rect 11250 3040 11290 3060
rect 11190 3020 11290 3040
rect 13210 3040 13250 3060
rect 13290 3040 13310 4440
rect 13210 3020 13310 3040
rect 11190 3000 13310 3020
rect 14790 4460 16910 4480
rect 14790 4440 14890 4460
rect 14790 3040 14810 4440
rect 14850 4420 14890 4440
rect 16810 4440 16910 4460
rect 16810 4420 16850 4440
rect 14850 4400 16850 4420
rect 14850 3580 14870 4400
rect 14966 4277 14982 4311
rect 15016 4277 15032 4311
rect 15479 4270 15495 4304
rect 15529 4270 15545 4304
rect 15671 4270 15687 4304
rect 15721 4270 15737 4304
rect 15863 4270 15879 4304
rect 15913 4270 15929 4304
rect 16055 4270 16071 4304
rect 16105 4270 16121 4304
rect 16247 4270 16263 4304
rect 16297 4270 16313 4304
rect 16439 4270 16455 4304
rect 16489 4270 16505 4304
rect 16666 4277 16682 4311
rect 16716 4277 16732 4311
rect 14860 3490 14870 3580
rect 14850 3100 14870 3490
rect 14938 4218 14972 4234
rect 14938 3226 14972 3242
rect 15026 4218 15060 4234
rect 15351 4211 15385 4227
rect 15166 3877 15182 3911
rect 15216 3877 15232 3911
rect 15026 3226 15060 3242
rect 15138 3818 15172 3834
rect 15138 3226 15172 3242
rect 15226 3818 15260 3834
rect 15226 3226 15260 3242
rect 15351 3219 15385 3235
rect 15447 4211 15481 4227
rect 15447 3219 15481 3235
rect 15543 4211 15577 4227
rect 15543 3219 15577 3235
rect 15639 4211 15673 4227
rect 15639 3219 15673 3235
rect 15735 4211 15769 4227
rect 15735 3219 15769 3235
rect 15831 4211 15865 4227
rect 15831 3219 15865 3235
rect 15927 4211 15961 4227
rect 15927 3219 15961 3235
rect 16023 4211 16057 4227
rect 16023 3219 16057 3235
rect 16119 4211 16153 4227
rect 16119 3219 16153 3235
rect 16215 4211 16249 4227
rect 16215 3219 16249 3235
rect 16311 4211 16345 4227
rect 16311 3219 16345 3235
rect 16407 4211 16441 4227
rect 16407 3219 16441 3235
rect 16503 4211 16537 4227
rect 16503 3219 16537 3235
rect 16638 4218 16672 4234
rect 16638 3226 16672 3242
rect 16726 4218 16760 4234
rect 16726 3226 16760 3242
rect 14966 3149 14982 3183
rect 15016 3149 15032 3183
rect 15166 3149 15182 3183
rect 15216 3149 15232 3183
rect 15383 3142 15399 3176
rect 15433 3142 15449 3176
rect 15575 3142 15591 3176
rect 15625 3142 15641 3176
rect 15767 3142 15783 3176
rect 15817 3142 15833 3176
rect 15959 3142 15975 3176
rect 16009 3142 16025 3176
rect 16151 3142 16167 3176
rect 16201 3142 16217 3176
rect 16343 3142 16359 3176
rect 16393 3142 16409 3176
rect 16666 3149 16682 3183
rect 16716 3149 16732 3183
rect 14850 3080 14890 3100
rect 16830 3080 16850 4400
rect 14850 3060 16850 3080
rect 14850 3040 14890 3060
rect 14790 3020 14890 3040
rect 16810 3040 16850 3060
rect 16890 3040 16910 4440
rect 16810 3020 16910 3040
rect 14790 3000 16910 3020
rect 18290 4460 20410 4480
rect 18290 4440 18390 4460
rect 18290 3040 18310 4440
rect 18350 4420 18390 4440
rect 20310 4440 20410 4460
rect 20310 4420 20350 4440
rect 18350 4400 20350 4420
rect 18350 3580 18370 4400
rect 18466 4277 18482 4311
rect 18516 4277 18532 4311
rect 18979 4270 18995 4304
rect 19029 4270 19045 4304
rect 19171 4270 19187 4304
rect 19221 4270 19237 4304
rect 19363 4270 19379 4304
rect 19413 4270 19429 4304
rect 19555 4270 19571 4304
rect 19605 4270 19621 4304
rect 19747 4270 19763 4304
rect 19797 4270 19813 4304
rect 19939 4270 19955 4304
rect 19989 4270 20005 4304
rect 20166 4277 20182 4311
rect 20216 4277 20232 4311
rect 18360 3490 18370 3580
rect 18350 3100 18370 3490
rect 18438 4218 18472 4234
rect 18438 3226 18472 3242
rect 18526 4218 18560 4234
rect 18851 4211 18885 4227
rect 18666 3877 18682 3911
rect 18716 3877 18732 3911
rect 18526 3226 18560 3242
rect 18638 3818 18672 3834
rect 18638 3226 18672 3242
rect 18726 3818 18760 3834
rect 18726 3226 18760 3242
rect 18851 3219 18885 3235
rect 18947 4211 18981 4227
rect 18947 3219 18981 3235
rect 19043 4211 19077 4227
rect 19043 3219 19077 3235
rect 19139 4211 19173 4227
rect 19139 3219 19173 3235
rect 19235 4211 19269 4227
rect 19235 3219 19269 3235
rect 19331 4211 19365 4227
rect 19331 3219 19365 3235
rect 19427 4211 19461 4227
rect 19427 3219 19461 3235
rect 19523 4211 19557 4227
rect 19523 3219 19557 3235
rect 19619 4211 19653 4227
rect 19619 3219 19653 3235
rect 19715 4211 19749 4227
rect 19715 3219 19749 3235
rect 19811 4211 19845 4227
rect 19811 3219 19845 3235
rect 19907 4211 19941 4227
rect 19907 3219 19941 3235
rect 20003 4211 20037 4227
rect 20003 3219 20037 3235
rect 20138 4218 20172 4234
rect 20138 3226 20172 3242
rect 20226 4218 20260 4234
rect 20226 3226 20260 3242
rect 18466 3149 18482 3183
rect 18516 3149 18532 3183
rect 18666 3149 18682 3183
rect 18716 3149 18732 3183
rect 18883 3142 18899 3176
rect 18933 3142 18949 3176
rect 19075 3142 19091 3176
rect 19125 3142 19141 3176
rect 19267 3142 19283 3176
rect 19317 3142 19333 3176
rect 19459 3142 19475 3176
rect 19509 3142 19525 3176
rect 19651 3142 19667 3176
rect 19701 3142 19717 3176
rect 19843 3142 19859 3176
rect 19893 3142 19909 3176
rect 20166 3149 20182 3183
rect 20216 3149 20232 3183
rect 18350 3080 18390 3100
rect 20330 3080 20350 4400
rect 18350 3060 20350 3080
rect 18350 3040 18390 3060
rect 18290 3020 18390 3040
rect 20310 3040 20350 3060
rect 20390 3040 20410 4440
rect 20310 3020 20410 3040
rect 18290 3000 20410 3020
rect 21990 4460 24110 4480
rect 21990 4440 22090 4460
rect 21990 3040 22010 4440
rect 22050 4420 22090 4440
rect 24010 4440 24110 4460
rect 24010 4420 24050 4440
rect 22050 4400 24050 4420
rect 22050 3580 22070 4400
rect 22166 4277 22182 4311
rect 22216 4277 22232 4311
rect 22679 4270 22695 4304
rect 22729 4270 22745 4304
rect 22871 4270 22887 4304
rect 22921 4270 22937 4304
rect 23063 4270 23079 4304
rect 23113 4270 23129 4304
rect 23255 4270 23271 4304
rect 23305 4270 23321 4304
rect 23447 4270 23463 4304
rect 23497 4270 23513 4304
rect 23639 4270 23655 4304
rect 23689 4270 23705 4304
rect 23866 4277 23882 4311
rect 23916 4277 23932 4311
rect 22060 3490 22070 3580
rect 22050 3100 22070 3490
rect 22138 4218 22172 4234
rect 22138 3226 22172 3242
rect 22226 4218 22260 4234
rect 22551 4211 22585 4227
rect 22366 3877 22382 3911
rect 22416 3877 22432 3911
rect 22226 3226 22260 3242
rect 22338 3818 22372 3834
rect 22338 3226 22372 3242
rect 22426 3818 22460 3834
rect 22426 3226 22460 3242
rect 22551 3219 22585 3235
rect 22647 4211 22681 4227
rect 22647 3219 22681 3235
rect 22743 4211 22777 4227
rect 22743 3219 22777 3235
rect 22839 4211 22873 4227
rect 22839 3219 22873 3235
rect 22935 4211 22969 4227
rect 22935 3219 22969 3235
rect 23031 4211 23065 4227
rect 23031 3219 23065 3235
rect 23127 4211 23161 4227
rect 23127 3219 23161 3235
rect 23223 4211 23257 4227
rect 23223 3219 23257 3235
rect 23319 4211 23353 4227
rect 23319 3219 23353 3235
rect 23415 4211 23449 4227
rect 23415 3219 23449 3235
rect 23511 4211 23545 4227
rect 23511 3219 23545 3235
rect 23607 4211 23641 4227
rect 23607 3219 23641 3235
rect 23703 4211 23737 4227
rect 23703 3219 23737 3235
rect 23838 4218 23872 4234
rect 23838 3226 23872 3242
rect 23926 4218 23960 4234
rect 23926 3226 23960 3242
rect 22166 3149 22182 3183
rect 22216 3149 22232 3183
rect 22366 3149 22382 3183
rect 22416 3149 22432 3183
rect 22583 3142 22599 3176
rect 22633 3142 22649 3176
rect 22775 3142 22791 3176
rect 22825 3142 22841 3176
rect 22967 3142 22983 3176
rect 23017 3142 23033 3176
rect 23159 3142 23175 3176
rect 23209 3142 23225 3176
rect 23351 3142 23367 3176
rect 23401 3142 23417 3176
rect 23543 3142 23559 3176
rect 23593 3142 23609 3176
rect 23866 3149 23882 3183
rect 23916 3149 23932 3183
rect 22050 3080 22090 3100
rect 24030 3080 24050 4400
rect 22050 3060 24050 3080
rect 22050 3040 22090 3060
rect 21990 3020 22090 3040
rect 24010 3040 24050 3060
rect 24090 3040 24110 4440
rect 24010 3020 24110 3040
rect 21990 3000 24110 3020
rect 25790 4460 27910 4480
rect 25790 4440 25890 4460
rect 25790 3040 25810 4440
rect 25850 4420 25890 4440
rect 27810 4440 27910 4460
rect 27810 4420 27850 4440
rect 25850 4400 27850 4420
rect 25850 3580 25870 4400
rect 25966 4277 25982 4311
rect 26016 4277 26032 4311
rect 26479 4270 26495 4304
rect 26529 4270 26545 4304
rect 26671 4270 26687 4304
rect 26721 4270 26737 4304
rect 26863 4270 26879 4304
rect 26913 4270 26929 4304
rect 27055 4270 27071 4304
rect 27105 4270 27121 4304
rect 27247 4270 27263 4304
rect 27297 4270 27313 4304
rect 27439 4270 27455 4304
rect 27489 4270 27505 4304
rect 27666 4277 27682 4311
rect 27716 4277 27732 4311
rect 25860 3490 25870 3580
rect 25850 3100 25870 3490
rect 25938 4218 25972 4234
rect 25938 3226 25972 3242
rect 26026 4218 26060 4234
rect 26351 4211 26385 4227
rect 26166 3877 26182 3911
rect 26216 3877 26232 3911
rect 26026 3226 26060 3242
rect 26138 3818 26172 3834
rect 26138 3226 26172 3242
rect 26226 3818 26260 3834
rect 26226 3226 26260 3242
rect 26351 3219 26385 3235
rect 26447 4211 26481 4227
rect 26447 3219 26481 3235
rect 26543 4211 26577 4227
rect 26543 3219 26577 3235
rect 26639 4211 26673 4227
rect 26639 3219 26673 3235
rect 26735 4211 26769 4227
rect 26735 3219 26769 3235
rect 26831 4211 26865 4227
rect 26831 3219 26865 3235
rect 26927 4211 26961 4227
rect 26927 3219 26961 3235
rect 27023 4211 27057 4227
rect 27023 3219 27057 3235
rect 27119 4211 27153 4227
rect 27119 3219 27153 3235
rect 27215 4211 27249 4227
rect 27215 3219 27249 3235
rect 27311 4211 27345 4227
rect 27311 3219 27345 3235
rect 27407 4211 27441 4227
rect 27407 3219 27441 3235
rect 27503 4211 27537 4227
rect 27503 3219 27537 3235
rect 27638 4218 27672 4234
rect 27638 3226 27672 3242
rect 27726 4218 27760 4234
rect 27726 3226 27760 3242
rect 25966 3149 25982 3183
rect 26016 3149 26032 3183
rect 26166 3149 26182 3183
rect 26216 3149 26232 3183
rect 26383 3142 26399 3176
rect 26433 3142 26449 3176
rect 26575 3142 26591 3176
rect 26625 3142 26641 3176
rect 26767 3142 26783 3176
rect 26817 3142 26833 3176
rect 26959 3142 26975 3176
rect 27009 3142 27025 3176
rect 27151 3142 27167 3176
rect 27201 3142 27217 3176
rect 27343 3142 27359 3176
rect 27393 3142 27409 3176
rect 27666 3149 27682 3183
rect 27716 3149 27732 3183
rect 25850 3080 25890 3100
rect 27830 3080 27850 4400
rect 25850 3060 27850 3080
rect 25850 3040 25890 3060
rect 25790 3020 25890 3040
rect 27810 3040 27850 3060
rect 27890 3040 27910 4440
rect 29560 4110 29580 4750
rect 29620 4110 29640 4750
rect 29918 4596 29934 4630
rect 30102 4596 30118 4630
rect 30298 4596 30314 4630
rect 30482 4596 30498 4630
rect 30698 4596 30714 4630
rect 30882 4596 30898 4630
rect 31078 4596 31094 4630
rect 31262 4596 31278 4630
rect 31336 4596 31352 4630
rect 31520 4596 31536 4630
rect 31594 4596 31610 4630
rect 31778 4596 31794 4630
rect 31852 4596 31868 4630
rect 32036 4596 32052 4630
rect 32110 4596 32126 4630
rect 32294 4596 32310 4630
rect 32368 4596 32384 4630
rect 32552 4596 32568 4630
rect 32626 4596 32642 4630
rect 32810 4596 32826 4630
rect 32884 4596 32900 4630
rect 33068 4596 33084 4630
rect 33142 4596 33158 4630
rect 33326 4596 33342 4630
rect 33518 4596 33534 4630
rect 33702 4596 33718 4630
rect 29872 4546 29906 4562
rect 29872 4354 29906 4370
rect 30130 4546 30164 4562
rect 30130 4354 30164 4370
rect 30252 4546 30286 4562
rect 30252 4354 30286 4370
rect 30510 4546 30544 4562
rect 30510 4354 30544 4370
rect 30652 4546 30686 4562
rect 30652 4354 30686 4370
rect 30910 4546 30944 4562
rect 30910 4354 30944 4370
rect 31032 4546 31066 4562
rect 31032 4354 31066 4370
rect 31290 4546 31324 4562
rect 31290 4354 31324 4370
rect 31548 4546 31582 4562
rect 31548 4354 31582 4370
rect 31806 4546 31840 4562
rect 31806 4354 31840 4370
rect 32064 4546 32098 4562
rect 32064 4354 32098 4370
rect 32322 4546 32356 4562
rect 32322 4354 32356 4370
rect 32580 4546 32614 4562
rect 32580 4354 32614 4370
rect 32838 4546 32872 4562
rect 32838 4354 32872 4370
rect 33096 4546 33130 4562
rect 33096 4354 33130 4370
rect 33354 4546 33388 4562
rect 33354 4354 33388 4370
rect 33472 4546 33506 4562
rect 33472 4354 33506 4370
rect 33730 4546 33764 4562
rect 33730 4354 33764 4370
rect 29918 4286 29934 4320
rect 30102 4286 30118 4320
rect 30298 4286 30314 4320
rect 30482 4286 30498 4320
rect 30698 4286 30714 4320
rect 30882 4286 30898 4320
rect 31078 4286 31094 4320
rect 31262 4286 31278 4320
rect 31336 4286 31352 4320
rect 31520 4286 31536 4320
rect 31594 4286 31610 4320
rect 31778 4286 31794 4320
rect 31852 4286 31868 4320
rect 32036 4286 32052 4320
rect 32110 4286 32126 4320
rect 32294 4286 32310 4320
rect 32368 4286 32384 4320
rect 32552 4286 32568 4320
rect 32626 4286 32642 4320
rect 32810 4286 32826 4320
rect 32884 4286 32900 4320
rect 33068 4286 33084 4320
rect 33142 4286 33158 4320
rect 33326 4286 33342 4320
rect 33518 4286 33534 4320
rect 33702 4286 33718 4320
rect 34720 4130 34740 4750
rect 34780 4130 34800 4790
rect 34720 4110 34800 4130
rect 29560 4090 34800 4110
rect 29560 4050 29660 4090
rect 34720 4050 34800 4090
rect 29560 4030 34800 4050
rect 27810 3020 27910 3040
rect 25790 3000 27910 3020
rect 1280 2900 3410 2930
rect 440 2690 620 2706
rect 440 2494 620 2510
rect 1280 2670 1310 2900
rect 1350 2860 1390 2900
rect 3310 2890 3410 2900
rect 3310 2860 3350 2890
rect 1350 2840 3350 2860
rect 1350 2670 1370 2840
rect 1470 2746 1486 2780
rect 1520 2746 1536 2780
rect 1670 2746 1686 2780
rect 1720 2746 1736 2780
rect 1983 2739 1999 2773
rect 2033 2739 2049 2773
rect 2175 2739 2191 2773
rect 2225 2739 2241 2773
rect 2367 2739 2383 2773
rect 2417 2739 2433 2773
rect 2559 2739 2575 2773
rect 2609 2739 2625 2773
rect 2751 2739 2767 2773
rect 2801 2739 2817 2773
rect 2943 2739 2959 2773
rect 2993 2739 3009 2773
rect 3150 2746 3166 2780
rect 3200 2746 3216 2780
rect 1280 2540 1300 2670
rect 1360 2540 1370 2670
rect 1280 1520 1310 2540
rect 1350 1570 1370 2540
rect 1442 2696 1476 2712
rect 1442 1704 1476 1720
rect 1530 2696 1564 2712
rect 1642 2696 1676 2712
rect 1642 2504 1676 2520
rect 1730 2696 1764 2712
rect 1730 2504 1764 2520
rect 1855 2689 1889 2705
rect 1670 2436 1686 2470
rect 1720 2436 1736 2470
rect 1530 1704 1564 1720
rect 1855 1697 1889 1713
rect 1951 2689 1985 2705
rect 1951 1697 1985 1713
rect 2047 2689 2081 2705
rect 2047 1697 2081 1713
rect 2143 2689 2177 2705
rect 2143 1697 2177 1713
rect 2239 2689 2273 2705
rect 2239 1697 2273 1713
rect 2335 2689 2369 2705
rect 2335 1697 2369 1713
rect 2431 2689 2465 2705
rect 2431 1697 2465 1713
rect 2527 2689 2561 2705
rect 2527 1697 2561 1713
rect 2623 2689 2657 2705
rect 2623 1697 2657 1713
rect 2719 2689 2753 2705
rect 2719 1697 2753 1713
rect 2815 2689 2849 2705
rect 2815 1697 2849 1713
rect 2911 2689 2945 2705
rect 2911 1697 2945 1713
rect 3007 2689 3041 2705
rect 3007 1697 3041 1713
rect 3122 2696 3156 2712
rect 3122 1704 3156 1720
rect 3210 2696 3244 2712
rect 3210 1704 3244 1720
rect 1470 1636 1486 1670
rect 1520 1636 1536 1670
rect 1887 1629 1903 1663
rect 1937 1629 1953 1663
rect 2079 1629 2095 1663
rect 2129 1629 2145 1663
rect 2271 1629 2287 1663
rect 2321 1629 2337 1663
rect 2463 1629 2479 1663
rect 2513 1629 2529 1663
rect 2655 1629 2671 1663
rect 2705 1629 2721 1663
rect 2847 1629 2863 1663
rect 2897 1629 2913 1663
rect 3150 1636 3166 1670
rect 3200 1636 3216 1670
rect 3330 1570 3350 2840
rect 1350 1540 3350 1570
rect 1350 1520 1390 1540
rect 1280 1500 1390 1520
rect 3310 1510 3350 1540
rect 3390 1510 3410 2890
rect 3310 1500 3410 1510
rect 1280 1480 3410 1500
rect 4580 2900 6710 2930
rect 4580 2670 4610 2900
rect 4650 2860 4690 2900
rect 6610 2890 6710 2900
rect 6610 2860 6650 2890
rect 4650 2840 6650 2860
rect 4650 2670 4670 2840
rect 4770 2746 4786 2780
rect 4820 2746 4836 2780
rect 4970 2746 4986 2780
rect 5020 2746 5036 2780
rect 5283 2739 5299 2773
rect 5333 2739 5349 2773
rect 5475 2739 5491 2773
rect 5525 2739 5541 2773
rect 5667 2739 5683 2773
rect 5717 2739 5733 2773
rect 5859 2739 5875 2773
rect 5909 2739 5925 2773
rect 6051 2739 6067 2773
rect 6101 2739 6117 2773
rect 6243 2739 6259 2773
rect 6293 2739 6309 2773
rect 6450 2746 6466 2780
rect 6500 2746 6516 2780
rect 4580 2540 4600 2670
rect 4660 2540 4670 2670
rect 4580 1520 4610 2540
rect 4650 1570 4670 2540
rect 4742 2696 4776 2712
rect 4742 1704 4776 1720
rect 4830 2696 4864 2712
rect 4942 2696 4976 2712
rect 4942 2504 4976 2520
rect 5030 2696 5064 2712
rect 5030 2504 5064 2520
rect 5155 2689 5189 2705
rect 4970 2436 4986 2470
rect 5020 2436 5036 2470
rect 4830 1704 4864 1720
rect 5155 1697 5189 1713
rect 5251 2689 5285 2705
rect 5251 1697 5285 1713
rect 5347 2689 5381 2705
rect 5347 1697 5381 1713
rect 5443 2689 5477 2705
rect 5443 1697 5477 1713
rect 5539 2689 5573 2705
rect 5539 1697 5573 1713
rect 5635 2689 5669 2705
rect 5635 1697 5669 1713
rect 5731 2689 5765 2705
rect 5731 1697 5765 1713
rect 5827 2689 5861 2705
rect 5827 1697 5861 1713
rect 5923 2689 5957 2705
rect 5923 1697 5957 1713
rect 6019 2689 6053 2705
rect 6019 1697 6053 1713
rect 6115 2689 6149 2705
rect 6115 1697 6149 1713
rect 6211 2689 6245 2705
rect 6211 1697 6245 1713
rect 6307 2689 6341 2705
rect 6307 1697 6341 1713
rect 6422 2696 6456 2712
rect 6422 1704 6456 1720
rect 6510 2696 6544 2712
rect 6510 1704 6544 1720
rect 4770 1636 4786 1670
rect 4820 1636 4836 1670
rect 5187 1629 5203 1663
rect 5237 1629 5253 1663
rect 5379 1629 5395 1663
rect 5429 1629 5445 1663
rect 5571 1629 5587 1663
rect 5621 1629 5637 1663
rect 5763 1629 5779 1663
rect 5813 1629 5829 1663
rect 5955 1629 5971 1663
rect 6005 1629 6021 1663
rect 6147 1629 6163 1663
rect 6197 1629 6213 1663
rect 6450 1636 6466 1670
rect 6500 1636 6516 1670
rect 6630 1570 6650 2840
rect 4650 1540 6650 1570
rect 4650 1520 4690 1540
rect 4580 1500 4690 1520
rect 6610 1510 6650 1540
rect 6690 1510 6710 2890
rect 6610 1500 6710 1510
rect 4580 1480 6710 1500
rect 7880 2900 10010 2930
rect 7880 2670 7910 2900
rect 7950 2860 7990 2900
rect 9910 2890 10010 2900
rect 9910 2860 9950 2890
rect 7950 2840 9950 2860
rect 7950 2670 7970 2840
rect 8070 2746 8086 2780
rect 8120 2746 8136 2780
rect 8270 2746 8286 2780
rect 8320 2746 8336 2780
rect 8583 2739 8599 2773
rect 8633 2739 8649 2773
rect 8775 2739 8791 2773
rect 8825 2739 8841 2773
rect 8967 2739 8983 2773
rect 9017 2739 9033 2773
rect 9159 2739 9175 2773
rect 9209 2739 9225 2773
rect 9351 2739 9367 2773
rect 9401 2739 9417 2773
rect 9543 2739 9559 2773
rect 9593 2739 9609 2773
rect 9750 2746 9766 2780
rect 9800 2746 9816 2780
rect 7880 2540 7900 2670
rect 7960 2540 7970 2670
rect 7880 1520 7910 2540
rect 7950 1570 7970 2540
rect 8042 2696 8076 2712
rect 8042 1704 8076 1720
rect 8130 2696 8164 2712
rect 8242 2696 8276 2712
rect 8242 2504 8276 2520
rect 8330 2696 8364 2712
rect 8330 2504 8364 2520
rect 8455 2689 8489 2705
rect 8270 2436 8286 2470
rect 8320 2436 8336 2470
rect 8130 1704 8164 1720
rect 8455 1697 8489 1713
rect 8551 2689 8585 2705
rect 8551 1697 8585 1713
rect 8647 2689 8681 2705
rect 8647 1697 8681 1713
rect 8743 2689 8777 2705
rect 8743 1697 8777 1713
rect 8839 2689 8873 2705
rect 8839 1697 8873 1713
rect 8935 2689 8969 2705
rect 8935 1697 8969 1713
rect 9031 2689 9065 2705
rect 9031 1697 9065 1713
rect 9127 2689 9161 2705
rect 9127 1697 9161 1713
rect 9223 2689 9257 2705
rect 9223 1697 9257 1713
rect 9319 2689 9353 2705
rect 9319 1697 9353 1713
rect 9415 2689 9449 2705
rect 9415 1697 9449 1713
rect 9511 2689 9545 2705
rect 9511 1697 9545 1713
rect 9607 2689 9641 2705
rect 9607 1697 9641 1713
rect 9722 2696 9756 2712
rect 9722 1704 9756 1720
rect 9810 2696 9844 2712
rect 9810 1704 9844 1720
rect 8070 1636 8086 1670
rect 8120 1636 8136 1670
rect 8487 1629 8503 1663
rect 8537 1629 8553 1663
rect 8679 1629 8695 1663
rect 8729 1629 8745 1663
rect 8871 1629 8887 1663
rect 8921 1629 8937 1663
rect 9063 1629 9079 1663
rect 9113 1629 9129 1663
rect 9255 1629 9271 1663
rect 9305 1629 9321 1663
rect 9447 1629 9463 1663
rect 9497 1629 9513 1663
rect 9750 1636 9766 1670
rect 9800 1636 9816 1670
rect 9930 1570 9950 2840
rect 7950 1540 9950 1570
rect 7950 1520 7990 1540
rect 7880 1500 7990 1520
rect 9910 1510 9950 1540
rect 9990 1510 10010 2890
rect 9910 1500 10010 1510
rect 7880 1480 10010 1500
rect 11180 2900 13310 2930
rect 11180 2670 11210 2900
rect 11250 2860 11290 2900
rect 13210 2890 13310 2900
rect 13210 2860 13250 2890
rect 11250 2840 13250 2860
rect 11250 2670 11270 2840
rect 11370 2746 11386 2780
rect 11420 2746 11436 2780
rect 11570 2746 11586 2780
rect 11620 2746 11636 2780
rect 11883 2739 11899 2773
rect 11933 2739 11949 2773
rect 12075 2739 12091 2773
rect 12125 2739 12141 2773
rect 12267 2739 12283 2773
rect 12317 2739 12333 2773
rect 12459 2739 12475 2773
rect 12509 2739 12525 2773
rect 12651 2739 12667 2773
rect 12701 2739 12717 2773
rect 12843 2739 12859 2773
rect 12893 2739 12909 2773
rect 13050 2746 13066 2780
rect 13100 2746 13116 2780
rect 11180 2540 11200 2670
rect 11260 2540 11270 2670
rect 11180 1520 11210 2540
rect 11250 1570 11270 2540
rect 11342 2696 11376 2712
rect 11342 1704 11376 1720
rect 11430 2696 11464 2712
rect 11542 2696 11576 2712
rect 11542 2504 11576 2520
rect 11630 2696 11664 2712
rect 11630 2504 11664 2520
rect 11755 2689 11789 2705
rect 11570 2436 11586 2470
rect 11620 2436 11636 2470
rect 11430 1704 11464 1720
rect 11755 1697 11789 1713
rect 11851 2689 11885 2705
rect 11851 1697 11885 1713
rect 11947 2689 11981 2705
rect 11947 1697 11981 1713
rect 12043 2689 12077 2705
rect 12043 1697 12077 1713
rect 12139 2689 12173 2705
rect 12139 1697 12173 1713
rect 12235 2689 12269 2705
rect 12235 1697 12269 1713
rect 12331 2689 12365 2705
rect 12331 1697 12365 1713
rect 12427 2689 12461 2705
rect 12427 1697 12461 1713
rect 12523 2689 12557 2705
rect 12523 1697 12557 1713
rect 12619 2689 12653 2705
rect 12619 1697 12653 1713
rect 12715 2689 12749 2705
rect 12715 1697 12749 1713
rect 12811 2689 12845 2705
rect 12811 1697 12845 1713
rect 12907 2689 12941 2705
rect 12907 1697 12941 1713
rect 13022 2696 13056 2712
rect 13022 1704 13056 1720
rect 13110 2696 13144 2712
rect 13110 1704 13144 1720
rect 11370 1636 11386 1670
rect 11420 1636 11436 1670
rect 11787 1629 11803 1663
rect 11837 1629 11853 1663
rect 11979 1629 11995 1663
rect 12029 1629 12045 1663
rect 12171 1629 12187 1663
rect 12221 1629 12237 1663
rect 12363 1629 12379 1663
rect 12413 1629 12429 1663
rect 12555 1629 12571 1663
rect 12605 1629 12621 1663
rect 12747 1629 12763 1663
rect 12797 1629 12813 1663
rect 13050 1636 13066 1670
rect 13100 1636 13116 1670
rect 13230 1570 13250 2840
rect 11250 1540 13250 1570
rect 11250 1520 11290 1540
rect 11180 1500 11290 1520
rect 13210 1510 13250 1540
rect 13290 1510 13310 2890
rect 13210 1500 13310 1510
rect 11180 1480 13310 1500
rect 14780 2900 16910 2930
rect 14780 2670 14810 2900
rect 14850 2860 14890 2900
rect 16810 2890 16910 2900
rect 16810 2860 16850 2890
rect 14850 2840 16850 2860
rect 14850 2670 14870 2840
rect 14970 2746 14986 2780
rect 15020 2746 15036 2780
rect 15170 2746 15186 2780
rect 15220 2746 15236 2780
rect 15483 2739 15499 2773
rect 15533 2739 15549 2773
rect 15675 2739 15691 2773
rect 15725 2739 15741 2773
rect 15867 2739 15883 2773
rect 15917 2739 15933 2773
rect 16059 2739 16075 2773
rect 16109 2739 16125 2773
rect 16251 2739 16267 2773
rect 16301 2739 16317 2773
rect 16443 2739 16459 2773
rect 16493 2739 16509 2773
rect 16650 2746 16666 2780
rect 16700 2746 16716 2780
rect 14780 2540 14800 2670
rect 14860 2540 14870 2670
rect 14780 1520 14810 2540
rect 14850 1570 14870 2540
rect 14942 2696 14976 2712
rect 14942 1704 14976 1720
rect 15030 2696 15064 2712
rect 15142 2696 15176 2712
rect 15142 2504 15176 2520
rect 15230 2696 15264 2712
rect 15230 2504 15264 2520
rect 15355 2689 15389 2705
rect 15170 2436 15186 2470
rect 15220 2436 15236 2470
rect 15030 1704 15064 1720
rect 15355 1697 15389 1713
rect 15451 2689 15485 2705
rect 15451 1697 15485 1713
rect 15547 2689 15581 2705
rect 15547 1697 15581 1713
rect 15643 2689 15677 2705
rect 15643 1697 15677 1713
rect 15739 2689 15773 2705
rect 15739 1697 15773 1713
rect 15835 2689 15869 2705
rect 15835 1697 15869 1713
rect 15931 2689 15965 2705
rect 15931 1697 15965 1713
rect 16027 2689 16061 2705
rect 16027 1697 16061 1713
rect 16123 2689 16157 2705
rect 16123 1697 16157 1713
rect 16219 2689 16253 2705
rect 16219 1697 16253 1713
rect 16315 2689 16349 2705
rect 16315 1697 16349 1713
rect 16411 2689 16445 2705
rect 16411 1697 16445 1713
rect 16507 2689 16541 2705
rect 16507 1697 16541 1713
rect 16622 2696 16656 2712
rect 16622 1704 16656 1720
rect 16710 2696 16744 2712
rect 16710 1704 16744 1720
rect 14970 1636 14986 1670
rect 15020 1636 15036 1670
rect 15387 1629 15403 1663
rect 15437 1629 15453 1663
rect 15579 1629 15595 1663
rect 15629 1629 15645 1663
rect 15771 1629 15787 1663
rect 15821 1629 15837 1663
rect 15963 1629 15979 1663
rect 16013 1629 16029 1663
rect 16155 1629 16171 1663
rect 16205 1629 16221 1663
rect 16347 1629 16363 1663
rect 16397 1629 16413 1663
rect 16650 1636 16666 1670
rect 16700 1636 16716 1670
rect 16830 1570 16850 2840
rect 14850 1540 16850 1570
rect 14850 1520 14890 1540
rect 14780 1500 14890 1520
rect 16810 1510 16850 1540
rect 16890 1510 16910 2890
rect 16810 1500 16910 1510
rect 14780 1480 16910 1500
rect 18280 2900 20410 2930
rect 18280 2670 18310 2900
rect 18350 2860 18390 2900
rect 20310 2890 20410 2900
rect 20310 2860 20350 2890
rect 18350 2840 20350 2860
rect 18350 2670 18370 2840
rect 18470 2746 18486 2780
rect 18520 2746 18536 2780
rect 18670 2746 18686 2780
rect 18720 2746 18736 2780
rect 18983 2739 18999 2773
rect 19033 2739 19049 2773
rect 19175 2739 19191 2773
rect 19225 2739 19241 2773
rect 19367 2739 19383 2773
rect 19417 2739 19433 2773
rect 19559 2739 19575 2773
rect 19609 2739 19625 2773
rect 19751 2739 19767 2773
rect 19801 2739 19817 2773
rect 19943 2739 19959 2773
rect 19993 2739 20009 2773
rect 20150 2746 20166 2780
rect 20200 2746 20216 2780
rect 18280 2540 18300 2670
rect 18360 2540 18370 2670
rect 18280 1520 18310 2540
rect 18350 1570 18370 2540
rect 18442 2696 18476 2712
rect 18442 1704 18476 1720
rect 18530 2696 18564 2712
rect 18642 2696 18676 2712
rect 18642 2504 18676 2520
rect 18730 2696 18764 2712
rect 18730 2504 18764 2520
rect 18855 2689 18889 2705
rect 18670 2436 18686 2470
rect 18720 2436 18736 2470
rect 18530 1704 18564 1720
rect 18855 1697 18889 1713
rect 18951 2689 18985 2705
rect 18951 1697 18985 1713
rect 19047 2689 19081 2705
rect 19047 1697 19081 1713
rect 19143 2689 19177 2705
rect 19143 1697 19177 1713
rect 19239 2689 19273 2705
rect 19239 1697 19273 1713
rect 19335 2689 19369 2705
rect 19335 1697 19369 1713
rect 19431 2689 19465 2705
rect 19431 1697 19465 1713
rect 19527 2689 19561 2705
rect 19527 1697 19561 1713
rect 19623 2689 19657 2705
rect 19623 1697 19657 1713
rect 19719 2689 19753 2705
rect 19719 1697 19753 1713
rect 19815 2689 19849 2705
rect 19815 1697 19849 1713
rect 19911 2689 19945 2705
rect 19911 1697 19945 1713
rect 20007 2689 20041 2705
rect 20007 1697 20041 1713
rect 20122 2696 20156 2712
rect 20122 1704 20156 1720
rect 20210 2696 20244 2712
rect 20210 1704 20244 1720
rect 18470 1636 18486 1670
rect 18520 1636 18536 1670
rect 18887 1629 18903 1663
rect 18937 1629 18953 1663
rect 19079 1629 19095 1663
rect 19129 1629 19145 1663
rect 19271 1629 19287 1663
rect 19321 1629 19337 1663
rect 19463 1629 19479 1663
rect 19513 1629 19529 1663
rect 19655 1629 19671 1663
rect 19705 1629 19721 1663
rect 19847 1629 19863 1663
rect 19897 1629 19913 1663
rect 20150 1636 20166 1670
rect 20200 1636 20216 1670
rect 20330 1570 20350 2840
rect 18350 1540 20350 1570
rect 18350 1520 18390 1540
rect 18280 1500 18390 1520
rect 20310 1510 20350 1540
rect 20390 1510 20410 2890
rect 20310 1500 20410 1510
rect 18280 1480 20410 1500
rect 21980 2900 24110 2930
rect 21980 2670 22010 2900
rect 22050 2860 22090 2900
rect 24010 2890 24110 2900
rect 24010 2860 24050 2890
rect 22050 2840 24050 2860
rect 22050 2670 22070 2840
rect 22170 2746 22186 2780
rect 22220 2746 22236 2780
rect 22370 2746 22386 2780
rect 22420 2746 22436 2780
rect 22683 2739 22699 2773
rect 22733 2739 22749 2773
rect 22875 2739 22891 2773
rect 22925 2739 22941 2773
rect 23067 2739 23083 2773
rect 23117 2739 23133 2773
rect 23259 2739 23275 2773
rect 23309 2739 23325 2773
rect 23451 2739 23467 2773
rect 23501 2739 23517 2773
rect 23643 2739 23659 2773
rect 23693 2739 23709 2773
rect 23850 2746 23866 2780
rect 23900 2746 23916 2780
rect 21980 2540 22000 2670
rect 22060 2540 22070 2670
rect 21980 1520 22010 2540
rect 22050 1570 22070 2540
rect 22142 2696 22176 2712
rect 22142 1704 22176 1720
rect 22230 2696 22264 2712
rect 22342 2696 22376 2712
rect 22342 2504 22376 2520
rect 22430 2696 22464 2712
rect 22430 2504 22464 2520
rect 22555 2689 22589 2705
rect 22370 2436 22386 2470
rect 22420 2436 22436 2470
rect 22230 1704 22264 1720
rect 22555 1697 22589 1713
rect 22651 2689 22685 2705
rect 22651 1697 22685 1713
rect 22747 2689 22781 2705
rect 22747 1697 22781 1713
rect 22843 2689 22877 2705
rect 22843 1697 22877 1713
rect 22939 2689 22973 2705
rect 22939 1697 22973 1713
rect 23035 2689 23069 2705
rect 23035 1697 23069 1713
rect 23131 2689 23165 2705
rect 23131 1697 23165 1713
rect 23227 2689 23261 2705
rect 23227 1697 23261 1713
rect 23323 2689 23357 2705
rect 23323 1697 23357 1713
rect 23419 2689 23453 2705
rect 23419 1697 23453 1713
rect 23515 2689 23549 2705
rect 23515 1697 23549 1713
rect 23611 2689 23645 2705
rect 23611 1697 23645 1713
rect 23707 2689 23741 2705
rect 23707 1697 23741 1713
rect 23822 2696 23856 2712
rect 23822 1704 23856 1720
rect 23910 2696 23944 2712
rect 23910 1704 23944 1720
rect 22170 1636 22186 1670
rect 22220 1636 22236 1670
rect 22587 1629 22603 1663
rect 22637 1629 22653 1663
rect 22779 1629 22795 1663
rect 22829 1629 22845 1663
rect 22971 1629 22987 1663
rect 23021 1629 23037 1663
rect 23163 1629 23179 1663
rect 23213 1629 23229 1663
rect 23355 1629 23371 1663
rect 23405 1629 23421 1663
rect 23547 1629 23563 1663
rect 23597 1629 23613 1663
rect 23850 1636 23866 1670
rect 23900 1636 23916 1670
rect 24030 1570 24050 2840
rect 22050 1540 24050 1570
rect 22050 1520 22090 1540
rect 21980 1500 22090 1520
rect 24010 1510 24050 1540
rect 24090 1510 24110 2890
rect 24010 1500 24110 1510
rect 21980 1480 24110 1500
rect 25780 2900 27910 2930
rect 25780 2670 25810 2900
rect 25850 2860 25890 2900
rect 27810 2890 27910 2900
rect 27810 2860 27850 2890
rect 25850 2840 27850 2860
rect 25850 2670 25870 2840
rect 25970 2746 25986 2780
rect 26020 2746 26036 2780
rect 26170 2746 26186 2780
rect 26220 2746 26236 2780
rect 26483 2739 26499 2773
rect 26533 2739 26549 2773
rect 26675 2739 26691 2773
rect 26725 2739 26741 2773
rect 26867 2739 26883 2773
rect 26917 2739 26933 2773
rect 27059 2739 27075 2773
rect 27109 2739 27125 2773
rect 27251 2739 27267 2773
rect 27301 2739 27317 2773
rect 27443 2739 27459 2773
rect 27493 2739 27509 2773
rect 27650 2746 27666 2780
rect 27700 2746 27716 2780
rect 25780 2540 25800 2670
rect 25860 2540 25870 2670
rect 25780 1520 25810 2540
rect 25850 1570 25870 2540
rect 25942 2696 25976 2712
rect 25942 1704 25976 1720
rect 26030 2696 26064 2712
rect 26142 2696 26176 2712
rect 26142 2504 26176 2520
rect 26230 2696 26264 2712
rect 26230 2504 26264 2520
rect 26355 2689 26389 2705
rect 26170 2436 26186 2470
rect 26220 2436 26236 2470
rect 26030 1704 26064 1720
rect 26355 1697 26389 1713
rect 26451 2689 26485 2705
rect 26451 1697 26485 1713
rect 26547 2689 26581 2705
rect 26547 1697 26581 1713
rect 26643 2689 26677 2705
rect 26643 1697 26677 1713
rect 26739 2689 26773 2705
rect 26739 1697 26773 1713
rect 26835 2689 26869 2705
rect 26835 1697 26869 1713
rect 26931 2689 26965 2705
rect 26931 1697 26965 1713
rect 27027 2689 27061 2705
rect 27027 1697 27061 1713
rect 27123 2689 27157 2705
rect 27123 1697 27157 1713
rect 27219 2689 27253 2705
rect 27219 1697 27253 1713
rect 27315 2689 27349 2705
rect 27315 1697 27349 1713
rect 27411 2689 27445 2705
rect 27411 1697 27445 1713
rect 27507 2689 27541 2705
rect 27507 1697 27541 1713
rect 27622 2696 27656 2712
rect 27622 1704 27656 1720
rect 27710 2696 27744 2712
rect 27710 1704 27744 1720
rect 25970 1636 25986 1670
rect 26020 1636 26036 1670
rect 26387 1629 26403 1663
rect 26437 1629 26453 1663
rect 26579 1629 26595 1663
rect 26629 1629 26645 1663
rect 26771 1629 26787 1663
rect 26821 1629 26837 1663
rect 26963 1629 26979 1663
rect 27013 1629 27029 1663
rect 27155 1629 27171 1663
rect 27205 1629 27221 1663
rect 27347 1629 27363 1663
rect 27397 1629 27413 1663
rect 27650 1636 27666 1670
rect 27700 1636 27716 1670
rect 27830 1570 27850 2840
rect 25850 1540 27850 1570
rect 25850 1520 25890 1540
rect 25780 1500 25890 1520
rect 27810 1510 27850 1540
rect 27890 1510 27910 2890
rect 27810 1500 27910 1510
rect 25780 1480 27910 1500
<< viali >>
rect 4977 27391 5011 27425
rect 5069 27391 5103 27425
rect 5161 27391 5195 27425
rect 5253 27391 5287 27425
rect 5345 27391 5379 27425
rect 5437 27391 5471 27425
rect 5529 27391 5563 27425
rect 5621 27391 5655 27425
rect 5713 27391 5747 27425
rect 5805 27391 5839 27425
rect 5897 27391 5931 27425
rect 5989 27391 6023 27425
rect 6081 27391 6115 27425
rect 6173 27391 6207 27425
rect 6265 27391 6299 27425
rect 6357 27391 6391 27425
rect 6449 27391 6483 27425
rect 6541 27391 6575 27425
rect 6633 27391 6667 27425
rect 6725 27391 6759 27425
rect 6817 27391 6851 27425
rect 6909 27391 6943 27425
rect 7001 27391 7035 27425
rect 7093 27391 7127 27425
rect 7185 27391 7219 27425
rect 7277 27391 7311 27425
rect 7369 27391 7403 27425
rect 7461 27391 7495 27425
rect 7553 27391 7587 27425
rect 7645 27391 7679 27425
rect 7737 27391 7771 27425
rect 7829 27391 7863 27425
rect 7921 27391 7955 27425
rect 8013 27391 8047 27425
rect 8105 27391 8139 27425
rect 8197 27391 8231 27425
rect 8289 27391 8323 27425
rect 8381 27391 8415 27425
rect 8473 27391 8507 27425
rect 8565 27391 8599 27425
rect 8657 27391 8691 27425
rect 8749 27391 8783 27425
rect 8841 27391 8875 27425
rect 8933 27391 8967 27425
rect 9025 27391 9059 27425
rect 9117 27391 9151 27425
rect 9209 27391 9243 27425
rect 9301 27391 9335 27425
rect 9393 27391 9427 27425
rect 9485 27391 9519 27425
rect 9577 27391 9611 27425
rect 9669 27391 9703 27425
rect 9761 27391 9795 27425
rect 9853 27391 9887 27425
rect 9945 27391 9979 27425
rect 10037 27391 10071 27425
rect 10129 27391 10163 27425
rect 10221 27391 10255 27425
rect 10313 27391 10347 27425
rect 10405 27391 10439 27425
rect 10497 27391 10531 27425
rect 10589 27391 10623 27425
rect 10681 27391 10715 27425
rect 10773 27391 10807 27425
rect 10865 27391 10899 27425
rect 10957 27391 10991 27425
rect 11049 27391 11083 27425
rect 11141 27391 11175 27425
rect 11233 27391 11267 27425
rect 11325 27391 11359 27425
rect 11417 27391 11451 27425
rect 11509 27391 11543 27425
rect 11601 27391 11635 27425
rect 11693 27391 11727 27425
rect 11785 27391 11819 27425
rect 11877 27391 11911 27425
rect 11969 27391 12003 27425
rect 12061 27391 12095 27425
rect 12153 27391 12187 27425
rect 12245 27391 12279 27425
rect 12337 27391 12371 27425
rect 12429 27391 12463 27425
rect 12521 27391 12555 27425
rect 12613 27391 12647 27425
rect 12705 27391 12739 27425
rect 12797 27391 12831 27425
rect 12889 27391 12923 27425
rect 12981 27391 13015 27425
rect 13073 27391 13107 27425
rect 13165 27391 13199 27425
rect 13257 27391 13291 27425
rect 13349 27391 13383 27425
rect 13441 27391 13475 27425
rect 13533 27391 13567 27425
rect 13625 27391 13659 27425
rect 13717 27391 13751 27425
rect 13809 27391 13843 27425
rect 13901 27391 13935 27425
rect 13993 27391 14027 27425
rect 14085 27391 14119 27425
rect 14177 27391 14211 27425
rect 14269 27391 14303 27425
rect 14361 27391 14395 27425
rect 14453 27391 14487 27425
rect 14545 27391 14579 27425
rect 14637 27391 14671 27425
rect 14729 27391 14763 27425
rect 14821 27391 14855 27425
rect 14913 27391 14947 27425
rect 15005 27391 15039 27425
rect 15097 27391 15131 27425
rect 15189 27391 15223 27425
rect 15281 27391 15315 27425
rect 15373 27391 15407 27425
rect 15465 27391 15499 27425
rect 15557 27391 15591 27425
rect 15649 27391 15683 27425
rect 15741 27391 15775 27425
rect 15833 27391 15867 27425
rect 15925 27391 15959 27425
rect 16017 27391 16051 27425
rect 16109 27391 16143 27425
rect 16201 27391 16235 27425
rect 16293 27391 16327 27425
rect 16385 27391 16419 27425
rect 16477 27391 16511 27425
rect 16569 27391 16603 27425
rect 16661 27391 16695 27425
rect 16753 27391 16787 27425
rect 16845 27391 16879 27425
rect 16937 27391 16971 27425
rect 17029 27391 17063 27425
rect 17121 27391 17155 27425
rect 17213 27391 17247 27425
rect 17305 27391 17339 27425
rect 17397 27391 17431 27425
rect 17489 27391 17523 27425
rect 17581 27391 17615 27425
rect 17673 27391 17707 27425
rect 17765 27391 17799 27425
rect 17857 27391 17891 27425
rect 17949 27391 17983 27425
rect 18041 27391 18075 27425
rect 18133 27391 18167 27425
rect 18225 27391 18259 27425
rect 18317 27391 18351 27425
rect 18409 27391 18443 27425
rect 18501 27391 18535 27425
rect 18593 27391 18627 27425
rect 18685 27391 18719 27425
rect 18777 27391 18811 27425
rect 18869 27391 18903 27425
rect 18961 27391 18995 27425
rect 19053 27391 19087 27425
rect 19145 27391 19179 27425
rect 19237 27391 19271 27425
rect 19329 27391 19363 27425
rect 19421 27391 19455 27425
rect 19513 27391 19547 27425
rect 19605 27391 19639 27425
rect 19697 27391 19731 27425
rect 19789 27391 19823 27425
rect 19881 27391 19915 27425
rect 19973 27391 20007 27425
rect 20065 27391 20099 27425
rect 20157 27391 20191 27425
rect 5897 27221 5931 27255
rect 5805 26958 5835 26983
rect 5835 26958 5839 26983
rect 5805 26949 5839 26958
rect 10129 27159 10137 27187
rect 10137 27159 10163 27187
rect 10129 27153 10163 27159
rect 10313 26965 10347 26983
rect 10313 26949 10341 26965
rect 10341 26949 10347 26965
rect 18869 27221 18903 27255
rect 18777 26958 18807 26983
rect 18807 26958 18811 26983
rect 18777 26949 18811 26958
rect 4977 26847 5011 26881
rect 5069 26847 5103 26881
rect 5161 26847 5195 26881
rect 5253 26847 5287 26881
rect 5345 26847 5379 26881
rect 5437 26847 5471 26881
rect 5529 26847 5563 26881
rect 5621 26847 5655 26881
rect 5713 26847 5747 26881
rect 5805 26847 5839 26881
rect 5897 26847 5931 26881
rect 5989 26847 6023 26881
rect 6081 26847 6115 26881
rect 6173 26847 6207 26881
rect 6265 26847 6299 26881
rect 6357 26847 6391 26881
rect 6449 26847 6483 26881
rect 6541 26847 6575 26881
rect 6633 26847 6667 26881
rect 6725 26847 6759 26881
rect 6817 26847 6851 26881
rect 6909 26847 6943 26881
rect 7001 26847 7035 26881
rect 7093 26847 7127 26881
rect 7185 26847 7219 26881
rect 7277 26847 7311 26881
rect 7369 26847 7403 26881
rect 7461 26847 7495 26881
rect 7553 26847 7587 26881
rect 7645 26847 7679 26881
rect 7737 26847 7771 26881
rect 7829 26847 7863 26881
rect 7921 26847 7955 26881
rect 8013 26847 8047 26881
rect 8105 26847 8139 26881
rect 8197 26847 8231 26881
rect 8289 26847 8323 26881
rect 8381 26847 8415 26881
rect 8473 26847 8507 26881
rect 8565 26847 8599 26881
rect 8657 26847 8691 26881
rect 8749 26847 8783 26881
rect 8841 26847 8875 26881
rect 8933 26847 8967 26881
rect 9025 26847 9059 26881
rect 9117 26847 9151 26881
rect 9209 26847 9243 26881
rect 9301 26847 9335 26881
rect 9393 26847 9427 26881
rect 9485 26847 9519 26881
rect 9577 26847 9611 26881
rect 9669 26847 9703 26881
rect 9761 26847 9795 26881
rect 9853 26847 9887 26881
rect 9945 26847 9979 26881
rect 10037 26847 10071 26881
rect 10129 26847 10163 26881
rect 10221 26847 10255 26881
rect 10313 26847 10347 26881
rect 10405 26847 10439 26881
rect 10497 26847 10531 26881
rect 10589 26847 10623 26881
rect 10681 26847 10715 26881
rect 10773 26847 10807 26881
rect 10865 26847 10899 26881
rect 10957 26847 10991 26881
rect 11049 26847 11083 26881
rect 11141 26847 11175 26881
rect 11233 26847 11267 26881
rect 11325 26847 11359 26881
rect 11417 26847 11451 26881
rect 11509 26847 11543 26881
rect 11601 26847 11635 26881
rect 11693 26847 11727 26881
rect 11785 26847 11819 26881
rect 11877 26847 11911 26881
rect 11969 26847 12003 26881
rect 12061 26847 12095 26881
rect 12153 26847 12187 26881
rect 12245 26847 12279 26881
rect 12337 26847 12371 26881
rect 12429 26847 12463 26881
rect 12521 26847 12555 26881
rect 12613 26847 12647 26881
rect 12705 26847 12739 26881
rect 12797 26847 12831 26881
rect 12889 26847 12923 26881
rect 12981 26847 13015 26881
rect 13073 26847 13107 26881
rect 13165 26847 13199 26881
rect 13257 26847 13291 26881
rect 13349 26847 13383 26881
rect 13441 26847 13475 26881
rect 13533 26847 13567 26881
rect 13625 26847 13659 26881
rect 13717 26847 13751 26881
rect 13809 26847 13843 26881
rect 13901 26847 13935 26881
rect 13993 26847 14027 26881
rect 14085 26847 14119 26881
rect 14177 26847 14211 26881
rect 14269 26847 14303 26881
rect 14361 26847 14395 26881
rect 14453 26847 14487 26881
rect 14545 26847 14579 26881
rect 14637 26847 14671 26881
rect 14729 26847 14763 26881
rect 14821 26847 14855 26881
rect 14913 26847 14947 26881
rect 15005 26847 15039 26881
rect 15097 26847 15131 26881
rect 15189 26847 15223 26881
rect 15281 26847 15315 26881
rect 15373 26847 15407 26881
rect 15465 26847 15499 26881
rect 15557 26847 15591 26881
rect 15649 26847 15683 26881
rect 15741 26847 15775 26881
rect 15833 26847 15867 26881
rect 15925 26847 15959 26881
rect 16017 26847 16051 26881
rect 16109 26847 16143 26881
rect 16201 26847 16235 26881
rect 16293 26847 16327 26881
rect 16385 26847 16419 26881
rect 16477 26847 16511 26881
rect 16569 26847 16603 26881
rect 16661 26847 16695 26881
rect 16753 26847 16787 26881
rect 16845 26847 16879 26881
rect 16937 26847 16971 26881
rect 17029 26847 17063 26881
rect 17121 26847 17155 26881
rect 17213 26847 17247 26881
rect 17305 26847 17339 26881
rect 17397 26847 17431 26881
rect 17489 26847 17523 26881
rect 17581 26847 17615 26881
rect 17673 26847 17707 26881
rect 17765 26847 17799 26881
rect 17857 26847 17891 26881
rect 17949 26847 17983 26881
rect 18041 26847 18075 26881
rect 18133 26847 18167 26881
rect 18225 26847 18259 26881
rect 18317 26847 18351 26881
rect 18409 26847 18443 26881
rect 18501 26847 18535 26881
rect 18593 26847 18627 26881
rect 18685 26847 18719 26881
rect 18777 26847 18811 26881
rect 18869 26847 18903 26881
rect 18961 26847 18995 26881
rect 19053 26847 19087 26881
rect 19145 26847 19179 26881
rect 19237 26847 19271 26881
rect 19329 26847 19363 26881
rect 19421 26847 19455 26881
rect 19513 26847 19547 26881
rect 19605 26847 19639 26881
rect 19697 26847 19731 26881
rect 19789 26847 19823 26881
rect 19881 26847 19915 26881
rect 19973 26847 20007 26881
rect 20065 26847 20099 26881
rect 20157 26847 20191 26881
rect 4977 26303 5011 26337
rect 5069 26303 5103 26337
rect 5161 26303 5195 26337
rect 5253 26303 5287 26337
rect 5345 26303 5379 26337
rect 5437 26303 5471 26337
rect 5529 26303 5563 26337
rect 5621 26303 5655 26337
rect 5713 26303 5747 26337
rect 5805 26303 5839 26337
rect 5897 26303 5931 26337
rect 5989 26303 6023 26337
rect 6081 26303 6115 26337
rect 6173 26303 6207 26337
rect 6265 26303 6299 26337
rect 6357 26303 6391 26337
rect 6449 26303 6483 26337
rect 6541 26303 6575 26337
rect 6633 26303 6667 26337
rect 6725 26303 6759 26337
rect 6817 26303 6851 26337
rect 6909 26303 6943 26337
rect 7001 26303 7035 26337
rect 7093 26303 7127 26337
rect 7185 26303 7219 26337
rect 7277 26303 7311 26337
rect 7369 26303 7403 26337
rect 7461 26303 7495 26337
rect 7553 26303 7587 26337
rect 7645 26303 7679 26337
rect 7737 26303 7771 26337
rect 7829 26303 7863 26337
rect 7921 26303 7955 26337
rect 8013 26303 8047 26337
rect 8105 26303 8139 26337
rect 8197 26303 8231 26337
rect 8289 26303 8323 26337
rect 8381 26303 8415 26337
rect 8473 26303 8507 26337
rect 8565 26303 8599 26337
rect 8657 26303 8691 26337
rect 8749 26303 8783 26337
rect 8841 26303 8875 26337
rect 8933 26303 8967 26337
rect 9025 26303 9059 26337
rect 9117 26303 9151 26337
rect 9209 26303 9243 26337
rect 9301 26303 9335 26337
rect 9393 26303 9427 26337
rect 9485 26303 9519 26337
rect 9577 26303 9611 26337
rect 9669 26303 9703 26337
rect 9761 26303 9795 26337
rect 9853 26303 9887 26337
rect 9945 26303 9979 26337
rect 10037 26303 10071 26337
rect 10129 26303 10163 26337
rect 10221 26303 10255 26337
rect 10313 26303 10347 26337
rect 10405 26303 10439 26337
rect 10497 26303 10531 26337
rect 10589 26303 10623 26337
rect 10681 26303 10715 26337
rect 10773 26303 10807 26337
rect 10865 26303 10899 26337
rect 10957 26303 10991 26337
rect 11049 26303 11083 26337
rect 11141 26303 11175 26337
rect 11233 26303 11267 26337
rect 11325 26303 11359 26337
rect 11417 26303 11451 26337
rect 11509 26303 11543 26337
rect 11601 26303 11635 26337
rect 11693 26303 11727 26337
rect 11785 26303 11819 26337
rect 11877 26303 11911 26337
rect 11969 26303 12003 26337
rect 12061 26303 12095 26337
rect 12153 26303 12187 26337
rect 12245 26303 12279 26337
rect 12337 26303 12371 26337
rect 12429 26303 12463 26337
rect 12521 26303 12555 26337
rect 12613 26303 12647 26337
rect 12705 26303 12739 26337
rect 12797 26303 12831 26337
rect 12889 26303 12923 26337
rect 12981 26303 13015 26337
rect 13073 26303 13107 26337
rect 13165 26303 13199 26337
rect 13257 26303 13291 26337
rect 13349 26303 13383 26337
rect 13441 26303 13475 26337
rect 13533 26303 13567 26337
rect 13625 26303 13659 26337
rect 13717 26303 13751 26337
rect 13809 26303 13843 26337
rect 13901 26303 13935 26337
rect 13993 26303 14027 26337
rect 14085 26303 14119 26337
rect 14177 26303 14211 26337
rect 14269 26303 14303 26337
rect 14361 26303 14395 26337
rect 14453 26303 14487 26337
rect 14545 26303 14579 26337
rect 14637 26303 14671 26337
rect 14729 26303 14763 26337
rect 14821 26303 14855 26337
rect 14913 26303 14947 26337
rect 15005 26303 15039 26337
rect 15097 26303 15131 26337
rect 15189 26303 15223 26337
rect 15281 26303 15315 26337
rect 15373 26303 15407 26337
rect 15465 26303 15499 26337
rect 15557 26303 15591 26337
rect 15649 26303 15683 26337
rect 15741 26303 15775 26337
rect 15833 26303 15867 26337
rect 15925 26303 15959 26337
rect 16017 26303 16051 26337
rect 16109 26303 16143 26337
rect 16201 26303 16235 26337
rect 16293 26303 16327 26337
rect 16385 26303 16419 26337
rect 16477 26303 16511 26337
rect 16569 26303 16603 26337
rect 16661 26303 16695 26337
rect 16753 26303 16787 26337
rect 16845 26303 16879 26337
rect 16937 26303 16971 26337
rect 17029 26303 17063 26337
rect 17121 26303 17155 26337
rect 17213 26303 17247 26337
rect 17305 26303 17339 26337
rect 17397 26303 17431 26337
rect 17489 26303 17523 26337
rect 17581 26303 17615 26337
rect 17673 26303 17707 26337
rect 17765 26303 17799 26337
rect 17857 26303 17891 26337
rect 17949 26303 17983 26337
rect 18041 26303 18075 26337
rect 18133 26303 18167 26337
rect 18225 26303 18259 26337
rect 18317 26303 18351 26337
rect 18409 26303 18443 26337
rect 18501 26303 18535 26337
rect 18593 26303 18627 26337
rect 18685 26303 18719 26337
rect 18777 26303 18811 26337
rect 18869 26303 18903 26337
rect 18961 26303 18995 26337
rect 19053 26303 19087 26337
rect 19145 26303 19179 26337
rect 19237 26303 19271 26337
rect 19329 26303 19363 26337
rect 19421 26303 19455 26337
rect 19513 26303 19547 26337
rect 19605 26303 19639 26337
rect 19697 26303 19731 26337
rect 19789 26303 19823 26337
rect 19881 26303 19915 26337
rect 19973 26303 20007 26337
rect 20065 26303 20099 26337
rect 20157 26303 20191 26337
rect 4977 25759 5011 25793
rect 5069 25759 5103 25793
rect 5161 25759 5195 25793
rect 5253 25759 5287 25793
rect 5345 25759 5379 25793
rect 5437 25759 5471 25793
rect 5529 25759 5563 25793
rect 5621 25759 5655 25793
rect 5713 25759 5747 25793
rect 5805 25759 5839 25793
rect 5897 25759 5931 25793
rect 5989 25759 6023 25793
rect 6081 25759 6115 25793
rect 6173 25759 6207 25793
rect 6265 25759 6299 25793
rect 6357 25759 6391 25793
rect 6449 25759 6483 25793
rect 6541 25759 6575 25793
rect 6633 25759 6667 25793
rect 6725 25759 6759 25793
rect 6817 25759 6851 25793
rect 6909 25759 6943 25793
rect 7001 25759 7035 25793
rect 7093 25759 7127 25793
rect 7185 25759 7219 25793
rect 7277 25759 7311 25793
rect 7369 25759 7403 25793
rect 7461 25759 7495 25793
rect 7553 25759 7587 25793
rect 7645 25759 7679 25793
rect 7737 25759 7771 25793
rect 7829 25759 7863 25793
rect 7921 25759 7955 25793
rect 8013 25759 8047 25793
rect 8105 25759 8139 25793
rect 8197 25759 8231 25793
rect 8289 25759 8323 25793
rect 8381 25759 8415 25793
rect 8473 25759 8507 25793
rect 8565 25759 8599 25793
rect 8657 25759 8691 25793
rect 8749 25759 8783 25793
rect 8841 25759 8875 25793
rect 8933 25759 8967 25793
rect 9025 25759 9059 25793
rect 9117 25759 9151 25793
rect 9209 25759 9243 25793
rect 9301 25759 9335 25793
rect 9393 25759 9427 25793
rect 9485 25759 9519 25793
rect 9577 25759 9611 25793
rect 9669 25759 9703 25793
rect 9761 25759 9795 25793
rect 9853 25759 9887 25793
rect 9945 25759 9979 25793
rect 10037 25759 10071 25793
rect 10129 25759 10163 25793
rect 10221 25759 10255 25793
rect 10313 25759 10347 25793
rect 10405 25759 10439 25793
rect 10497 25759 10531 25793
rect 10589 25759 10623 25793
rect 10681 25759 10715 25793
rect 10773 25759 10807 25793
rect 10865 25759 10899 25793
rect 10957 25759 10991 25793
rect 11049 25759 11083 25793
rect 11141 25759 11175 25793
rect 11233 25759 11267 25793
rect 11325 25759 11359 25793
rect 11417 25759 11451 25793
rect 11509 25759 11543 25793
rect 11601 25759 11635 25793
rect 11693 25759 11727 25793
rect 11785 25759 11819 25793
rect 11877 25759 11911 25793
rect 11969 25759 12003 25793
rect 12061 25759 12095 25793
rect 12153 25759 12187 25793
rect 12245 25759 12279 25793
rect 12337 25759 12371 25793
rect 12429 25759 12463 25793
rect 12521 25759 12555 25793
rect 12613 25759 12647 25793
rect 12705 25759 12739 25793
rect 12797 25759 12831 25793
rect 12889 25759 12923 25793
rect 12981 25759 13015 25793
rect 13073 25759 13107 25793
rect 13165 25759 13199 25793
rect 13257 25759 13291 25793
rect 13349 25759 13383 25793
rect 13441 25759 13475 25793
rect 13533 25759 13567 25793
rect 13625 25759 13659 25793
rect 13717 25759 13751 25793
rect 13809 25759 13843 25793
rect 13901 25759 13935 25793
rect 13993 25759 14027 25793
rect 14085 25759 14119 25793
rect 14177 25759 14211 25793
rect 14269 25759 14303 25793
rect 14361 25759 14395 25793
rect 14453 25759 14487 25793
rect 14545 25759 14579 25793
rect 14637 25759 14671 25793
rect 14729 25759 14763 25793
rect 14821 25759 14855 25793
rect 14913 25759 14947 25793
rect 15005 25759 15039 25793
rect 15097 25759 15131 25793
rect 15189 25759 15223 25793
rect 15281 25759 15315 25793
rect 15373 25759 15407 25793
rect 15465 25759 15499 25793
rect 15557 25759 15591 25793
rect 15649 25759 15683 25793
rect 15741 25759 15775 25793
rect 15833 25759 15867 25793
rect 15925 25759 15959 25793
rect 16017 25759 16051 25793
rect 16109 25759 16143 25793
rect 16201 25759 16235 25793
rect 16293 25759 16327 25793
rect 16385 25759 16419 25793
rect 16477 25759 16511 25793
rect 16569 25759 16603 25793
rect 16661 25759 16695 25793
rect 16753 25759 16787 25793
rect 16845 25759 16879 25793
rect 16937 25759 16971 25793
rect 17029 25759 17063 25793
rect 17121 25759 17155 25793
rect 17213 25759 17247 25793
rect 17305 25759 17339 25793
rect 17397 25759 17431 25793
rect 17489 25759 17523 25793
rect 17581 25759 17615 25793
rect 17673 25759 17707 25793
rect 17765 25759 17799 25793
rect 17857 25759 17891 25793
rect 17949 25759 17983 25793
rect 18041 25759 18075 25793
rect 18133 25759 18167 25793
rect 18225 25759 18259 25793
rect 18317 25759 18351 25793
rect 18409 25759 18443 25793
rect 18501 25759 18535 25793
rect 18593 25759 18627 25793
rect 18685 25759 18719 25793
rect 18777 25759 18811 25793
rect 18869 25759 18903 25793
rect 18961 25759 18995 25793
rect 19053 25759 19087 25793
rect 19145 25759 19179 25793
rect 19237 25759 19271 25793
rect 19329 25759 19363 25793
rect 19421 25759 19455 25793
rect 19513 25759 19547 25793
rect 19605 25759 19639 25793
rect 19697 25759 19731 25793
rect 19789 25759 19823 25793
rect 19881 25759 19915 25793
rect 19973 25759 20007 25793
rect 20065 25759 20099 25793
rect 20157 25759 20191 25793
rect 4977 25215 5011 25249
rect 5069 25215 5103 25249
rect 5161 25215 5195 25249
rect 5253 25215 5287 25249
rect 5345 25215 5379 25249
rect 5437 25215 5471 25249
rect 5529 25215 5563 25249
rect 5621 25215 5655 25249
rect 5713 25215 5747 25249
rect 5805 25215 5839 25249
rect 5897 25215 5931 25249
rect 5989 25215 6023 25249
rect 6081 25215 6115 25249
rect 6173 25215 6207 25249
rect 6265 25215 6299 25249
rect 6357 25215 6391 25249
rect 6449 25215 6483 25249
rect 6541 25215 6575 25249
rect 6633 25215 6667 25249
rect 6725 25215 6759 25249
rect 6817 25215 6851 25249
rect 6909 25215 6943 25249
rect 7001 25215 7035 25249
rect 7093 25215 7127 25249
rect 7185 25215 7219 25249
rect 7277 25215 7311 25249
rect 7369 25215 7403 25249
rect 7461 25215 7495 25249
rect 7553 25215 7587 25249
rect 7645 25215 7679 25249
rect 7737 25215 7771 25249
rect 7829 25215 7863 25249
rect 7921 25215 7955 25249
rect 8013 25215 8047 25249
rect 8105 25215 8139 25249
rect 8197 25215 8231 25249
rect 8289 25215 8323 25249
rect 8381 25215 8415 25249
rect 8473 25215 8507 25249
rect 8565 25215 8599 25249
rect 8657 25215 8691 25249
rect 8749 25215 8783 25249
rect 8841 25215 8875 25249
rect 8933 25215 8967 25249
rect 9025 25215 9059 25249
rect 9117 25215 9151 25249
rect 9209 25215 9243 25249
rect 9301 25215 9335 25249
rect 9393 25215 9427 25249
rect 9485 25215 9519 25249
rect 9577 25215 9611 25249
rect 9669 25215 9703 25249
rect 9761 25215 9795 25249
rect 9853 25215 9887 25249
rect 9945 25215 9979 25249
rect 10037 25215 10071 25249
rect 10129 25215 10163 25249
rect 10221 25215 10255 25249
rect 10313 25215 10347 25249
rect 10405 25215 10439 25249
rect 10497 25215 10531 25249
rect 10589 25215 10623 25249
rect 10681 25215 10715 25249
rect 10773 25215 10807 25249
rect 10865 25215 10899 25249
rect 10957 25215 10991 25249
rect 11049 25215 11083 25249
rect 11141 25215 11175 25249
rect 11233 25215 11267 25249
rect 11325 25215 11359 25249
rect 11417 25215 11451 25249
rect 11509 25215 11543 25249
rect 11601 25215 11635 25249
rect 11693 25215 11727 25249
rect 11785 25215 11819 25249
rect 11877 25215 11911 25249
rect 11969 25215 12003 25249
rect 12061 25215 12095 25249
rect 12153 25215 12187 25249
rect 12245 25215 12279 25249
rect 12337 25215 12371 25249
rect 12429 25215 12463 25249
rect 12521 25215 12555 25249
rect 12613 25215 12647 25249
rect 12705 25215 12739 25249
rect 12797 25215 12831 25249
rect 12889 25215 12923 25249
rect 12981 25215 13015 25249
rect 13073 25215 13107 25249
rect 13165 25215 13199 25249
rect 13257 25215 13291 25249
rect 13349 25215 13383 25249
rect 13441 25215 13475 25249
rect 13533 25215 13567 25249
rect 13625 25215 13659 25249
rect 13717 25215 13751 25249
rect 13809 25215 13843 25249
rect 13901 25215 13935 25249
rect 13993 25215 14027 25249
rect 14085 25215 14119 25249
rect 14177 25215 14211 25249
rect 14269 25215 14303 25249
rect 14361 25215 14395 25249
rect 14453 25215 14487 25249
rect 14545 25215 14579 25249
rect 14637 25215 14671 25249
rect 14729 25215 14763 25249
rect 14821 25215 14855 25249
rect 14913 25215 14947 25249
rect 15005 25215 15039 25249
rect 15097 25215 15131 25249
rect 15189 25215 15223 25249
rect 15281 25215 15315 25249
rect 15373 25215 15407 25249
rect 15465 25215 15499 25249
rect 15557 25215 15591 25249
rect 15649 25215 15683 25249
rect 15741 25215 15775 25249
rect 15833 25215 15867 25249
rect 15925 25215 15959 25249
rect 16017 25215 16051 25249
rect 16109 25215 16143 25249
rect 16201 25215 16235 25249
rect 16293 25215 16327 25249
rect 16385 25215 16419 25249
rect 16477 25215 16511 25249
rect 16569 25215 16603 25249
rect 16661 25215 16695 25249
rect 16753 25215 16787 25249
rect 16845 25215 16879 25249
rect 16937 25215 16971 25249
rect 17029 25215 17063 25249
rect 17121 25215 17155 25249
rect 17213 25215 17247 25249
rect 17305 25215 17339 25249
rect 17397 25215 17431 25249
rect 17489 25215 17523 25249
rect 17581 25215 17615 25249
rect 17673 25215 17707 25249
rect 17765 25215 17799 25249
rect 17857 25215 17891 25249
rect 17949 25215 17983 25249
rect 18041 25215 18075 25249
rect 18133 25215 18167 25249
rect 18225 25215 18259 25249
rect 18317 25215 18351 25249
rect 18409 25215 18443 25249
rect 18501 25215 18535 25249
rect 18593 25215 18627 25249
rect 18685 25215 18719 25249
rect 18777 25215 18811 25249
rect 18869 25215 18903 25249
rect 18961 25215 18995 25249
rect 19053 25215 19087 25249
rect 19145 25215 19179 25249
rect 19237 25215 19271 25249
rect 19329 25215 19363 25249
rect 19421 25215 19455 25249
rect 19513 25215 19547 25249
rect 19605 25215 19639 25249
rect 19697 25215 19731 25249
rect 19789 25215 19823 25249
rect 19881 25215 19915 25249
rect 19973 25215 20007 25249
rect 20065 25215 20099 25249
rect 20157 25215 20191 25249
rect 4977 24671 5011 24705
rect 5069 24671 5103 24705
rect 5161 24671 5195 24705
rect 5253 24671 5287 24705
rect 5345 24671 5379 24705
rect 5437 24671 5471 24705
rect 5529 24671 5563 24705
rect 5621 24671 5655 24705
rect 5713 24671 5747 24705
rect 5805 24671 5839 24705
rect 5897 24671 5931 24705
rect 5989 24671 6023 24705
rect 6081 24671 6115 24705
rect 6173 24671 6207 24705
rect 6265 24671 6299 24705
rect 6357 24671 6391 24705
rect 6449 24671 6483 24705
rect 6541 24671 6575 24705
rect 6633 24671 6667 24705
rect 6725 24671 6759 24705
rect 6817 24671 6851 24705
rect 6909 24671 6943 24705
rect 7001 24671 7035 24705
rect 7093 24671 7127 24705
rect 7185 24671 7219 24705
rect 7277 24671 7311 24705
rect 7369 24671 7403 24705
rect 7461 24671 7495 24705
rect 7553 24671 7587 24705
rect 7645 24671 7679 24705
rect 7737 24671 7771 24705
rect 7829 24671 7863 24705
rect 7921 24671 7955 24705
rect 8013 24671 8047 24705
rect 8105 24671 8139 24705
rect 8197 24671 8231 24705
rect 8289 24671 8323 24705
rect 8381 24671 8415 24705
rect 8473 24671 8507 24705
rect 8565 24671 8599 24705
rect 8657 24671 8691 24705
rect 8749 24671 8783 24705
rect 8841 24671 8875 24705
rect 8933 24671 8967 24705
rect 9025 24671 9059 24705
rect 9117 24671 9151 24705
rect 9209 24671 9243 24705
rect 9301 24671 9335 24705
rect 9393 24671 9427 24705
rect 9485 24671 9519 24705
rect 9577 24671 9611 24705
rect 9669 24671 9703 24705
rect 9761 24671 9795 24705
rect 9853 24671 9887 24705
rect 9945 24671 9979 24705
rect 10037 24671 10071 24705
rect 10129 24671 10163 24705
rect 10221 24671 10255 24705
rect 10313 24671 10347 24705
rect 10405 24671 10439 24705
rect 10497 24671 10531 24705
rect 10589 24671 10623 24705
rect 10681 24671 10715 24705
rect 10773 24671 10807 24705
rect 10865 24671 10899 24705
rect 10957 24671 10991 24705
rect 11049 24671 11083 24705
rect 11141 24671 11175 24705
rect 11233 24671 11267 24705
rect 11325 24671 11359 24705
rect 11417 24671 11451 24705
rect 11509 24671 11543 24705
rect 11601 24671 11635 24705
rect 11693 24671 11727 24705
rect 11785 24671 11819 24705
rect 11877 24671 11911 24705
rect 11969 24671 12003 24705
rect 12061 24671 12095 24705
rect 12153 24671 12187 24705
rect 12245 24671 12279 24705
rect 12337 24671 12371 24705
rect 12429 24671 12463 24705
rect 12521 24671 12555 24705
rect 12613 24671 12647 24705
rect 12705 24671 12739 24705
rect 12797 24671 12831 24705
rect 12889 24671 12923 24705
rect 12981 24671 13015 24705
rect 13073 24671 13107 24705
rect 13165 24671 13199 24705
rect 13257 24671 13291 24705
rect 13349 24671 13383 24705
rect 13441 24671 13475 24705
rect 13533 24671 13567 24705
rect 13625 24671 13659 24705
rect 13717 24671 13751 24705
rect 13809 24671 13843 24705
rect 13901 24671 13935 24705
rect 13993 24671 14027 24705
rect 14085 24671 14119 24705
rect 14177 24671 14211 24705
rect 14269 24671 14303 24705
rect 14361 24671 14395 24705
rect 14453 24671 14487 24705
rect 14545 24671 14579 24705
rect 14637 24671 14671 24705
rect 14729 24671 14763 24705
rect 14821 24671 14855 24705
rect 14913 24671 14947 24705
rect 15005 24671 15039 24705
rect 15097 24671 15131 24705
rect 15189 24671 15223 24705
rect 15281 24671 15315 24705
rect 15373 24671 15407 24705
rect 15465 24671 15499 24705
rect 15557 24671 15591 24705
rect 15649 24671 15683 24705
rect 15741 24671 15775 24705
rect 15833 24671 15867 24705
rect 15925 24671 15959 24705
rect 16017 24671 16051 24705
rect 16109 24671 16143 24705
rect 16201 24671 16235 24705
rect 16293 24671 16327 24705
rect 16385 24671 16419 24705
rect 16477 24671 16511 24705
rect 16569 24671 16603 24705
rect 16661 24671 16695 24705
rect 16753 24671 16787 24705
rect 16845 24671 16879 24705
rect 16937 24671 16971 24705
rect 17029 24671 17063 24705
rect 17121 24671 17155 24705
rect 17213 24671 17247 24705
rect 17305 24671 17339 24705
rect 17397 24671 17431 24705
rect 17489 24671 17523 24705
rect 17581 24671 17615 24705
rect 17673 24671 17707 24705
rect 17765 24671 17799 24705
rect 17857 24671 17891 24705
rect 17949 24671 17983 24705
rect 18041 24671 18075 24705
rect 18133 24671 18167 24705
rect 18225 24671 18259 24705
rect 18317 24671 18351 24705
rect 18409 24671 18443 24705
rect 18501 24671 18535 24705
rect 18593 24671 18627 24705
rect 18685 24671 18719 24705
rect 18777 24671 18811 24705
rect 18869 24671 18903 24705
rect 18961 24671 18995 24705
rect 19053 24671 19087 24705
rect 19145 24671 19179 24705
rect 19237 24671 19271 24705
rect 19329 24671 19363 24705
rect 19421 24671 19455 24705
rect 19513 24671 19547 24705
rect 19605 24671 19639 24705
rect 19697 24671 19731 24705
rect 19789 24671 19823 24705
rect 19881 24671 19915 24705
rect 19973 24671 20007 24705
rect 20065 24671 20099 24705
rect 20157 24671 20191 24705
rect 4977 24127 5011 24161
rect 5069 24127 5103 24161
rect 5161 24127 5195 24161
rect 5253 24127 5287 24161
rect 5345 24127 5379 24161
rect 5437 24127 5471 24161
rect 5529 24127 5563 24161
rect 5621 24127 5655 24161
rect 5713 24127 5747 24161
rect 5805 24127 5839 24161
rect 5897 24127 5931 24161
rect 5989 24127 6023 24161
rect 6081 24127 6115 24161
rect 6173 24127 6207 24161
rect 6265 24127 6299 24161
rect 6357 24127 6391 24161
rect 6449 24127 6483 24161
rect 6541 24127 6575 24161
rect 6633 24127 6667 24161
rect 6725 24127 6759 24161
rect 6817 24127 6851 24161
rect 6909 24127 6943 24161
rect 7001 24127 7035 24161
rect 7093 24127 7127 24161
rect 7185 24127 7219 24161
rect 7277 24127 7311 24161
rect 7369 24127 7403 24161
rect 7461 24127 7495 24161
rect 7553 24127 7587 24161
rect 7645 24127 7679 24161
rect 7737 24127 7771 24161
rect 7829 24127 7863 24161
rect 7921 24127 7955 24161
rect 8013 24127 8047 24161
rect 8105 24127 8139 24161
rect 8197 24127 8231 24161
rect 8289 24127 8323 24161
rect 8381 24127 8415 24161
rect 8473 24127 8507 24161
rect 8565 24127 8599 24161
rect 8657 24127 8691 24161
rect 8749 24127 8783 24161
rect 8841 24127 8875 24161
rect 8933 24127 8967 24161
rect 9025 24127 9059 24161
rect 9117 24127 9151 24161
rect 9209 24127 9243 24161
rect 9301 24127 9335 24161
rect 9393 24127 9427 24161
rect 9485 24127 9519 24161
rect 9577 24127 9611 24161
rect 9669 24127 9703 24161
rect 9761 24127 9795 24161
rect 9853 24127 9887 24161
rect 9945 24127 9979 24161
rect 10037 24127 10071 24161
rect 10129 24127 10163 24161
rect 10221 24127 10255 24161
rect 10313 24127 10347 24161
rect 10405 24127 10439 24161
rect 10497 24127 10531 24161
rect 10589 24127 10623 24161
rect 10681 24127 10715 24161
rect 10773 24127 10807 24161
rect 10865 24127 10899 24161
rect 10957 24127 10991 24161
rect 11049 24127 11083 24161
rect 11141 24127 11175 24161
rect 11233 24127 11267 24161
rect 11325 24127 11359 24161
rect 11417 24127 11451 24161
rect 11509 24127 11543 24161
rect 11601 24127 11635 24161
rect 11693 24127 11727 24161
rect 11785 24127 11819 24161
rect 11877 24127 11911 24161
rect 11969 24127 12003 24161
rect 12061 24127 12095 24161
rect 12153 24127 12187 24161
rect 12245 24127 12279 24161
rect 12337 24127 12371 24161
rect 12429 24127 12463 24161
rect 12521 24127 12555 24161
rect 12613 24127 12647 24161
rect 12705 24127 12739 24161
rect 12797 24127 12831 24161
rect 12889 24127 12923 24161
rect 12981 24127 13015 24161
rect 13073 24127 13107 24161
rect 13165 24127 13199 24161
rect 13257 24127 13291 24161
rect 13349 24127 13383 24161
rect 13441 24127 13475 24161
rect 13533 24127 13567 24161
rect 13625 24127 13659 24161
rect 13717 24127 13751 24161
rect 13809 24127 13843 24161
rect 13901 24127 13935 24161
rect 13993 24127 14027 24161
rect 14085 24127 14119 24161
rect 14177 24127 14211 24161
rect 14269 24127 14303 24161
rect 14361 24127 14395 24161
rect 14453 24127 14487 24161
rect 14545 24127 14579 24161
rect 14637 24127 14671 24161
rect 14729 24127 14763 24161
rect 14821 24127 14855 24161
rect 14913 24127 14947 24161
rect 15005 24127 15039 24161
rect 15097 24127 15131 24161
rect 15189 24127 15223 24161
rect 15281 24127 15315 24161
rect 15373 24127 15407 24161
rect 15465 24127 15499 24161
rect 15557 24127 15591 24161
rect 15649 24127 15683 24161
rect 15741 24127 15775 24161
rect 15833 24127 15867 24161
rect 15925 24127 15959 24161
rect 16017 24127 16051 24161
rect 16109 24127 16143 24161
rect 16201 24127 16235 24161
rect 16293 24127 16327 24161
rect 16385 24127 16419 24161
rect 16477 24127 16511 24161
rect 16569 24127 16603 24161
rect 16661 24127 16695 24161
rect 16753 24127 16787 24161
rect 16845 24127 16879 24161
rect 16937 24127 16971 24161
rect 17029 24127 17063 24161
rect 17121 24127 17155 24161
rect 17213 24127 17247 24161
rect 17305 24127 17339 24161
rect 17397 24127 17431 24161
rect 17489 24127 17523 24161
rect 17581 24127 17615 24161
rect 17673 24127 17707 24161
rect 17765 24127 17799 24161
rect 17857 24127 17891 24161
rect 17949 24127 17983 24161
rect 18041 24127 18075 24161
rect 18133 24127 18167 24161
rect 18225 24127 18259 24161
rect 18317 24127 18351 24161
rect 18409 24127 18443 24161
rect 18501 24127 18535 24161
rect 18593 24127 18627 24161
rect 18685 24127 18719 24161
rect 18777 24127 18811 24161
rect 18869 24127 18903 24161
rect 18961 24127 18995 24161
rect 19053 24127 19087 24161
rect 19145 24127 19179 24161
rect 19237 24127 19271 24161
rect 19329 24127 19363 24161
rect 19421 24127 19455 24161
rect 19513 24127 19547 24161
rect 19605 24127 19639 24161
rect 19697 24127 19731 24161
rect 19789 24127 19823 24161
rect 19881 24127 19915 24161
rect 19973 24127 20007 24161
rect 20065 24127 20099 24161
rect 20157 24127 20191 24161
rect 4977 23583 5011 23617
rect 5069 23583 5103 23617
rect 5161 23583 5195 23617
rect 5253 23583 5287 23617
rect 5345 23583 5379 23617
rect 5437 23583 5471 23617
rect 5529 23583 5563 23617
rect 5621 23583 5655 23617
rect 5713 23583 5747 23617
rect 5805 23583 5839 23617
rect 5897 23583 5931 23617
rect 5989 23583 6023 23617
rect 6081 23583 6115 23617
rect 6173 23583 6207 23617
rect 6265 23583 6299 23617
rect 6357 23583 6391 23617
rect 6449 23583 6483 23617
rect 6541 23583 6575 23617
rect 6633 23583 6667 23617
rect 6725 23583 6759 23617
rect 6817 23583 6851 23617
rect 6909 23583 6943 23617
rect 7001 23583 7035 23617
rect 7093 23583 7127 23617
rect 7185 23583 7219 23617
rect 7277 23583 7311 23617
rect 7369 23583 7403 23617
rect 7461 23583 7495 23617
rect 7553 23583 7587 23617
rect 7645 23583 7679 23617
rect 7737 23583 7771 23617
rect 7829 23583 7863 23617
rect 7921 23583 7955 23617
rect 8013 23583 8047 23617
rect 8105 23583 8139 23617
rect 8197 23583 8231 23617
rect 8289 23583 8323 23617
rect 8381 23583 8415 23617
rect 8473 23583 8507 23617
rect 8565 23583 8599 23617
rect 8657 23583 8691 23617
rect 8749 23583 8783 23617
rect 8841 23583 8875 23617
rect 8933 23583 8967 23617
rect 9025 23583 9059 23617
rect 9117 23583 9151 23617
rect 9209 23583 9243 23617
rect 9301 23583 9335 23617
rect 9393 23583 9427 23617
rect 9485 23583 9519 23617
rect 9577 23583 9611 23617
rect 9669 23583 9703 23617
rect 9761 23583 9795 23617
rect 9853 23583 9887 23617
rect 9945 23583 9979 23617
rect 10037 23583 10071 23617
rect 10129 23583 10163 23617
rect 10221 23583 10255 23617
rect 10313 23583 10347 23617
rect 10405 23583 10439 23617
rect 10497 23583 10531 23617
rect 10589 23583 10623 23617
rect 10681 23583 10715 23617
rect 10773 23583 10807 23617
rect 10865 23583 10899 23617
rect 10957 23583 10991 23617
rect 11049 23583 11083 23617
rect 11141 23583 11175 23617
rect 11233 23583 11267 23617
rect 11325 23583 11359 23617
rect 11417 23583 11451 23617
rect 11509 23583 11543 23617
rect 11601 23583 11635 23617
rect 11693 23583 11727 23617
rect 11785 23583 11819 23617
rect 11877 23583 11911 23617
rect 11969 23583 12003 23617
rect 12061 23583 12095 23617
rect 12153 23583 12187 23617
rect 12245 23583 12279 23617
rect 12337 23583 12371 23617
rect 12429 23583 12463 23617
rect 12521 23583 12555 23617
rect 12613 23583 12647 23617
rect 12705 23583 12739 23617
rect 12797 23583 12831 23617
rect 12889 23583 12923 23617
rect 12981 23583 13015 23617
rect 13073 23583 13107 23617
rect 13165 23583 13199 23617
rect 13257 23583 13291 23617
rect 13349 23583 13383 23617
rect 13441 23583 13475 23617
rect 13533 23583 13567 23617
rect 13625 23583 13659 23617
rect 13717 23583 13751 23617
rect 13809 23583 13843 23617
rect 13901 23583 13935 23617
rect 13993 23583 14027 23617
rect 14085 23583 14119 23617
rect 14177 23583 14211 23617
rect 14269 23583 14303 23617
rect 14361 23583 14395 23617
rect 14453 23583 14487 23617
rect 14545 23583 14579 23617
rect 14637 23583 14671 23617
rect 14729 23583 14763 23617
rect 14821 23583 14855 23617
rect 14913 23583 14947 23617
rect 15005 23583 15039 23617
rect 15097 23583 15131 23617
rect 15189 23583 15223 23617
rect 15281 23583 15315 23617
rect 15373 23583 15407 23617
rect 15465 23583 15499 23617
rect 15557 23583 15591 23617
rect 15649 23583 15683 23617
rect 15741 23583 15775 23617
rect 15833 23583 15867 23617
rect 15925 23583 15959 23617
rect 16017 23583 16051 23617
rect 16109 23583 16143 23617
rect 16201 23583 16235 23617
rect 16293 23583 16327 23617
rect 16385 23583 16419 23617
rect 16477 23583 16511 23617
rect 16569 23583 16603 23617
rect 16661 23583 16695 23617
rect 16753 23583 16787 23617
rect 16845 23583 16879 23617
rect 16937 23583 16971 23617
rect 17029 23583 17063 23617
rect 17121 23583 17155 23617
rect 17213 23583 17247 23617
rect 17305 23583 17339 23617
rect 17397 23583 17431 23617
rect 17489 23583 17523 23617
rect 17581 23583 17615 23617
rect 17673 23583 17707 23617
rect 17765 23583 17799 23617
rect 17857 23583 17891 23617
rect 17949 23583 17983 23617
rect 18041 23583 18075 23617
rect 18133 23583 18167 23617
rect 18225 23583 18259 23617
rect 18317 23583 18351 23617
rect 18409 23583 18443 23617
rect 18501 23583 18535 23617
rect 18593 23583 18627 23617
rect 18685 23583 18719 23617
rect 18777 23583 18811 23617
rect 18869 23583 18903 23617
rect 18961 23583 18995 23617
rect 19053 23583 19087 23617
rect 19145 23583 19179 23617
rect 19237 23583 19271 23617
rect 19329 23583 19363 23617
rect 19421 23583 19455 23617
rect 19513 23583 19547 23617
rect 19605 23583 19639 23617
rect 19697 23583 19731 23617
rect 19789 23583 19823 23617
rect 19881 23583 19915 23617
rect 19973 23583 20007 23617
rect 20065 23583 20099 23617
rect 20157 23583 20191 23617
rect 4977 23039 5011 23073
rect 5069 23039 5103 23073
rect 5161 23039 5195 23073
rect 5253 23039 5287 23073
rect 5345 23039 5379 23073
rect 5437 23039 5471 23073
rect 5529 23039 5563 23073
rect 5621 23039 5655 23073
rect 5713 23039 5747 23073
rect 5805 23039 5839 23073
rect 5897 23039 5931 23073
rect 5989 23039 6023 23073
rect 6081 23039 6115 23073
rect 6173 23039 6207 23073
rect 6265 23039 6299 23073
rect 6357 23039 6391 23073
rect 6449 23039 6483 23073
rect 6541 23039 6575 23073
rect 6633 23039 6667 23073
rect 6725 23039 6759 23073
rect 6817 23039 6851 23073
rect 6909 23039 6943 23073
rect 7001 23039 7035 23073
rect 7093 23039 7127 23073
rect 7185 23039 7219 23073
rect 7277 23039 7311 23073
rect 7369 23039 7403 23073
rect 7461 23039 7495 23073
rect 7553 23039 7587 23073
rect 7645 23039 7679 23073
rect 7737 23039 7771 23073
rect 7829 23039 7863 23073
rect 7921 23039 7955 23073
rect 8013 23039 8047 23073
rect 8105 23039 8139 23073
rect 8197 23039 8231 23073
rect 8289 23039 8323 23073
rect 8381 23039 8415 23073
rect 8473 23039 8507 23073
rect 8565 23039 8599 23073
rect 8657 23039 8691 23073
rect 8749 23039 8783 23073
rect 8841 23039 8875 23073
rect 8933 23039 8967 23073
rect 9025 23039 9059 23073
rect 9117 23039 9151 23073
rect 9209 23039 9243 23073
rect 9301 23039 9335 23073
rect 9393 23039 9427 23073
rect 9485 23039 9519 23073
rect 9577 23039 9611 23073
rect 9669 23039 9703 23073
rect 9761 23039 9795 23073
rect 9853 23039 9887 23073
rect 9945 23039 9979 23073
rect 10037 23039 10071 23073
rect 10129 23039 10163 23073
rect 10221 23039 10255 23073
rect 10313 23039 10347 23073
rect 10405 23039 10439 23073
rect 10497 23039 10531 23073
rect 10589 23039 10623 23073
rect 10681 23039 10715 23073
rect 10773 23039 10807 23073
rect 10865 23039 10899 23073
rect 10957 23039 10991 23073
rect 11049 23039 11083 23073
rect 11141 23039 11175 23073
rect 11233 23039 11267 23073
rect 11325 23039 11359 23073
rect 11417 23039 11451 23073
rect 11509 23039 11543 23073
rect 11601 23039 11635 23073
rect 11693 23039 11727 23073
rect 11785 23039 11819 23073
rect 11877 23039 11911 23073
rect 11969 23039 12003 23073
rect 12061 23039 12095 23073
rect 12153 23039 12187 23073
rect 12245 23039 12279 23073
rect 12337 23039 12371 23073
rect 12429 23039 12463 23073
rect 12521 23039 12555 23073
rect 12613 23039 12647 23073
rect 12705 23039 12739 23073
rect 12797 23039 12831 23073
rect 12889 23039 12923 23073
rect 12981 23039 13015 23073
rect 13073 23039 13107 23073
rect 13165 23039 13199 23073
rect 13257 23039 13291 23073
rect 13349 23039 13383 23073
rect 13441 23039 13475 23073
rect 13533 23039 13567 23073
rect 13625 23039 13659 23073
rect 13717 23039 13751 23073
rect 13809 23039 13843 23073
rect 13901 23039 13935 23073
rect 13993 23039 14027 23073
rect 14085 23039 14119 23073
rect 14177 23039 14211 23073
rect 14269 23039 14303 23073
rect 14361 23039 14395 23073
rect 14453 23039 14487 23073
rect 14545 23039 14579 23073
rect 14637 23039 14671 23073
rect 14729 23039 14763 23073
rect 14821 23039 14855 23073
rect 14913 23039 14947 23073
rect 15005 23039 15039 23073
rect 15097 23039 15131 23073
rect 15189 23039 15223 23073
rect 15281 23039 15315 23073
rect 15373 23039 15407 23073
rect 15465 23039 15499 23073
rect 15557 23039 15591 23073
rect 15649 23039 15683 23073
rect 15741 23039 15775 23073
rect 15833 23039 15867 23073
rect 15925 23039 15959 23073
rect 16017 23039 16051 23073
rect 16109 23039 16143 23073
rect 16201 23039 16235 23073
rect 16293 23039 16327 23073
rect 16385 23039 16419 23073
rect 16477 23039 16511 23073
rect 16569 23039 16603 23073
rect 16661 23039 16695 23073
rect 16753 23039 16787 23073
rect 16845 23039 16879 23073
rect 16937 23039 16971 23073
rect 17029 23039 17063 23073
rect 17121 23039 17155 23073
rect 17213 23039 17247 23073
rect 17305 23039 17339 23073
rect 17397 23039 17431 23073
rect 17489 23039 17523 23073
rect 17581 23039 17615 23073
rect 17673 23039 17707 23073
rect 17765 23039 17799 23073
rect 17857 23039 17891 23073
rect 17949 23039 17983 23073
rect 18041 23039 18075 23073
rect 18133 23039 18167 23073
rect 18225 23039 18259 23073
rect 18317 23039 18351 23073
rect 18409 23039 18443 23073
rect 18501 23039 18535 23073
rect 18593 23039 18627 23073
rect 18685 23039 18719 23073
rect 18777 23039 18811 23073
rect 18869 23039 18903 23073
rect 18961 23039 18995 23073
rect 19053 23039 19087 23073
rect 19145 23039 19179 23073
rect 19237 23039 19271 23073
rect 19329 23039 19363 23073
rect 19421 23039 19455 23073
rect 19513 23039 19547 23073
rect 19605 23039 19639 23073
rect 19697 23039 19731 23073
rect 19789 23039 19823 23073
rect 19881 23039 19915 23073
rect 19973 23039 20007 23073
rect 20065 23039 20099 23073
rect 20157 23039 20191 23073
rect 4977 22495 5011 22529
rect 5069 22495 5103 22529
rect 5161 22495 5195 22529
rect 5253 22495 5287 22529
rect 5345 22495 5379 22529
rect 5437 22495 5471 22529
rect 5529 22495 5563 22529
rect 5621 22495 5655 22529
rect 5713 22495 5747 22529
rect 5805 22495 5839 22529
rect 5897 22495 5931 22529
rect 5989 22495 6023 22529
rect 6081 22495 6115 22529
rect 6173 22495 6207 22529
rect 6265 22495 6299 22529
rect 6357 22495 6391 22529
rect 6449 22495 6483 22529
rect 6541 22495 6575 22529
rect 6633 22495 6667 22529
rect 6725 22495 6759 22529
rect 6817 22495 6851 22529
rect 6909 22495 6943 22529
rect 7001 22495 7035 22529
rect 7093 22495 7127 22529
rect 7185 22495 7219 22529
rect 7277 22495 7311 22529
rect 7369 22495 7403 22529
rect 7461 22495 7495 22529
rect 7553 22495 7587 22529
rect 7645 22495 7679 22529
rect 7737 22495 7771 22529
rect 7829 22495 7863 22529
rect 7921 22495 7955 22529
rect 8013 22495 8047 22529
rect 8105 22495 8139 22529
rect 8197 22495 8231 22529
rect 8289 22495 8323 22529
rect 8381 22495 8415 22529
rect 8473 22495 8507 22529
rect 8565 22495 8599 22529
rect 8657 22495 8691 22529
rect 8749 22495 8783 22529
rect 8841 22495 8875 22529
rect 8933 22495 8967 22529
rect 9025 22495 9059 22529
rect 9117 22495 9151 22529
rect 9209 22495 9243 22529
rect 9301 22495 9335 22529
rect 9393 22495 9427 22529
rect 9485 22495 9519 22529
rect 9577 22495 9611 22529
rect 9669 22495 9703 22529
rect 9761 22495 9795 22529
rect 9853 22495 9887 22529
rect 9945 22495 9979 22529
rect 10037 22495 10071 22529
rect 10129 22495 10163 22529
rect 10221 22495 10255 22529
rect 10313 22495 10347 22529
rect 10405 22495 10439 22529
rect 10497 22495 10531 22529
rect 10589 22495 10623 22529
rect 10681 22495 10715 22529
rect 10773 22495 10807 22529
rect 10865 22495 10899 22529
rect 10957 22495 10991 22529
rect 11049 22495 11083 22529
rect 11141 22495 11175 22529
rect 11233 22495 11267 22529
rect 11325 22495 11359 22529
rect 11417 22495 11451 22529
rect 11509 22495 11543 22529
rect 11601 22495 11635 22529
rect 11693 22495 11727 22529
rect 11785 22495 11819 22529
rect 11877 22495 11911 22529
rect 11969 22495 12003 22529
rect 12061 22495 12095 22529
rect 12153 22495 12187 22529
rect 12245 22495 12279 22529
rect 12337 22495 12371 22529
rect 12429 22495 12463 22529
rect 12521 22495 12555 22529
rect 12613 22495 12647 22529
rect 12705 22495 12739 22529
rect 12797 22495 12831 22529
rect 12889 22495 12923 22529
rect 12981 22495 13015 22529
rect 13073 22495 13107 22529
rect 13165 22495 13199 22529
rect 13257 22495 13291 22529
rect 13349 22495 13383 22529
rect 13441 22495 13475 22529
rect 13533 22495 13567 22529
rect 13625 22495 13659 22529
rect 13717 22495 13751 22529
rect 13809 22495 13843 22529
rect 13901 22495 13935 22529
rect 13993 22495 14027 22529
rect 14085 22495 14119 22529
rect 14177 22495 14211 22529
rect 14269 22495 14303 22529
rect 14361 22495 14395 22529
rect 14453 22495 14487 22529
rect 14545 22495 14579 22529
rect 14637 22495 14671 22529
rect 14729 22495 14763 22529
rect 14821 22495 14855 22529
rect 14913 22495 14947 22529
rect 15005 22495 15039 22529
rect 15097 22495 15131 22529
rect 15189 22495 15223 22529
rect 15281 22495 15315 22529
rect 15373 22495 15407 22529
rect 15465 22495 15499 22529
rect 15557 22495 15591 22529
rect 15649 22495 15683 22529
rect 15741 22495 15775 22529
rect 15833 22495 15867 22529
rect 15925 22495 15959 22529
rect 16017 22495 16051 22529
rect 16109 22495 16143 22529
rect 16201 22495 16235 22529
rect 16293 22495 16327 22529
rect 16385 22495 16419 22529
rect 16477 22495 16511 22529
rect 16569 22495 16603 22529
rect 16661 22495 16695 22529
rect 16753 22495 16787 22529
rect 16845 22495 16879 22529
rect 16937 22495 16971 22529
rect 17029 22495 17063 22529
rect 17121 22495 17155 22529
rect 17213 22495 17247 22529
rect 17305 22495 17339 22529
rect 17397 22495 17431 22529
rect 17489 22495 17523 22529
rect 17581 22495 17615 22529
rect 17673 22495 17707 22529
rect 17765 22495 17799 22529
rect 17857 22495 17891 22529
rect 17949 22495 17983 22529
rect 18041 22495 18075 22529
rect 18133 22495 18167 22529
rect 18225 22495 18259 22529
rect 18317 22495 18351 22529
rect 18409 22495 18443 22529
rect 18501 22495 18535 22529
rect 18593 22495 18627 22529
rect 18685 22495 18719 22529
rect 18777 22495 18811 22529
rect 18869 22495 18903 22529
rect 18961 22495 18995 22529
rect 19053 22495 19087 22529
rect 19145 22495 19179 22529
rect 19237 22495 19271 22529
rect 19329 22495 19363 22529
rect 19421 22495 19455 22529
rect 19513 22495 19547 22529
rect 19605 22495 19639 22529
rect 19697 22495 19731 22529
rect 19789 22495 19823 22529
rect 19881 22495 19915 22529
rect 19973 22495 20007 22529
rect 20065 22495 20099 22529
rect 20157 22495 20191 22529
rect 4977 21951 5011 21985
rect 5069 21951 5103 21985
rect 5161 21951 5195 21985
rect 5253 21951 5287 21985
rect 5345 21951 5379 21985
rect 5437 21951 5471 21985
rect 5529 21951 5563 21985
rect 5621 21951 5655 21985
rect 5713 21951 5747 21985
rect 5805 21951 5839 21985
rect 5897 21951 5931 21985
rect 5989 21951 6023 21985
rect 6081 21951 6115 21985
rect 6173 21951 6207 21985
rect 6265 21951 6299 21985
rect 6357 21951 6391 21985
rect 6449 21951 6483 21985
rect 6541 21951 6575 21985
rect 6633 21951 6667 21985
rect 6725 21951 6759 21985
rect 6817 21951 6851 21985
rect 6909 21951 6943 21985
rect 7001 21951 7035 21985
rect 7093 21951 7127 21985
rect 7185 21951 7219 21985
rect 7277 21951 7311 21985
rect 7369 21951 7403 21985
rect 7461 21951 7495 21985
rect 7553 21951 7587 21985
rect 7645 21951 7679 21985
rect 7737 21951 7771 21985
rect 7829 21951 7863 21985
rect 7921 21951 7955 21985
rect 8013 21951 8047 21985
rect 8105 21951 8139 21985
rect 8197 21951 8231 21985
rect 8289 21951 8323 21985
rect 8381 21951 8415 21985
rect 8473 21951 8507 21985
rect 8565 21951 8599 21985
rect 8657 21951 8691 21985
rect 8749 21951 8783 21985
rect 8841 21951 8875 21985
rect 8933 21951 8967 21985
rect 9025 21951 9059 21985
rect 9117 21951 9151 21985
rect 9209 21951 9243 21985
rect 9301 21951 9335 21985
rect 9393 21951 9427 21985
rect 9485 21951 9519 21985
rect 9577 21951 9611 21985
rect 9669 21951 9703 21985
rect 9761 21951 9795 21985
rect 9853 21951 9887 21985
rect 9945 21951 9979 21985
rect 10037 21951 10071 21985
rect 10129 21951 10163 21985
rect 10221 21951 10255 21985
rect 10313 21951 10347 21985
rect 10405 21951 10439 21985
rect 10497 21951 10531 21985
rect 10589 21951 10623 21985
rect 10681 21951 10715 21985
rect 10773 21951 10807 21985
rect 10865 21951 10899 21985
rect 10957 21951 10991 21985
rect 11049 21951 11083 21985
rect 11141 21951 11175 21985
rect 11233 21951 11267 21985
rect 11325 21951 11359 21985
rect 11417 21951 11451 21985
rect 11509 21951 11543 21985
rect 11601 21951 11635 21985
rect 11693 21951 11727 21985
rect 11785 21951 11819 21985
rect 11877 21951 11911 21985
rect 11969 21951 12003 21985
rect 12061 21951 12095 21985
rect 12153 21951 12187 21985
rect 12245 21951 12279 21985
rect 12337 21951 12371 21985
rect 12429 21951 12463 21985
rect 12521 21951 12555 21985
rect 12613 21951 12647 21985
rect 12705 21951 12739 21985
rect 12797 21951 12831 21985
rect 12889 21951 12923 21985
rect 12981 21951 13015 21985
rect 13073 21951 13107 21985
rect 13165 21951 13199 21985
rect 13257 21951 13291 21985
rect 13349 21951 13383 21985
rect 13441 21951 13475 21985
rect 13533 21951 13567 21985
rect 13625 21951 13659 21985
rect 13717 21951 13751 21985
rect 13809 21951 13843 21985
rect 13901 21951 13935 21985
rect 13993 21951 14027 21985
rect 14085 21951 14119 21985
rect 14177 21951 14211 21985
rect 14269 21951 14303 21985
rect 14361 21951 14395 21985
rect 14453 21951 14487 21985
rect 14545 21951 14579 21985
rect 14637 21951 14671 21985
rect 14729 21951 14763 21985
rect 14821 21951 14855 21985
rect 14913 21951 14947 21985
rect 15005 21951 15039 21985
rect 15097 21951 15131 21985
rect 15189 21951 15223 21985
rect 15281 21951 15315 21985
rect 15373 21951 15407 21985
rect 15465 21951 15499 21985
rect 15557 21951 15591 21985
rect 15649 21951 15683 21985
rect 15741 21951 15775 21985
rect 15833 21951 15867 21985
rect 15925 21951 15959 21985
rect 16017 21951 16051 21985
rect 16109 21951 16143 21985
rect 16201 21951 16235 21985
rect 16293 21951 16327 21985
rect 16385 21951 16419 21985
rect 16477 21951 16511 21985
rect 16569 21951 16603 21985
rect 16661 21951 16695 21985
rect 16753 21951 16787 21985
rect 16845 21951 16879 21985
rect 16937 21951 16971 21985
rect 17029 21951 17063 21985
rect 17121 21951 17155 21985
rect 17213 21951 17247 21985
rect 17305 21951 17339 21985
rect 17397 21951 17431 21985
rect 17489 21951 17523 21985
rect 17581 21951 17615 21985
rect 17673 21951 17707 21985
rect 17765 21951 17799 21985
rect 17857 21951 17891 21985
rect 17949 21951 17983 21985
rect 18041 21951 18075 21985
rect 18133 21951 18167 21985
rect 18225 21951 18259 21985
rect 18317 21951 18351 21985
rect 18409 21951 18443 21985
rect 18501 21951 18535 21985
rect 18593 21951 18627 21985
rect 18685 21951 18719 21985
rect 18777 21951 18811 21985
rect 18869 21951 18903 21985
rect 18961 21951 18995 21985
rect 19053 21951 19087 21985
rect 19145 21951 19179 21985
rect 19237 21951 19271 21985
rect 19329 21951 19363 21985
rect 19421 21951 19455 21985
rect 19513 21951 19547 21985
rect 19605 21951 19639 21985
rect 19697 21951 19731 21985
rect 19789 21951 19823 21985
rect 19881 21951 19915 21985
rect 19973 21951 20007 21985
rect 20065 21951 20099 21985
rect 20157 21951 20191 21985
rect 4977 21407 5011 21441
rect 5069 21407 5103 21441
rect 5161 21407 5195 21441
rect 5253 21407 5287 21441
rect 5345 21407 5379 21441
rect 5437 21407 5471 21441
rect 5529 21407 5563 21441
rect 5621 21407 5655 21441
rect 5713 21407 5747 21441
rect 5805 21407 5839 21441
rect 5897 21407 5931 21441
rect 5989 21407 6023 21441
rect 6081 21407 6115 21441
rect 6173 21407 6207 21441
rect 6265 21407 6299 21441
rect 6357 21407 6391 21441
rect 6449 21407 6483 21441
rect 6541 21407 6575 21441
rect 6633 21407 6667 21441
rect 6725 21407 6759 21441
rect 6817 21407 6851 21441
rect 6909 21407 6943 21441
rect 7001 21407 7035 21441
rect 7093 21407 7127 21441
rect 7185 21407 7219 21441
rect 7277 21407 7311 21441
rect 7369 21407 7403 21441
rect 7461 21407 7495 21441
rect 7553 21407 7587 21441
rect 7645 21407 7679 21441
rect 7737 21407 7771 21441
rect 7829 21407 7863 21441
rect 7921 21407 7955 21441
rect 8013 21407 8047 21441
rect 8105 21407 8139 21441
rect 8197 21407 8231 21441
rect 8289 21407 8323 21441
rect 8381 21407 8415 21441
rect 8473 21407 8507 21441
rect 8565 21407 8599 21441
rect 8657 21407 8691 21441
rect 8749 21407 8783 21441
rect 8841 21407 8875 21441
rect 8933 21407 8967 21441
rect 9025 21407 9059 21441
rect 9117 21407 9151 21441
rect 9209 21407 9243 21441
rect 9301 21407 9335 21441
rect 9393 21407 9427 21441
rect 9485 21407 9519 21441
rect 9577 21407 9611 21441
rect 9669 21407 9703 21441
rect 9761 21407 9795 21441
rect 9853 21407 9887 21441
rect 9945 21407 9979 21441
rect 10037 21407 10071 21441
rect 10129 21407 10163 21441
rect 10221 21407 10255 21441
rect 10313 21407 10347 21441
rect 10405 21407 10439 21441
rect 10497 21407 10531 21441
rect 10589 21407 10623 21441
rect 10681 21407 10715 21441
rect 10773 21407 10807 21441
rect 10865 21407 10899 21441
rect 10957 21407 10991 21441
rect 11049 21407 11083 21441
rect 11141 21407 11175 21441
rect 11233 21407 11267 21441
rect 11325 21407 11359 21441
rect 11417 21407 11451 21441
rect 11509 21407 11543 21441
rect 11601 21407 11635 21441
rect 11693 21407 11727 21441
rect 11785 21407 11819 21441
rect 11877 21407 11911 21441
rect 11969 21407 12003 21441
rect 12061 21407 12095 21441
rect 12153 21407 12187 21441
rect 12245 21407 12279 21441
rect 12337 21407 12371 21441
rect 12429 21407 12463 21441
rect 12521 21407 12555 21441
rect 12613 21407 12647 21441
rect 12705 21407 12739 21441
rect 12797 21407 12831 21441
rect 12889 21407 12923 21441
rect 12981 21407 13015 21441
rect 13073 21407 13107 21441
rect 13165 21407 13199 21441
rect 13257 21407 13291 21441
rect 13349 21407 13383 21441
rect 13441 21407 13475 21441
rect 13533 21407 13567 21441
rect 13625 21407 13659 21441
rect 13717 21407 13751 21441
rect 13809 21407 13843 21441
rect 13901 21407 13935 21441
rect 13993 21407 14027 21441
rect 14085 21407 14119 21441
rect 14177 21407 14211 21441
rect 14269 21407 14303 21441
rect 14361 21407 14395 21441
rect 14453 21407 14487 21441
rect 14545 21407 14579 21441
rect 14637 21407 14671 21441
rect 14729 21407 14763 21441
rect 14821 21407 14855 21441
rect 14913 21407 14947 21441
rect 15005 21407 15039 21441
rect 15097 21407 15131 21441
rect 15189 21407 15223 21441
rect 15281 21407 15315 21441
rect 15373 21407 15407 21441
rect 15465 21407 15499 21441
rect 15557 21407 15591 21441
rect 15649 21407 15683 21441
rect 15741 21407 15775 21441
rect 15833 21407 15867 21441
rect 15925 21407 15959 21441
rect 16017 21407 16051 21441
rect 16109 21407 16143 21441
rect 16201 21407 16235 21441
rect 16293 21407 16327 21441
rect 16385 21407 16419 21441
rect 16477 21407 16511 21441
rect 16569 21407 16603 21441
rect 16661 21407 16695 21441
rect 16753 21407 16787 21441
rect 16845 21407 16879 21441
rect 16937 21407 16971 21441
rect 17029 21407 17063 21441
rect 17121 21407 17155 21441
rect 17213 21407 17247 21441
rect 17305 21407 17339 21441
rect 17397 21407 17431 21441
rect 17489 21407 17523 21441
rect 17581 21407 17615 21441
rect 17673 21407 17707 21441
rect 17765 21407 17799 21441
rect 17857 21407 17891 21441
rect 17949 21407 17983 21441
rect 18041 21407 18075 21441
rect 18133 21407 18167 21441
rect 18225 21407 18259 21441
rect 18317 21407 18351 21441
rect 18409 21407 18443 21441
rect 18501 21407 18535 21441
rect 18593 21407 18627 21441
rect 18685 21407 18719 21441
rect 18777 21407 18811 21441
rect 18869 21407 18903 21441
rect 18961 21407 18995 21441
rect 19053 21407 19087 21441
rect 19145 21407 19179 21441
rect 19237 21407 19271 21441
rect 19329 21407 19363 21441
rect 19421 21407 19455 21441
rect 19513 21407 19547 21441
rect 19605 21407 19639 21441
rect 19697 21407 19731 21441
rect 19789 21407 19823 21441
rect 19881 21407 19915 21441
rect 19973 21407 20007 21441
rect 20065 21407 20099 21441
rect 20157 21407 20191 21441
rect 4977 20863 5011 20897
rect 5069 20863 5103 20897
rect 5161 20863 5195 20897
rect 5253 20863 5287 20897
rect 5345 20863 5379 20897
rect 5437 20863 5471 20897
rect 5529 20863 5563 20897
rect 5621 20863 5655 20897
rect 5713 20863 5747 20897
rect 5805 20863 5839 20897
rect 5897 20863 5931 20897
rect 5989 20863 6023 20897
rect 6081 20863 6115 20897
rect 6173 20863 6207 20897
rect 6265 20863 6299 20897
rect 6357 20863 6391 20897
rect 6449 20863 6483 20897
rect 6541 20863 6575 20897
rect 6633 20863 6667 20897
rect 6725 20863 6759 20897
rect 6817 20863 6851 20897
rect 6909 20863 6943 20897
rect 7001 20863 7035 20897
rect 7093 20863 7127 20897
rect 7185 20863 7219 20897
rect 7277 20863 7311 20897
rect 7369 20863 7403 20897
rect 7461 20863 7495 20897
rect 7553 20863 7587 20897
rect 7645 20863 7679 20897
rect 7737 20863 7771 20897
rect 7829 20863 7863 20897
rect 7921 20863 7955 20897
rect 8013 20863 8047 20897
rect 8105 20863 8139 20897
rect 8197 20863 8231 20897
rect 8289 20863 8323 20897
rect 8381 20863 8415 20897
rect 8473 20863 8507 20897
rect 8565 20863 8599 20897
rect 8657 20863 8691 20897
rect 8749 20863 8783 20897
rect 8841 20863 8875 20897
rect 8933 20863 8967 20897
rect 9025 20863 9059 20897
rect 9117 20863 9151 20897
rect 9209 20863 9243 20897
rect 9301 20863 9335 20897
rect 9393 20863 9427 20897
rect 9485 20863 9519 20897
rect 9577 20863 9611 20897
rect 9669 20863 9703 20897
rect 9761 20863 9795 20897
rect 9853 20863 9887 20897
rect 9945 20863 9979 20897
rect 10037 20863 10071 20897
rect 10129 20863 10163 20897
rect 10221 20863 10255 20897
rect 10313 20863 10347 20897
rect 10405 20863 10439 20897
rect 10497 20863 10531 20897
rect 10589 20863 10623 20897
rect 10681 20863 10715 20897
rect 10773 20863 10807 20897
rect 10865 20863 10899 20897
rect 10957 20863 10991 20897
rect 11049 20863 11083 20897
rect 11141 20863 11175 20897
rect 11233 20863 11267 20897
rect 11325 20863 11359 20897
rect 11417 20863 11451 20897
rect 11509 20863 11543 20897
rect 11601 20863 11635 20897
rect 11693 20863 11727 20897
rect 11785 20863 11819 20897
rect 11877 20863 11911 20897
rect 11969 20863 12003 20897
rect 12061 20863 12095 20897
rect 12153 20863 12187 20897
rect 12245 20863 12279 20897
rect 12337 20863 12371 20897
rect 12429 20863 12463 20897
rect 12521 20863 12555 20897
rect 12613 20863 12647 20897
rect 12705 20863 12739 20897
rect 12797 20863 12831 20897
rect 12889 20863 12923 20897
rect 12981 20863 13015 20897
rect 13073 20863 13107 20897
rect 13165 20863 13199 20897
rect 13257 20863 13291 20897
rect 13349 20863 13383 20897
rect 13441 20863 13475 20897
rect 13533 20863 13567 20897
rect 13625 20863 13659 20897
rect 13717 20863 13751 20897
rect 13809 20863 13843 20897
rect 13901 20863 13935 20897
rect 13993 20863 14027 20897
rect 14085 20863 14119 20897
rect 14177 20863 14211 20897
rect 14269 20863 14303 20897
rect 14361 20863 14395 20897
rect 14453 20863 14487 20897
rect 14545 20863 14579 20897
rect 14637 20863 14671 20897
rect 14729 20863 14763 20897
rect 14821 20863 14855 20897
rect 14913 20863 14947 20897
rect 15005 20863 15039 20897
rect 15097 20863 15131 20897
rect 15189 20863 15223 20897
rect 15281 20863 15315 20897
rect 15373 20863 15407 20897
rect 15465 20863 15499 20897
rect 15557 20863 15591 20897
rect 15649 20863 15683 20897
rect 15741 20863 15775 20897
rect 15833 20863 15867 20897
rect 15925 20863 15959 20897
rect 16017 20863 16051 20897
rect 16109 20863 16143 20897
rect 16201 20863 16235 20897
rect 16293 20863 16327 20897
rect 16385 20863 16419 20897
rect 16477 20863 16511 20897
rect 16569 20863 16603 20897
rect 16661 20863 16695 20897
rect 16753 20863 16787 20897
rect 16845 20863 16879 20897
rect 16937 20863 16971 20897
rect 17029 20863 17063 20897
rect 17121 20863 17155 20897
rect 17213 20863 17247 20897
rect 17305 20863 17339 20897
rect 17397 20863 17431 20897
rect 17489 20863 17523 20897
rect 17581 20863 17615 20897
rect 17673 20863 17707 20897
rect 17765 20863 17799 20897
rect 17857 20863 17891 20897
rect 17949 20863 17983 20897
rect 18041 20863 18075 20897
rect 18133 20863 18167 20897
rect 18225 20863 18259 20897
rect 18317 20863 18351 20897
rect 18409 20863 18443 20897
rect 18501 20863 18535 20897
rect 18593 20863 18627 20897
rect 18685 20863 18719 20897
rect 18777 20863 18811 20897
rect 18869 20863 18903 20897
rect 18961 20863 18995 20897
rect 19053 20863 19087 20897
rect 19145 20863 19179 20897
rect 19237 20863 19271 20897
rect 19329 20863 19363 20897
rect 19421 20863 19455 20897
rect 19513 20863 19547 20897
rect 19605 20863 19639 20897
rect 19697 20863 19731 20897
rect 19789 20863 19823 20897
rect 19881 20863 19915 20897
rect 19973 20863 20007 20897
rect 20065 20863 20099 20897
rect 20157 20863 20191 20897
rect 4977 20319 5011 20353
rect 5069 20319 5103 20353
rect 5161 20319 5195 20353
rect 5253 20319 5287 20353
rect 5345 20319 5379 20353
rect 5437 20319 5471 20353
rect 5529 20319 5563 20353
rect 5621 20319 5655 20353
rect 5713 20319 5747 20353
rect 5805 20319 5839 20353
rect 5897 20319 5931 20353
rect 5989 20319 6023 20353
rect 6081 20319 6115 20353
rect 6173 20319 6207 20353
rect 6265 20319 6299 20353
rect 6357 20319 6391 20353
rect 6449 20319 6483 20353
rect 6541 20319 6575 20353
rect 6633 20319 6667 20353
rect 6725 20319 6759 20353
rect 6817 20319 6851 20353
rect 6909 20319 6943 20353
rect 7001 20319 7035 20353
rect 7093 20319 7127 20353
rect 7185 20319 7219 20353
rect 7277 20319 7311 20353
rect 7369 20319 7403 20353
rect 7461 20319 7495 20353
rect 7553 20319 7587 20353
rect 7645 20319 7679 20353
rect 7737 20319 7771 20353
rect 7829 20319 7863 20353
rect 7921 20319 7955 20353
rect 8013 20319 8047 20353
rect 8105 20319 8139 20353
rect 8197 20319 8231 20353
rect 8289 20319 8323 20353
rect 8381 20319 8415 20353
rect 8473 20319 8507 20353
rect 8565 20319 8599 20353
rect 8657 20319 8691 20353
rect 8749 20319 8783 20353
rect 8841 20319 8875 20353
rect 8933 20319 8967 20353
rect 9025 20319 9059 20353
rect 9117 20319 9151 20353
rect 9209 20319 9243 20353
rect 9301 20319 9335 20353
rect 9393 20319 9427 20353
rect 9485 20319 9519 20353
rect 9577 20319 9611 20353
rect 9669 20319 9703 20353
rect 9761 20319 9795 20353
rect 9853 20319 9887 20353
rect 9945 20319 9979 20353
rect 10037 20319 10071 20353
rect 10129 20319 10163 20353
rect 10221 20319 10255 20353
rect 10313 20319 10347 20353
rect 10405 20319 10439 20353
rect 10497 20319 10531 20353
rect 10589 20319 10623 20353
rect 10681 20319 10715 20353
rect 10773 20319 10807 20353
rect 10865 20319 10899 20353
rect 10957 20319 10991 20353
rect 11049 20319 11083 20353
rect 11141 20319 11175 20353
rect 11233 20319 11267 20353
rect 11325 20319 11359 20353
rect 11417 20319 11451 20353
rect 11509 20319 11543 20353
rect 11601 20319 11635 20353
rect 11693 20319 11727 20353
rect 11785 20319 11819 20353
rect 11877 20319 11911 20353
rect 11969 20319 12003 20353
rect 12061 20319 12095 20353
rect 12153 20319 12187 20353
rect 12245 20319 12279 20353
rect 12337 20319 12371 20353
rect 12429 20319 12463 20353
rect 12521 20319 12555 20353
rect 12613 20319 12647 20353
rect 12705 20319 12739 20353
rect 12797 20319 12831 20353
rect 12889 20319 12923 20353
rect 12981 20319 13015 20353
rect 13073 20319 13107 20353
rect 13165 20319 13199 20353
rect 13257 20319 13291 20353
rect 13349 20319 13383 20353
rect 13441 20319 13475 20353
rect 13533 20319 13567 20353
rect 13625 20319 13659 20353
rect 13717 20319 13751 20353
rect 13809 20319 13843 20353
rect 13901 20319 13935 20353
rect 13993 20319 14027 20353
rect 14085 20319 14119 20353
rect 14177 20319 14211 20353
rect 14269 20319 14303 20353
rect 14361 20319 14395 20353
rect 14453 20319 14487 20353
rect 14545 20319 14579 20353
rect 14637 20319 14671 20353
rect 14729 20319 14763 20353
rect 14821 20319 14855 20353
rect 14913 20319 14947 20353
rect 15005 20319 15039 20353
rect 15097 20319 15131 20353
rect 15189 20319 15223 20353
rect 15281 20319 15315 20353
rect 15373 20319 15407 20353
rect 15465 20319 15499 20353
rect 15557 20319 15591 20353
rect 15649 20319 15683 20353
rect 15741 20319 15775 20353
rect 15833 20319 15867 20353
rect 15925 20319 15959 20353
rect 16017 20319 16051 20353
rect 16109 20319 16143 20353
rect 16201 20319 16235 20353
rect 16293 20319 16327 20353
rect 16385 20319 16419 20353
rect 16477 20319 16511 20353
rect 16569 20319 16603 20353
rect 16661 20319 16695 20353
rect 16753 20319 16787 20353
rect 16845 20319 16879 20353
rect 16937 20319 16971 20353
rect 17029 20319 17063 20353
rect 17121 20319 17155 20353
rect 17213 20319 17247 20353
rect 17305 20319 17339 20353
rect 17397 20319 17431 20353
rect 17489 20319 17523 20353
rect 17581 20319 17615 20353
rect 17673 20319 17707 20353
rect 17765 20319 17799 20353
rect 17857 20319 17891 20353
rect 17949 20319 17983 20353
rect 18041 20319 18075 20353
rect 18133 20319 18167 20353
rect 18225 20319 18259 20353
rect 18317 20319 18351 20353
rect 18409 20319 18443 20353
rect 18501 20319 18535 20353
rect 18593 20319 18627 20353
rect 18685 20319 18719 20353
rect 18777 20319 18811 20353
rect 18869 20319 18903 20353
rect 18961 20319 18995 20353
rect 19053 20319 19087 20353
rect 19145 20319 19179 20353
rect 19237 20319 19271 20353
rect 19329 20319 19363 20353
rect 19421 20319 19455 20353
rect 19513 20319 19547 20353
rect 19605 20319 19639 20353
rect 19697 20319 19731 20353
rect 19789 20319 19823 20353
rect 19881 20319 19915 20353
rect 19973 20319 20007 20353
rect 20065 20319 20099 20353
rect 20157 20319 20191 20353
rect 4977 19775 5011 19809
rect 5069 19775 5103 19809
rect 5161 19775 5195 19809
rect 5253 19775 5287 19809
rect 5345 19775 5379 19809
rect 5437 19775 5471 19809
rect 5529 19775 5563 19809
rect 5621 19775 5655 19809
rect 5713 19775 5747 19809
rect 5805 19775 5839 19809
rect 5897 19775 5931 19809
rect 5989 19775 6023 19809
rect 6081 19775 6115 19809
rect 6173 19775 6207 19809
rect 6265 19775 6299 19809
rect 6357 19775 6391 19809
rect 6449 19775 6483 19809
rect 6541 19775 6575 19809
rect 6633 19775 6667 19809
rect 6725 19775 6759 19809
rect 6817 19775 6851 19809
rect 6909 19775 6943 19809
rect 7001 19775 7035 19809
rect 7093 19775 7127 19809
rect 7185 19775 7219 19809
rect 7277 19775 7311 19809
rect 7369 19775 7403 19809
rect 7461 19775 7495 19809
rect 7553 19775 7587 19809
rect 7645 19775 7679 19809
rect 7737 19775 7771 19809
rect 7829 19775 7863 19809
rect 7921 19775 7955 19809
rect 8013 19775 8047 19809
rect 8105 19775 8139 19809
rect 8197 19775 8231 19809
rect 8289 19775 8323 19809
rect 8381 19775 8415 19809
rect 8473 19775 8507 19809
rect 8565 19775 8599 19809
rect 8657 19775 8691 19809
rect 8749 19775 8783 19809
rect 8841 19775 8875 19809
rect 8933 19775 8967 19809
rect 9025 19775 9059 19809
rect 9117 19775 9151 19809
rect 9209 19775 9243 19809
rect 9301 19775 9335 19809
rect 9393 19775 9427 19809
rect 9485 19775 9519 19809
rect 9577 19775 9611 19809
rect 9669 19775 9703 19809
rect 9761 19775 9795 19809
rect 9853 19775 9887 19809
rect 9945 19775 9979 19809
rect 10037 19775 10071 19809
rect 10129 19775 10163 19809
rect 10221 19775 10255 19809
rect 10313 19775 10347 19809
rect 10405 19775 10439 19809
rect 10497 19775 10531 19809
rect 10589 19775 10623 19809
rect 10681 19775 10715 19809
rect 10773 19775 10807 19809
rect 10865 19775 10899 19809
rect 10957 19775 10991 19809
rect 11049 19775 11083 19809
rect 11141 19775 11175 19809
rect 11233 19775 11267 19809
rect 11325 19775 11359 19809
rect 11417 19775 11451 19809
rect 11509 19775 11543 19809
rect 11601 19775 11635 19809
rect 11693 19775 11727 19809
rect 11785 19775 11819 19809
rect 11877 19775 11911 19809
rect 11969 19775 12003 19809
rect 12061 19775 12095 19809
rect 12153 19775 12187 19809
rect 12245 19775 12279 19809
rect 12337 19775 12371 19809
rect 12429 19775 12463 19809
rect 12521 19775 12555 19809
rect 12613 19775 12647 19809
rect 12705 19775 12739 19809
rect 12797 19775 12831 19809
rect 12889 19775 12923 19809
rect 12981 19775 13015 19809
rect 13073 19775 13107 19809
rect 13165 19775 13199 19809
rect 13257 19775 13291 19809
rect 13349 19775 13383 19809
rect 13441 19775 13475 19809
rect 13533 19775 13567 19809
rect 13625 19775 13659 19809
rect 13717 19775 13751 19809
rect 13809 19775 13843 19809
rect 13901 19775 13935 19809
rect 13993 19775 14027 19809
rect 14085 19775 14119 19809
rect 14177 19775 14211 19809
rect 14269 19775 14303 19809
rect 14361 19775 14395 19809
rect 14453 19775 14487 19809
rect 14545 19775 14579 19809
rect 14637 19775 14671 19809
rect 14729 19775 14763 19809
rect 14821 19775 14855 19809
rect 14913 19775 14947 19809
rect 15005 19775 15039 19809
rect 15097 19775 15131 19809
rect 15189 19775 15223 19809
rect 15281 19775 15315 19809
rect 15373 19775 15407 19809
rect 15465 19775 15499 19809
rect 15557 19775 15591 19809
rect 15649 19775 15683 19809
rect 15741 19775 15775 19809
rect 15833 19775 15867 19809
rect 15925 19775 15959 19809
rect 16017 19775 16051 19809
rect 16109 19775 16143 19809
rect 16201 19775 16235 19809
rect 16293 19775 16327 19809
rect 16385 19775 16419 19809
rect 16477 19775 16511 19809
rect 16569 19775 16603 19809
rect 16661 19775 16695 19809
rect 16753 19775 16787 19809
rect 16845 19775 16879 19809
rect 16937 19775 16971 19809
rect 17029 19775 17063 19809
rect 17121 19775 17155 19809
rect 17213 19775 17247 19809
rect 17305 19775 17339 19809
rect 17397 19775 17431 19809
rect 17489 19775 17523 19809
rect 17581 19775 17615 19809
rect 17673 19775 17707 19809
rect 17765 19775 17799 19809
rect 17857 19775 17891 19809
rect 17949 19775 17983 19809
rect 18041 19775 18075 19809
rect 18133 19775 18167 19809
rect 18225 19775 18259 19809
rect 18317 19775 18351 19809
rect 18409 19775 18443 19809
rect 18501 19775 18535 19809
rect 18593 19775 18627 19809
rect 18685 19775 18719 19809
rect 18777 19775 18811 19809
rect 18869 19775 18903 19809
rect 18961 19775 18995 19809
rect 19053 19775 19087 19809
rect 19145 19775 19179 19809
rect 19237 19775 19271 19809
rect 19329 19775 19363 19809
rect 19421 19775 19455 19809
rect 19513 19775 19547 19809
rect 19605 19775 19639 19809
rect 19697 19775 19731 19809
rect 19789 19775 19823 19809
rect 19881 19775 19915 19809
rect 19973 19775 20007 19809
rect 20065 19775 20099 19809
rect 20157 19775 20191 19809
rect 4977 19231 5011 19265
rect 5069 19231 5103 19265
rect 5161 19231 5195 19265
rect 5253 19231 5287 19265
rect 5345 19231 5379 19265
rect 5437 19231 5471 19265
rect 5529 19231 5563 19265
rect 5621 19231 5655 19265
rect 5713 19231 5747 19265
rect 5805 19231 5839 19265
rect 5897 19231 5931 19265
rect 5989 19231 6023 19265
rect 6081 19231 6115 19265
rect 6173 19231 6207 19265
rect 6265 19231 6299 19265
rect 6357 19231 6391 19265
rect 6449 19231 6483 19265
rect 6541 19231 6575 19265
rect 6633 19231 6667 19265
rect 6725 19231 6759 19265
rect 6817 19231 6851 19265
rect 6909 19231 6943 19265
rect 7001 19231 7035 19265
rect 7093 19231 7127 19265
rect 7185 19231 7219 19265
rect 7277 19231 7311 19265
rect 7369 19231 7403 19265
rect 7461 19231 7495 19265
rect 7553 19231 7587 19265
rect 7645 19231 7679 19265
rect 7737 19231 7771 19265
rect 7829 19231 7863 19265
rect 7921 19231 7955 19265
rect 8013 19231 8047 19265
rect 8105 19231 8139 19265
rect 8197 19231 8231 19265
rect 8289 19231 8323 19265
rect 8381 19231 8415 19265
rect 8473 19231 8507 19265
rect 8565 19231 8599 19265
rect 8657 19231 8691 19265
rect 8749 19231 8783 19265
rect 8841 19231 8875 19265
rect 8933 19231 8967 19265
rect 9025 19231 9059 19265
rect 9117 19231 9151 19265
rect 9209 19231 9243 19265
rect 9301 19231 9335 19265
rect 9393 19231 9427 19265
rect 9485 19231 9519 19265
rect 9577 19231 9611 19265
rect 9669 19231 9703 19265
rect 9761 19231 9795 19265
rect 9853 19231 9887 19265
rect 9945 19231 9979 19265
rect 10037 19231 10071 19265
rect 10129 19231 10163 19265
rect 10221 19231 10255 19265
rect 10313 19231 10347 19265
rect 10405 19231 10439 19265
rect 10497 19231 10531 19265
rect 10589 19231 10623 19265
rect 10681 19231 10715 19265
rect 10773 19231 10807 19265
rect 10865 19231 10899 19265
rect 10957 19231 10991 19265
rect 11049 19231 11083 19265
rect 11141 19231 11175 19265
rect 11233 19231 11267 19265
rect 11325 19231 11359 19265
rect 11417 19231 11451 19265
rect 11509 19231 11543 19265
rect 11601 19231 11635 19265
rect 11693 19231 11727 19265
rect 11785 19231 11819 19265
rect 11877 19231 11911 19265
rect 11969 19231 12003 19265
rect 12061 19231 12095 19265
rect 12153 19231 12187 19265
rect 12245 19231 12279 19265
rect 12337 19231 12371 19265
rect 12429 19231 12463 19265
rect 12521 19231 12555 19265
rect 12613 19231 12647 19265
rect 12705 19231 12739 19265
rect 12797 19231 12831 19265
rect 12889 19231 12923 19265
rect 12981 19231 13015 19265
rect 13073 19231 13107 19265
rect 13165 19231 13199 19265
rect 13257 19231 13291 19265
rect 13349 19231 13383 19265
rect 13441 19231 13475 19265
rect 13533 19231 13567 19265
rect 13625 19231 13659 19265
rect 13717 19231 13751 19265
rect 13809 19231 13843 19265
rect 13901 19231 13935 19265
rect 13993 19231 14027 19265
rect 14085 19231 14119 19265
rect 14177 19231 14211 19265
rect 14269 19231 14303 19265
rect 14361 19231 14395 19265
rect 14453 19231 14487 19265
rect 14545 19231 14579 19265
rect 14637 19231 14671 19265
rect 14729 19231 14763 19265
rect 14821 19231 14855 19265
rect 14913 19231 14947 19265
rect 15005 19231 15039 19265
rect 15097 19231 15131 19265
rect 15189 19231 15223 19265
rect 15281 19231 15315 19265
rect 15373 19231 15407 19265
rect 15465 19231 15499 19265
rect 15557 19231 15591 19265
rect 15649 19231 15683 19265
rect 15741 19231 15775 19265
rect 15833 19231 15867 19265
rect 15925 19231 15959 19265
rect 16017 19231 16051 19265
rect 16109 19231 16143 19265
rect 16201 19231 16235 19265
rect 16293 19231 16327 19265
rect 16385 19231 16419 19265
rect 16477 19231 16511 19265
rect 16569 19231 16603 19265
rect 16661 19231 16695 19265
rect 16753 19231 16787 19265
rect 16845 19231 16879 19265
rect 16937 19231 16971 19265
rect 17029 19231 17063 19265
rect 17121 19231 17155 19265
rect 17213 19231 17247 19265
rect 17305 19231 17339 19265
rect 17397 19231 17431 19265
rect 17489 19231 17523 19265
rect 17581 19231 17615 19265
rect 17673 19231 17707 19265
rect 17765 19231 17799 19265
rect 17857 19231 17891 19265
rect 17949 19231 17983 19265
rect 18041 19231 18075 19265
rect 18133 19231 18167 19265
rect 18225 19231 18259 19265
rect 18317 19231 18351 19265
rect 18409 19231 18443 19265
rect 18501 19231 18535 19265
rect 18593 19231 18627 19265
rect 18685 19231 18719 19265
rect 18777 19231 18811 19265
rect 18869 19231 18903 19265
rect 18961 19231 18995 19265
rect 19053 19231 19087 19265
rect 19145 19231 19179 19265
rect 19237 19231 19271 19265
rect 19329 19231 19363 19265
rect 19421 19231 19455 19265
rect 19513 19231 19547 19265
rect 19605 19231 19639 19265
rect 19697 19231 19731 19265
rect 19789 19231 19823 19265
rect 19881 19231 19915 19265
rect 19973 19231 20007 19265
rect 20065 19231 20099 19265
rect 20157 19231 20191 19265
rect 4977 18687 5011 18721
rect 5069 18687 5103 18721
rect 5161 18687 5195 18721
rect 5253 18687 5287 18721
rect 5345 18687 5379 18721
rect 5437 18687 5471 18721
rect 5529 18687 5563 18721
rect 5621 18687 5655 18721
rect 5713 18687 5747 18721
rect 5805 18687 5839 18721
rect 5897 18687 5931 18721
rect 5989 18687 6023 18721
rect 6081 18687 6115 18721
rect 6173 18687 6207 18721
rect 6265 18687 6299 18721
rect 6357 18687 6391 18721
rect 6449 18687 6483 18721
rect 6541 18687 6575 18721
rect 6633 18687 6667 18721
rect 6725 18687 6759 18721
rect 6817 18687 6851 18721
rect 6909 18687 6943 18721
rect 7001 18687 7035 18721
rect 7093 18687 7127 18721
rect 7185 18687 7219 18721
rect 7277 18687 7311 18721
rect 7369 18687 7403 18721
rect 7461 18687 7495 18721
rect 7553 18687 7587 18721
rect 7645 18687 7679 18721
rect 7737 18687 7771 18721
rect 7829 18687 7863 18721
rect 7921 18687 7955 18721
rect 8013 18687 8047 18721
rect 8105 18687 8139 18721
rect 8197 18687 8231 18721
rect 8289 18687 8323 18721
rect 8381 18687 8415 18721
rect 8473 18687 8507 18721
rect 8565 18687 8599 18721
rect 8657 18687 8691 18721
rect 8749 18687 8783 18721
rect 8841 18687 8875 18721
rect 8933 18687 8967 18721
rect 9025 18687 9059 18721
rect 9117 18687 9151 18721
rect 9209 18687 9243 18721
rect 9301 18687 9335 18721
rect 9393 18687 9427 18721
rect 9485 18687 9519 18721
rect 9577 18687 9611 18721
rect 9669 18687 9703 18721
rect 9761 18687 9795 18721
rect 9853 18687 9887 18721
rect 9945 18687 9979 18721
rect 10037 18687 10071 18721
rect 10129 18687 10163 18721
rect 10221 18687 10255 18721
rect 10313 18687 10347 18721
rect 10405 18687 10439 18721
rect 10497 18687 10531 18721
rect 10589 18687 10623 18721
rect 10681 18687 10715 18721
rect 10773 18687 10807 18721
rect 10865 18687 10899 18721
rect 10957 18687 10991 18721
rect 11049 18687 11083 18721
rect 11141 18687 11175 18721
rect 11233 18687 11267 18721
rect 11325 18687 11359 18721
rect 11417 18687 11451 18721
rect 11509 18687 11543 18721
rect 11601 18687 11635 18721
rect 11693 18687 11727 18721
rect 11785 18687 11819 18721
rect 11877 18687 11911 18721
rect 11969 18687 12003 18721
rect 12061 18687 12095 18721
rect 12153 18687 12187 18721
rect 12245 18687 12279 18721
rect 12337 18687 12371 18721
rect 12429 18687 12463 18721
rect 12521 18687 12555 18721
rect 12613 18687 12647 18721
rect 12705 18687 12739 18721
rect 12797 18687 12831 18721
rect 12889 18687 12923 18721
rect 12981 18687 13015 18721
rect 13073 18687 13107 18721
rect 13165 18687 13199 18721
rect 13257 18687 13291 18721
rect 13349 18687 13383 18721
rect 13441 18687 13475 18721
rect 13533 18687 13567 18721
rect 13625 18687 13659 18721
rect 13717 18687 13751 18721
rect 13809 18687 13843 18721
rect 13901 18687 13935 18721
rect 13993 18687 14027 18721
rect 14085 18687 14119 18721
rect 14177 18687 14211 18721
rect 14269 18687 14303 18721
rect 14361 18687 14395 18721
rect 14453 18687 14487 18721
rect 14545 18687 14579 18721
rect 14637 18687 14671 18721
rect 14729 18687 14763 18721
rect 14821 18687 14855 18721
rect 14913 18687 14947 18721
rect 15005 18687 15039 18721
rect 15097 18687 15131 18721
rect 15189 18687 15223 18721
rect 15281 18687 15315 18721
rect 15373 18687 15407 18721
rect 15465 18687 15499 18721
rect 15557 18687 15591 18721
rect 15649 18687 15683 18721
rect 15741 18687 15775 18721
rect 15833 18687 15867 18721
rect 15925 18687 15959 18721
rect 16017 18687 16051 18721
rect 16109 18687 16143 18721
rect 16201 18687 16235 18721
rect 16293 18687 16327 18721
rect 16385 18687 16419 18721
rect 16477 18687 16511 18721
rect 16569 18687 16603 18721
rect 16661 18687 16695 18721
rect 16753 18687 16787 18721
rect 16845 18687 16879 18721
rect 16937 18687 16971 18721
rect 17029 18687 17063 18721
rect 17121 18687 17155 18721
rect 17213 18687 17247 18721
rect 17305 18687 17339 18721
rect 17397 18687 17431 18721
rect 17489 18687 17523 18721
rect 17581 18687 17615 18721
rect 17673 18687 17707 18721
rect 17765 18687 17799 18721
rect 17857 18687 17891 18721
rect 17949 18687 17983 18721
rect 18041 18687 18075 18721
rect 18133 18687 18167 18721
rect 18225 18687 18259 18721
rect 18317 18687 18351 18721
rect 18409 18687 18443 18721
rect 18501 18687 18535 18721
rect 18593 18687 18627 18721
rect 18685 18687 18719 18721
rect 18777 18687 18811 18721
rect 18869 18687 18903 18721
rect 18961 18687 18995 18721
rect 19053 18687 19087 18721
rect 19145 18687 19179 18721
rect 19237 18687 19271 18721
rect 19329 18687 19363 18721
rect 19421 18687 19455 18721
rect 19513 18687 19547 18721
rect 19605 18687 19639 18721
rect 19697 18687 19731 18721
rect 19789 18687 19823 18721
rect 19881 18687 19915 18721
rect 19973 18687 20007 18721
rect 20065 18687 20099 18721
rect 20157 18687 20191 18721
rect 4977 18143 5011 18177
rect 5069 18143 5103 18177
rect 5161 18143 5195 18177
rect 5253 18143 5287 18177
rect 5345 18143 5379 18177
rect 5437 18143 5471 18177
rect 5529 18143 5563 18177
rect 5621 18143 5655 18177
rect 5713 18143 5747 18177
rect 5805 18143 5839 18177
rect 5897 18143 5931 18177
rect 5989 18143 6023 18177
rect 6081 18143 6115 18177
rect 6173 18143 6207 18177
rect 6265 18143 6299 18177
rect 6357 18143 6391 18177
rect 6449 18143 6483 18177
rect 6541 18143 6575 18177
rect 6633 18143 6667 18177
rect 6725 18143 6759 18177
rect 6817 18143 6851 18177
rect 6909 18143 6943 18177
rect 7001 18143 7035 18177
rect 7093 18143 7127 18177
rect 7185 18143 7219 18177
rect 7277 18143 7311 18177
rect 7369 18143 7403 18177
rect 7461 18143 7495 18177
rect 7553 18143 7587 18177
rect 7645 18143 7679 18177
rect 7737 18143 7771 18177
rect 7829 18143 7863 18177
rect 7921 18143 7955 18177
rect 8013 18143 8047 18177
rect 8105 18143 8139 18177
rect 8197 18143 8231 18177
rect 8289 18143 8323 18177
rect 8381 18143 8415 18177
rect 8473 18143 8507 18177
rect 8565 18143 8599 18177
rect 8657 18143 8691 18177
rect 8749 18143 8783 18177
rect 8841 18143 8875 18177
rect 8933 18143 8967 18177
rect 9025 18143 9059 18177
rect 9117 18143 9151 18177
rect 9209 18143 9243 18177
rect 9301 18143 9335 18177
rect 9393 18143 9427 18177
rect 9485 18143 9519 18177
rect 9577 18143 9611 18177
rect 9669 18143 9703 18177
rect 9761 18143 9795 18177
rect 9853 18143 9887 18177
rect 9945 18143 9979 18177
rect 10037 18143 10071 18177
rect 10129 18143 10163 18177
rect 10221 18143 10255 18177
rect 10313 18143 10347 18177
rect 10405 18143 10439 18177
rect 10497 18143 10531 18177
rect 10589 18143 10623 18177
rect 10681 18143 10715 18177
rect 10773 18143 10807 18177
rect 10865 18143 10899 18177
rect 10957 18143 10991 18177
rect 11049 18143 11083 18177
rect 11141 18143 11175 18177
rect 11233 18143 11267 18177
rect 11325 18143 11359 18177
rect 11417 18143 11451 18177
rect 11509 18143 11543 18177
rect 11601 18143 11635 18177
rect 11693 18143 11727 18177
rect 11785 18143 11819 18177
rect 11877 18143 11911 18177
rect 11969 18143 12003 18177
rect 12061 18143 12095 18177
rect 12153 18143 12187 18177
rect 12245 18143 12279 18177
rect 12337 18143 12371 18177
rect 12429 18143 12463 18177
rect 12521 18143 12555 18177
rect 12613 18143 12647 18177
rect 12705 18143 12739 18177
rect 12797 18143 12831 18177
rect 12889 18143 12923 18177
rect 12981 18143 13015 18177
rect 13073 18143 13107 18177
rect 13165 18143 13199 18177
rect 13257 18143 13291 18177
rect 13349 18143 13383 18177
rect 13441 18143 13475 18177
rect 13533 18143 13567 18177
rect 13625 18143 13659 18177
rect 13717 18143 13751 18177
rect 13809 18143 13843 18177
rect 13901 18143 13935 18177
rect 13993 18143 14027 18177
rect 14085 18143 14119 18177
rect 14177 18143 14211 18177
rect 14269 18143 14303 18177
rect 14361 18143 14395 18177
rect 14453 18143 14487 18177
rect 14545 18143 14579 18177
rect 14637 18143 14671 18177
rect 14729 18143 14763 18177
rect 14821 18143 14855 18177
rect 14913 18143 14947 18177
rect 15005 18143 15039 18177
rect 15097 18143 15131 18177
rect 15189 18143 15223 18177
rect 15281 18143 15315 18177
rect 15373 18143 15407 18177
rect 15465 18143 15499 18177
rect 15557 18143 15591 18177
rect 15649 18143 15683 18177
rect 15741 18143 15775 18177
rect 15833 18143 15867 18177
rect 15925 18143 15959 18177
rect 16017 18143 16051 18177
rect 16109 18143 16143 18177
rect 16201 18143 16235 18177
rect 16293 18143 16327 18177
rect 16385 18143 16419 18177
rect 16477 18143 16511 18177
rect 16569 18143 16603 18177
rect 16661 18143 16695 18177
rect 16753 18143 16787 18177
rect 16845 18143 16879 18177
rect 16937 18143 16971 18177
rect 17029 18143 17063 18177
rect 17121 18143 17155 18177
rect 17213 18143 17247 18177
rect 17305 18143 17339 18177
rect 17397 18143 17431 18177
rect 17489 18143 17523 18177
rect 17581 18143 17615 18177
rect 17673 18143 17707 18177
rect 17765 18143 17799 18177
rect 17857 18143 17891 18177
rect 17949 18143 17983 18177
rect 18041 18143 18075 18177
rect 18133 18143 18167 18177
rect 18225 18143 18259 18177
rect 18317 18143 18351 18177
rect 18409 18143 18443 18177
rect 18501 18143 18535 18177
rect 18593 18143 18627 18177
rect 18685 18143 18719 18177
rect 18777 18143 18811 18177
rect 18869 18143 18903 18177
rect 18961 18143 18995 18177
rect 19053 18143 19087 18177
rect 19145 18143 19179 18177
rect 19237 18143 19271 18177
rect 19329 18143 19363 18177
rect 19421 18143 19455 18177
rect 19513 18143 19547 18177
rect 19605 18143 19639 18177
rect 19697 18143 19731 18177
rect 19789 18143 19823 18177
rect 19881 18143 19915 18177
rect 19973 18143 20007 18177
rect 20065 18143 20099 18177
rect 20157 18143 20191 18177
rect 4977 17599 5011 17633
rect 5069 17599 5103 17633
rect 5161 17599 5195 17633
rect 5253 17599 5287 17633
rect 5345 17599 5379 17633
rect 5437 17599 5471 17633
rect 5529 17599 5563 17633
rect 5621 17599 5655 17633
rect 5713 17599 5747 17633
rect 5805 17599 5839 17633
rect 5897 17599 5931 17633
rect 5989 17599 6023 17633
rect 6081 17599 6115 17633
rect 6173 17599 6207 17633
rect 6265 17599 6299 17633
rect 6357 17599 6391 17633
rect 6449 17599 6483 17633
rect 6541 17599 6575 17633
rect 6633 17599 6667 17633
rect 6725 17599 6759 17633
rect 6817 17599 6851 17633
rect 6909 17599 6943 17633
rect 7001 17599 7035 17633
rect 7093 17599 7127 17633
rect 7185 17599 7219 17633
rect 7277 17599 7311 17633
rect 7369 17599 7403 17633
rect 7461 17599 7495 17633
rect 7553 17599 7587 17633
rect 7645 17599 7679 17633
rect 7737 17599 7771 17633
rect 7829 17599 7863 17633
rect 7921 17599 7955 17633
rect 8013 17599 8047 17633
rect 8105 17599 8139 17633
rect 8197 17599 8231 17633
rect 8289 17599 8323 17633
rect 8381 17599 8415 17633
rect 8473 17599 8507 17633
rect 8565 17599 8599 17633
rect 8657 17599 8691 17633
rect 8749 17599 8783 17633
rect 8841 17599 8875 17633
rect 8933 17599 8967 17633
rect 9025 17599 9059 17633
rect 9117 17599 9151 17633
rect 9209 17599 9243 17633
rect 9301 17599 9335 17633
rect 9393 17599 9427 17633
rect 9485 17599 9519 17633
rect 9577 17599 9611 17633
rect 9669 17599 9703 17633
rect 9761 17599 9795 17633
rect 9853 17599 9887 17633
rect 9945 17599 9979 17633
rect 10037 17599 10071 17633
rect 10129 17599 10163 17633
rect 10221 17599 10255 17633
rect 10313 17599 10347 17633
rect 10405 17599 10439 17633
rect 10497 17599 10531 17633
rect 10589 17599 10623 17633
rect 10681 17599 10715 17633
rect 10773 17599 10807 17633
rect 10865 17599 10899 17633
rect 10957 17599 10991 17633
rect 11049 17599 11083 17633
rect 11141 17599 11175 17633
rect 11233 17599 11267 17633
rect 11325 17599 11359 17633
rect 11417 17599 11451 17633
rect 11509 17599 11543 17633
rect 11601 17599 11635 17633
rect 11693 17599 11727 17633
rect 11785 17599 11819 17633
rect 11877 17599 11911 17633
rect 11969 17599 12003 17633
rect 12061 17599 12095 17633
rect 12153 17599 12187 17633
rect 12245 17599 12279 17633
rect 12337 17599 12371 17633
rect 12429 17599 12463 17633
rect 12521 17599 12555 17633
rect 12613 17599 12647 17633
rect 12705 17599 12739 17633
rect 12797 17599 12831 17633
rect 12889 17599 12923 17633
rect 12981 17599 13015 17633
rect 13073 17599 13107 17633
rect 13165 17599 13199 17633
rect 13257 17599 13291 17633
rect 13349 17599 13383 17633
rect 13441 17599 13475 17633
rect 13533 17599 13567 17633
rect 13625 17599 13659 17633
rect 13717 17599 13751 17633
rect 13809 17599 13843 17633
rect 13901 17599 13935 17633
rect 13993 17599 14027 17633
rect 14085 17599 14119 17633
rect 14177 17599 14211 17633
rect 14269 17599 14303 17633
rect 14361 17599 14395 17633
rect 14453 17599 14487 17633
rect 14545 17599 14579 17633
rect 14637 17599 14671 17633
rect 14729 17599 14763 17633
rect 14821 17599 14855 17633
rect 14913 17599 14947 17633
rect 15005 17599 15039 17633
rect 15097 17599 15131 17633
rect 15189 17599 15223 17633
rect 15281 17599 15315 17633
rect 15373 17599 15407 17633
rect 15465 17599 15499 17633
rect 15557 17599 15591 17633
rect 15649 17599 15683 17633
rect 15741 17599 15775 17633
rect 15833 17599 15867 17633
rect 15925 17599 15959 17633
rect 16017 17599 16051 17633
rect 16109 17599 16143 17633
rect 16201 17599 16235 17633
rect 16293 17599 16327 17633
rect 16385 17599 16419 17633
rect 16477 17599 16511 17633
rect 16569 17599 16603 17633
rect 16661 17599 16695 17633
rect 16753 17599 16787 17633
rect 16845 17599 16879 17633
rect 16937 17599 16971 17633
rect 17029 17599 17063 17633
rect 17121 17599 17155 17633
rect 17213 17599 17247 17633
rect 17305 17599 17339 17633
rect 17397 17599 17431 17633
rect 17489 17599 17523 17633
rect 17581 17599 17615 17633
rect 17673 17599 17707 17633
rect 17765 17599 17799 17633
rect 17857 17599 17891 17633
rect 17949 17599 17983 17633
rect 18041 17599 18075 17633
rect 18133 17599 18167 17633
rect 18225 17599 18259 17633
rect 18317 17599 18351 17633
rect 18409 17599 18443 17633
rect 18501 17599 18535 17633
rect 18593 17599 18627 17633
rect 18685 17599 18719 17633
rect 18777 17599 18811 17633
rect 18869 17599 18903 17633
rect 18961 17599 18995 17633
rect 19053 17599 19087 17633
rect 19145 17599 19179 17633
rect 19237 17599 19271 17633
rect 19329 17599 19363 17633
rect 19421 17599 19455 17633
rect 19513 17599 19547 17633
rect 19605 17599 19639 17633
rect 19697 17599 19731 17633
rect 19789 17599 19823 17633
rect 19881 17599 19915 17633
rect 19973 17599 20007 17633
rect 20065 17599 20099 17633
rect 20157 17599 20191 17633
rect 4977 17055 5011 17089
rect 5069 17055 5103 17089
rect 5161 17055 5195 17089
rect 5253 17055 5287 17089
rect 5345 17055 5379 17089
rect 5437 17055 5471 17089
rect 5529 17055 5563 17089
rect 5621 17055 5655 17089
rect 5713 17055 5747 17089
rect 5805 17055 5839 17089
rect 5897 17055 5931 17089
rect 5989 17055 6023 17089
rect 6081 17055 6115 17089
rect 6173 17055 6207 17089
rect 6265 17055 6299 17089
rect 6357 17055 6391 17089
rect 6449 17055 6483 17089
rect 6541 17055 6575 17089
rect 6633 17055 6667 17089
rect 6725 17055 6759 17089
rect 6817 17055 6851 17089
rect 6909 17055 6943 17089
rect 7001 17055 7035 17089
rect 7093 17055 7127 17089
rect 7185 17055 7219 17089
rect 7277 17055 7311 17089
rect 7369 17055 7403 17089
rect 7461 17055 7495 17089
rect 7553 17055 7587 17089
rect 7645 17055 7679 17089
rect 7737 17055 7771 17089
rect 7829 17055 7863 17089
rect 7921 17055 7955 17089
rect 8013 17055 8047 17089
rect 8105 17055 8139 17089
rect 8197 17055 8231 17089
rect 8289 17055 8323 17089
rect 8381 17055 8415 17089
rect 8473 17055 8507 17089
rect 8565 17055 8599 17089
rect 8657 17055 8691 17089
rect 8749 17055 8783 17089
rect 8841 17055 8875 17089
rect 8933 17055 8967 17089
rect 9025 17055 9059 17089
rect 9117 17055 9151 17089
rect 9209 17055 9243 17089
rect 9301 17055 9335 17089
rect 9393 17055 9427 17089
rect 9485 17055 9519 17089
rect 9577 17055 9611 17089
rect 9669 17055 9703 17089
rect 9761 17055 9795 17089
rect 9853 17055 9887 17089
rect 9945 17055 9979 17089
rect 10037 17055 10071 17089
rect 10129 17055 10163 17089
rect 10221 17055 10255 17089
rect 10313 17055 10347 17089
rect 10405 17055 10439 17089
rect 10497 17055 10531 17089
rect 10589 17055 10623 17089
rect 10681 17055 10715 17089
rect 10773 17055 10807 17089
rect 10865 17055 10899 17089
rect 10957 17055 10991 17089
rect 11049 17055 11083 17089
rect 11141 17055 11175 17089
rect 11233 17055 11267 17089
rect 11325 17055 11359 17089
rect 11417 17055 11451 17089
rect 11509 17055 11543 17089
rect 11601 17055 11635 17089
rect 11693 17055 11727 17089
rect 11785 17055 11819 17089
rect 11877 17055 11911 17089
rect 11969 17055 12003 17089
rect 12061 17055 12095 17089
rect 12153 17055 12187 17089
rect 12245 17055 12279 17089
rect 12337 17055 12371 17089
rect 12429 17055 12463 17089
rect 12521 17055 12555 17089
rect 12613 17055 12647 17089
rect 12705 17055 12739 17089
rect 12797 17055 12831 17089
rect 12889 17055 12923 17089
rect 12981 17055 13015 17089
rect 13073 17055 13107 17089
rect 13165 17055 13199 17089
rect 13257 17055 13291 17089
rect 13349 17055 13383 17089
rect 13441 17055 13475 17089
rect 13533 17055 13567 17089
rect 13625 17055 13659 17089
rect 13717 17055 13751 17089
rect 13809 17055 13843 17089
rect 13901 17055 13935 17089
rect 13993 17055 14027 17089
rect 14085 17055 14119 17089
rect 14177 17055 14211 17089
rect 14269 17055 14303 17089
rect 14361 17055 14395 17089
rect 14453 17055 14487 17089
rect 14545 17055 14579 17089
rect 14637 17055 14671 17089
rect 14729 17055 14763 17089
rect 14821 17055 14855 17089
rect 14913 17055 14947 17089
rect 15005 17055 15039 17089
rect 15097 17055 15131 17089
rect 15189 17055 15223 17089
rect 15281 17055 15315 17089
rect 15373 17055 15407 17089
rect 15465 17055 15499 17089
rect 15557 17055 15591 17089
rect 15649 17055 15683 17089
rect 15741 17055 15775 17089
rect 15833 17055 15867 17089
rect 15925 17055 15959 17089
rect 16017 17055 16051 17089
rect 16109 17055 16143 17089
rect 16201 17055 16235 17089
rect 16293 17055 16327 17089
rect 16385 17055 16419 17089
rect 16477 17055 16511 17089
rect 16569 17055 16603 17089
rect 16661 17055 16695 17089
rect 16753 17055 16787 17089
rect 16845 17055 16879 17089
rect 16937 17055 16971 17089
rect 17029 17055 17063 17089
rect 17121 17055 17155 17089
rect 17213 17055 17247 17089
rect 17305 17055 17339 17089
rect 17397 17055 17431 17089
rect 17489 17055 17523 17089
rect 17581 17055 17615 17089
rect 17673 17055 17707 17089
rect 17765 17055 17799 17089
rect 17857 17055 17891 17089
rect 17949 17055 17983 17089
rect 18041 17055 18075 17089
rect 18133 17055 18167 17089
rect 18225 17055 18259 17089
rect 18317 17055 18351 17089
rect 18409 17055 18443 17089
rect 18501 17055 18535 17089
rect 18593 17055 18627 17089
rect 18685 17055 18719 17089
rect 18777 17055 18811 17089
rect 18869 17055 18903 17089
rect 18961 17055 18995 17089
rect 19053 17055 19087 17089
rect 19145 17055 19179 17089
rect 19237 17055 19271 17089
rect 19329 17055 19363 17089
rect 19421 17055 19455 17089
rect 19513 17055 19547 17089
rect 19605 17055 19639 17089
rect 19697 17055 19731 17089
rect 19789 17055 19823 17089
rect 19881 17055 19915 17089
rect 19973 17055 20007 17089
rect 20065 17055 20099 17089
rect 20157 17055 20191 17089
rect 4977 16511 5011 16545
rect 5069 16511 5103 16545
rect 5161 16511 5195 16545
rect 5253 16511 5287 16545
rect 5345 16511 5379 16545
rect 5437 16511 5471 16545
rect 5529 16511 5563 16545
rect 5621 16511 5655 16545
rect 5713 16511 5747 16545
rect 5805 16511 5839 16545
rect 5897 16511 5931 16545
rect 5989 16511 6023 16545
rect 6081 16511 6115 16545
rect 6173 16511 6207 16545
rect 6265 16511 6299 16545
rect 6357 16511 6391 16545
rect 6449 16511 6483 16545
rect 6541 16511 6575 16545
rect 6633 16511 6667 16545
rect 6725 16511 6759 16545
rect 6817 16511 6851 16545
rect 6909 16511 6943 16545
rect 7001 16511 7035 16545
rect 7093 16511 7127 16545
rect 7185 16511 7219 16545
rect 7277 16511 7311 16545
rect 7369 16511 7403 16545
rect 7461 16511 7495 16545
rect 7553 16511 7587 16545
rect 7645 16511 7679 16545
rect 7737 16511 7771 16545
rect 7829 16511 7863 16545
rect 7921 16511 7955 16545
rect 8013 16511 8047 16545
rect 8105 16511 8139 16545
rect 8197 16511 8231 16545
rect 8289 16511 8323 16545
rect 8381 16511 8415 16545
rect 8473 16511 8507 16545
rect 8565 16511 8599 16545
rect 8657 16511 8691 16545
rect 8749 16511 8783 16545
rect 8841 16511 8875 16545
rect 8933 16511 8967 16545
rect 9025 16511 9059 16545
rect 9117 16511 9151 16545
rect 9209 16511 9243 16545
rect 9301 16511 9335 16545
rect 9393 16511 9427 16545
rect 9485 16511 9519 16545
rect 9577 16511 9611 16545
rect 9669 16511 9703 16545
rect 9761 16511 9795 16545
rect 9853 16511 9887 16545
rect 9945 16511 9979 16545
rect 10037 16511 10071 16545
rect 10129 16511 10163 16545
rect 10221 16511 10255 16545
rect 10313 16511 10347 16545
rect 10405 16511 10439 16545
rect 10497 16511 10531 16545
rect 10589 16511 10623 16545
rect 10681 16511 10715 16545
rect 10773 16511 10807 16545
rect 10865 16511 10899 16545
rect 10957 16511 10991 16545
rect 11049 16511 11083 16545
rect 11141 16511 11175 16545
rect 11233 16511 11267 16545
rect 11325 16511 11359 16545
rect 11417 16511 11451 16545
rect 11509 16511 11543 16545
rect 11601 16511 11635 16545
rect 11693 16511 11727 16545
rect 11785 16511 11819 16545
rect 11877 16511 11911 16545
rect 11969 16511 12003 16545
rect 12061 16511 12095 16545
rect 12153 16511 12187 16545
rect 12245 16511 12279 16545
rect 12337 16511 12371 16545
rect 12429 16511 12463 16545
rect 12521 16511 12555 16545
rect 12613 16511 12647 16545
rect 12705 16511 12739 16545
rect 12797 16511 12831 16545
rect 12889 16511 12923 16545
rect 12981 16511 13015 16545
rect 13073 16511 13107 16545
rect 13165 16511 13199 16545
rect 13257 16511 13291 16545
rect 13349 16511 13383 16545
rect 13441 16511 13475 16545
rect 13533 16511 13567 16545
rect 13625 16511 13659 16545
rect 13717 16511 13751 16545
rect 13809 16511 13843 16545
rect 13901 16511 13935 16545
rect 13993 16511 14027 16545
rect 14085 16511 14119 16545
rect 14177 16511 14211 16545
rect 14269 16511 14303 16545
rect 14361 16511 14395 16545
rect 14453 16511 14487 16545
rect 14545 16511 14579 16545
rect 14637 16511 14671 16545
rect 14729 16511 14763 16545
rect 14821 16511 14855 16545
rect 14913 16511 14947 16545
rect 15005 16511 15039 16545
rect 15097 16511 15131 16545
rect 15189 16511 15223 16545
rect 15281 16511 15315 16545
rect 15373 16511 15407 16545
rect 15465 16511 15499 16545
rect 15557 16511 15591 16545
rect 15649 16511 15683 16545
rect 15741 16511 15775 16545
rect 15833 16511 15867 16545
rect 15925 16511 15959 16545
rect 16017 16511 16051 16545
rect 16109 16511 16143 16545
rect 16201 16511 16235 16545
rect 16293 16511 16327 16545
rect 16385 16511 16419 16545
rect 16477 16511 16511 16545
rect 16569 16511 16603 16545
rect 16661 16511 16695 16545
rect 16753 16511 16787 16545
rect 16845 16511 16879 16545
rect 16937 16511 16971 16545
rect 17029 16511 17063 16545
rect 17121 16511 17155 16545
rect 17213 16511 17247 16545
rect 17305 16511 17339 16545
rect 17397 16511 17431 16545
rect 17489 16511 17523 16545
rect 17581 16511 17615 16545
rect 17673 16511 17707 16545
rect 17765 16511 17799 16545
rect 17857 16511 17891 16545
rect 17949 16511 17983 16545
rect 18041 16511 18075 16545
rect 18133 16511 18167 16545
rect 18225 16511 18259 16545
rect 18317 16511 18351 16545
rect 18409 16511 18443 16545
rect 18501 16511 18535 16545
rect 18593 16511 18627 16545
rect 18685 16511 18719 16545
rect 18777 16511 18811 16545
rect 18869 16511 18903 16545
rect 18961 16511 18995 16545
rect 19053 16511 19087 16545
rect 19145 16511 19179 16545
rect 19237 16511 19271 16545
rect 19329 16511 19363 16545
rect 19421 16511 19455 16545
rect 19513 16511 19547 16545
rect 19605 16511 19639 16545
rect 19697 16511 19731 16545
rect 19789 16511 19823 16545
rect 19881 16511 19915 16545
rect 19973 16511 20007 16545
rect 20065 16511 20099 16545
rect 20157 16511 20191 16545
rect 4977 15967 5011 16001
rect 5069 15967 5103 16001
rect 5161 15967 5195 16001
rect 5253 15967 5287 16001
rect 5345 15967 5379 16001
rect 5437 15967 5471 16001
rect 5529 15967 5563 16001
rect 5621 15967 5655 16001
rect 5713 15967 5747 16001
rect 5805 15967 5839 16001
rect 5897 15967 5931 16001
rect 5989 15967 6023 16001
rect 6081 15967 6115 16001
rect 6173 15967 6207 16001
rect 6265 15967 6299 16001
rect 6357 15967 6391 16001
rect 6449 15967 6483 16001
rect 6541 15967 6575 16001
rect 6633 15967 6667 16001
rect 6725 15967 6759 16001
rect 6817 15967 6851 16001
rect 6909 15967 6943 16001
rect 7001 15967 7035 16001
rect 7093 15967 7127 16001
rect 7185 15967 7219 16001
rect 7277 15967 7311 16001
rect 7369 15967 7403 16001
rect 7461 15967 7495 16001
rect 7553 15967 7587 16001
rect 7645 15967 7679 16001
rect 7737 15967 7771 16001
rect 7829 15967 7863 16001
rect 7921 15967 7955 16001
rect 8013 15967 8047 16001
rect 8105 15967 8139 16001
rect 8197 15967 8231 16001
rect 8289 15967 8323 16001
rect 8381 15967 8415 16001
rect 8473 15967 8507 16001
rect 8565 15967 8599 16001
rect 8657 15967 8691 16001
rect 8749 15967 8783 16001
rect 8841 15967 8875 16001
rect 8933 15967 8967 16001
rect 9025 15967 9059 16001
rect 9117 15967 9151 16001
rect 9209 15967 9243 16001
rect 9301 15967 9335 16001
rect 9393 15967 9427 16001
rect 9485 15967 9519 16001
rect 9577 15967 9611 16001
rect 9669 15967 9703 16001
rect 9761 15967 9795 16001
rect 9853 15967 9887 16001
rect 9945 15967 9979 16001
rect 10037 15967 10071 16001
rect 10129 15967 10163 16001
rect 10221 15967 10255 16001
rect 10313 15967 10347 16001
rect 10405 15967 10439 16001
rect 10497 15967 10531 16001
rect 10589 15967 10623 16001
rect 10681 15967 10715 16001
rect 10773 15967 10807 16001
rect 10865 15967 10899 16001
rect 10957 15967 10991 16001
rect 11049 15967 11083 16001
rect 11141 15967 11175 16001
rect 11233 15967 11267 16001
rect 11325 15967 11359 16001
rect 11417 15967 11451 16001
rect 11509 15967 11543 16001
rect 11601 15967 11635 16001
rect 11693 15967 11727 16001
rect 11785 15967 11819 16001
rect 11877 15967 11911 16001
rect 11969 15967 12003 16001
rect 12061 15967 12095 16001
rect 12153 15967 12187 16001
rect 12245 15967 12279 16001
rect 12337 15967 12371 16001
rect 12429 15967 12463 16001
rect 12521 15967 12555 16001
rect 12613 15967 12647 16001
rect 12705 15967 12739 16001
rect 12797 15967 12831 16001
rect 12889 15967 12923 16001
rect 12981 15967 13015 16001
rect 13073 15967 13107 16001
rect 13165 15967 13199 16001
rect 13257 15967 13291 16001
rect 13349 15967 13383 16001
rect 13441 15967 13475 16001
rect 13533 15967 13567 16001
rect 13625 15967 13659 16001
rect 13717 15967 13751 16001
rect 13809 15967 13843 16001
rect 13901 15967 13935 16001
rect 13993 15967 14027 16001
rect 14085 15967 14119 16001
rect 14177 15967 14211 16001
rect 14269 15967 14303 16001
rect 14361 15967 14395 16001
rect 14453 15967 14487 16001
rect 14545 15967 14579 16001
rect 14637 15967 14671 16001
rect 14729 15967 14763 16001
rect 14821 15967 14855 16001
rect 14913 15967 14947 16001
rect 15005 15967 15039 16001
rect 15097 15967 15131 16001
rect 15189 15967 15223 16001
rect 15281 15967 15315 16001
rect 15373 15967 15407 16001
rect 15465 15967 15499 16001
rect 15557 15967 15591 16001
rect 15649 15967 15683 16001
rect 15741 15967 15775 16001
rect 15833 15967 15867 16001
rect 15925 15967 15959 16001
rect 16017 15967 16051 16001
rect 16109 15967 16143 16001
rect 16201 15967 16235 16001
rect 16293 15967 16327 16001
rect 16385 15967 16419 16001
rect 16477 15967 16511 16001
rect 16569 15967 16603 16001
rect 16661 15967 16695 16001
rect 16753 15967 16787 16001
rect 16845 15967 16879 16001
rect 16937 15967 16971 16001
rect 17029 15967 17063 16001
rect 17121 15967 17155 16001
rect 17213 15967 17247 16001
rect 17305 15967 17339 16001
rect 17397 15967 17431 16001
rect 17489 15967 17523 16001
rect 17581 15967 17615 16001
rect 17673 15967 17707 16001
rect 17765 15967 17799 16001
rect 17857 15967 17891 16001
rect 17949 15967 17983 16001
rect 18041 15967 18075 16001
rect 18133 15967 18167 16001
rect 18225 15967 18259 16001
rect 18317 15967 18351 16001
rect 18409 15967 18443 16001
rect 18501 15967 18535 16001
rect 18593 15967 18627 16001
rect 18685 15967 18719 16001
rect 18777 15967 18811 16001
rect 18869 15967 18903 16001
rect 18961 15967 18995 16001
rect 19053 15967 19087 16001
rect 19145 15967 19179 16001
rect 19237 15967 19271 16001
rect 19329 15967 19363 16001
rect 19421 15967 19455 16001
rect 19513 15967 19547 16001
rect 19605 15967 19639 16001
rect 19697 15967 19731 16001
rect 19789 15967 19823 16001
rect 19881 15967 19915 16001
rect 19973 15967 20007 16001
rect 20065 15967 20099 16001
rect 20157 15967 20191 16001
rect 4977 15423 5011 15457
rect 5069 15423 5103 15457
rect 5161 15423 5195 15457
rect 5253 15423 5287 15457
rect 5345 15423 5379 15457
rect 5437 15423 5471 15457
rect 5529 15423 5563 15457
rect 5621 15423 5655 15457
rect 5713 15423 5747 15457
rect 5805 15423 5839 15457
rect 5897 15423 5931 15457
rect 5989 15423 6023 15457
rect 6081 15423 6115 15457
rect 6173 15423 6207 15457
rect 6265 15423 6299 15457
rect 6357 15423 6391 15457
rect 6449 15423 6483 15457
rect 6541 15423 6575 15457
rect 6633 15423 6667 15457
rect 6725 15423 6759 15457
rect 6817 15423 6851 15457
rect 6909 15423 6943 15457
rect 7001 15423 7035 15457
rect 7093 15423 7127 15457
rect 7185 15423 7219 15457
rect 7277 15423 7311 15457
rect 7369 15423 7403 15457
rect 7461 15423 7495 15457
rect 7553 15423 7587 15457
rect 7645 15423 7679 15457
rect 7737 15423 7771 15457
rect 7829 15423 7863 15457
rect 7921 15423 7955 15457
rect 8013 15423 8047 15457
rect 8105 15423 8139 15457
rect 8197 15423 8231 15457
rect 8289 15423 8323 15457
rect 8381 15423 8415 15457
rect 8473 15423 8507 15457
rect 8565 15423 8599 15457
rect 8657 15423 8691 15457
rect 8749 15423 8783 15457
rect 8841 15423 8875 15457
rect 8933 15423 8967 15457
rect 9025 15423 9059 15457
rect 9117 15423 9151 15457
rect 9209 15423 9243 15457
rect 9301 15423 9335 15457
rect 9393 15423 9427 15457
rect 9485 15423 9519 15457
rect 9577 15423 9611 15457
rect 9669 15423 9703 15457
rect 9761 15423 9795 15457
rect 9853 15423 9887 15457
rect 9945 15423 9979 15457
rect 10037 15423 10071 15457
rect 10129 15423 10163 15457
rect 10221 15423 10255 15457
rect 10313 15423 10347 15457
rect 10405 15423 10439 15457
rect 10497 15423 10531 15457
rect 10589 15423 10623 15457
rect 10681 15423 10715 15457
rect 10773 15423 10807 15457
rect 10865 15423 10899 15457
rect 10957 15423 10991 15457
rect 11049 15423 11083 15457
rect 11141 15423 11175 15457
rect 11233 15423 11267 15457
rect 11325 15423 11359 15457
rect 11417 15423 11451 15457
rect 11509 15423 11543 15457
rect 11601 15423 11635 15457
rect 11693 15423 11727 15457
rect 11785 15423 11819 15457
rect 11877 15423 11911 15457
rect 11969 15423 12003 15457
rect 12061 15423 12095 15457
rect 12153 15423 12187 15457
rect 12245 15423 12279 15457
rect 12337 15423 12371 15457
rect 12429 15423 12463 15457
rect 12521 15423 12555 15457
rect 12613 15423 12647 15457
rect 12705 15423 12739 15457
rect 12797 15423 12831 15457
rect 12889 15423 12923 15457
rect 12981 15423 13015 15457
rect 13073 15423 13107 15457
rect 13165 15423 13199 15457
rect 13257 15423 13291 15457
rect 13349 15423 13383 15457
rect 13441 15423 13475 15457
rect 13533 15423 13567 15457
rect 13625 15423 13659 15457
rect 13717 15423 13751 15457
rect 13809 15423 13843 15457
rect 13901 15423 13935 15457
rect 13993 15423 14027 15457
rect 14085 15423 14119 15457
rect 14177 15423 14211 15457
rect 14269 15423 14303 15457
rect 14361 15423 14395 15457
rect 14453 15423 14487 15457
rect 14545 15423 14579 15457
rect 14637 15423 14671 15457
rect 14729 15423 14763 15457
rect 14821 15423 14855 15457
rect 14913 15423 14947 15457
rect 15005 15423 15039 15457
rect 15097 15423 15131 15457
rect 15189 15423 15223 15457
rect 15281 15423 15315 15457
rect 15373 15423 15407 15457
rect 15465 15423 15499 15457
rect 15557 15423 15591 15457
rect 15649 15423 15683 15457
rect 15741 15423 15775 15457
rect 15833 15423 15867 15457
rect 15925 15423 15959 15457
rect 16017 15423 16051 15457
rect 16109 15423 16143 15457
rect 16201 15423 16235 15457
rect 16293 15423 16327 15457
rect 16385 15423 16419 15457
rect 16477 15423 16511 15457
rect 16569 15423 16603 15457
rect 16661 15423 16695 15457
rect 16753 15423 16787 15457
rect 16845 15423 16879 15457
rect 16937 15423 16971 15457
rect 17029 15423 17063 15457
rect 17121 15423 17155 15457
rect 17213 15423 17247 15457
rect 17305 15423 17339 15457
rect 17397 15423 17431 15457
rect 17489 15423 17523 15457
rect 17581 15423 17615 15457
rect 17673 15423 17707 15457
rect 17765 15423 17799 15457
rect 17857 15423 17891 15457
rect 17949 15423 17983 15457
rect 18041 15423 18075 15457
rect 18133 15423 18167 15457
rect 18225 15423 18259 15457
rect 18317 15423 18351 15457
rect 18409 15423 18443 15457
rect 18501 15423 18535 15457
rect 18593 15423 18627 15457
rect 18685 15423 18719 15457
rect 18777 15423 18811 15457
rect 18869 15423 18903 15457
rect 18961 15423 18995 15457
rect 19053 15423 19087 15457
rect 19145 15423 19179 15457
rect 19237 15423 19271 15457
rect 19329 15423 19363 15457
rect 19421 15423 19455 15457
rect 19513 15423 19547 15457
rect 19605 15423 19639 15457
rect 19697 15423 19731 15457
rect 19789 15423 19823 15457
rect 19881 15423 19915 15457
rect 19973 15423 20007 15457
rect 20065 15423 20099 15457
rect 20157 15423 20191 15457
rect 12889 15117 12923 15151
rect 13441 14981 13450 15015
rect 13450 14981 13475 15015
rect 15373 15117 15407 15151
rect 16017 14981 16026 15015
rect 16026 14981 16051 15015
rect 4977 14879 5011 14913
rect 5069 14879 5103 14913
rect 5161 14879 5195 14913
rect 5253 14879 5287 14913
rect 5345 14879 5379 14913
rect 5437 14879 5471 14913
rect 5529 14879 5563 14913
rect 5621 14879 5655 14913
rect 5713 14879 5747 14913
rect 5805 14879 5839 14913
rect 5897 14879 5931 14913
rect 5989 14879 6023 14913
rect 6081 14879 6115 14913
rect 6173 14879 6207 14913
rect 6265 14879 6299 14913
rect 6357 14879 6391 14913
rect 6449 14879 6483 14913
rect 6541 14879 6575 14913
rect 6633 14879 6667 14913
rect 6725 14879 6759 14913
rect 6817 14879 6851 14913
rect 6909 14879 6943 14913
rect 7001 14879 7035 14913
rect 7093 14879 7127 14913
rect 7185 14879 7219 14913
rect 7277 14879 7311 14913
rect 7369 14879 7403 14913
rect 7461 14879 7495 14913
rect 7553 14879 7587 14913
rect 7645 14879 7679 14913
rect 7737 14879 7771 14913
rect 7829 14879 7863 14913
rect 7921 14879 7955 14913
rect 8013 14879 8047 14913
rect 8105 14879 8139 14913
rect 8197 14879 8231 14913
rect 8289 14879 8323 14913
rect 8381 14879 8415 14913
rect 8473 14879 8507 14913
rect 8565 14879 8599 14913
rect 8657 14879 8691 14913
rect 8749 14879 8783 14913
rect 8841 14879 8875 14913
rect 8933 14879 8967 14913
rect 9025 14879 9059 14913
rect 9117 14879 9151 14913
rect 9209 14879 9243 14913
rect 9301 14879 9335 14913
rect 9393 14879 9427 14913
rect 9485 14879 9519 14913
rect 9577 14879 9611 14913
rect 9669 14879 9703 14913
rect 9761 14879 9795 14913
rect 9853 14879 9887 14913
rect 9945 14879 9979 14913
rect 10037 14879 10071 14913
rect 10129 14879 10163 14913
rect 10221 14879 10255 14913
rect 10313 14879 10347 14913
rect 10405 14879 10439 14913
rect 10497 14879 10531 14913
rect 10589 14879 10623 14913
rect 10681 14879 10715 14913
rect 10773 14879 10807 14913
rect 10865 14879 10899 14913
rect 10957 14879 10991 14913
rect 11049 14879 11083 14913
rect 11141 14879 11175 14913
rect 11233 14879 11267 14913
rect 11325 14879 11359 14913
rect 11417 14879 11451 14913
rect 11509 14879 11543 14913
rect 11601 14879 11635 14913
rect 11693 14879 11727 14913
rect 11785 14879 11819 14913
rect 11877 14879 11911 14913
rect 11969 14879 12003 14913
rect 12061 14879 12095 14913
rect 12153 14879 12187 14913
rect 12245 14879 12279 14913
rect 12337 14879 12371 14913
rect 12429 14879 12463 14913
rect 12521 14879 12555 14913
rect 12613 14879 12647 14913
rect 12705 14879 12739 14913
rect 12797 14879 12831 14913
rect 12889 14879 12923 14913
rect 12981 14879 13015 14913
rect 13073 14879 13107 14913
rect 13165 14879 13199 14913
rect 13257 14879 13291 14913
rect 13349 14879 13383 14913
rect 13441 14879 13475 14913
rect 13533 14879 13567 14913
rect 13625 14879 13659 14913
rect 13717 14879 13751 14913
rect 13809 14879 13843 14913
rect 13901 14879 13935 14913
rect 13993 14879 14027 14913
rect 14085 14879 14119 14913
rect 14177 14879 14211 14913
rect 14269 14879 14303 14913
rect 14361 14879 14395 14913
rect 14453 14879 14487 14913
rect 14545 14879 14579 14913
rect 14637 14879 14671 14913
rect 14729 14879 14763 14913
rect 14821 14879 14855 14913
rect 14913 14879 14947 14913
rect 15005 14879 15039 14913
rect 15097 14879 15131 14913
rect 15189 14879 15223 14913
rect 15281 14879 15315 14913
rect 15373 14879 15407 14913
rect 15465 14879 15499 14913
rect 15557 14879 15591 14913
rect 15649 14879 15683 14913
rect 15741 14879 15775 14913
rect 15833 14879 15867 14913
rect 15925 14879 15959 14913
rect 16017 14879 16051 14913
rect 16109 14879 16143 14913
rect 16201 14879 16235 14913
rect 16293 14879 16327 14913
rect 16385 14879 16419 14913
rect 16477 14879 16511 14913
rect 16569 14879 16603 14913
rect 16661 14879 16695 14913
rect 16753 14879 16787 14913
rect 16845 14879 16879 14913
rect 16937 14879 16971 14913
rect 17029 14879 17063 14913
rect 17121 14879 17155 14913
rect 17213 14879 17247 14913
rect 17305 14879 17339 14913
rect 17397 14879 17431 14913
rect 17489 14879 17523 14913
rect 17581 14879 17615 14913
rect 17673 14879 17707 14913
rect 17765 14879 17799 14913
rect 17857 14879 17891 14913
rect 17949 14879 17983 14913
rect 18041 14879 18075 14913
rect 18133 14879 18167 14913
rect 18225 14879 18259 14913
rect 18317 14879 18351 14913
rect 18409 14879 18443 14913
rect 18501 14879 18535 14913
rect 18593 14879 18627 14913
rect 18685 14879 18719 14913
rect 18777 14879 18811 14913
rect 18869 14879 18903 14913
rect 18961 14879 18995 14913
rect 19053 14879 19087 14913
rect 19145 14879 19179 14913
rect 19237 14879 19271 14913
rect 19329 14879 19363 14913
rect 19421 14879 19455 14913
rect 19513 14879 19547 14913
rect 19605 14879 19639 14913
rect 19697 14879 19731 14913
rect 19789 14879 19823 14913
rect 19881 14879 19915 14913
rect 19973 14879 20007 14913
rect 20065 14879 20099 14913
rect 20157 14879 20191 14913
rect 10865 14641 10899 14675
rect 10957 14437 10991 14471
rect 11049 14573 11083 14607
rect 12889 14641 12923 14675
rect 11417 14464 11451 14471
rect 11417 14437 11445 14464
rect 11445 14437 11451 14464
rect 12981 14437 13015 14471
rect 13073 14573 13107 14607
rect 14453 14714 14481 14743
rect 14481 14714 14487 14743
rect 14453 14709 14487 14714
rect 14269 14601 14303 14607
rect 14269 14573 14277 14601
rect 14277 14573 14303 14601
rect 13441 14464 13475 14471
rect 13441 14437 13469 14464
rect 13469 14437 13475 14464
rect 15117 14717 15151 14743
rect 15117 14709 15120 14717
rect 15120 14709 15151 14717
rect 14545 14461 14551 14471
rect 14551 14461 14579 14471
rect 14901 14593 14935 14602
rect 14901 14568 14919 14593
rect 14919 14568 14935 14593
rect 14841 14505 14875 14539
rect 14545 14437 14579 14461
rect 15117 14591 15151 14607
rect 15117 14573 15125 14591
rect 15125 14573 15151 14591
rect 15741 14709 15775 14743
rect 15489 14521 15499 14539
rect 15499 14521 15523 14539
rect 15489 14505 15523 14521
rect 15561 14505 15595 14539
rect 15833 14573 15867 14607
rect 16119 14727 16153 14743
rect 16119 14709 16153 14727
rect 16017 14505 16051 14539
rect 16200 14582 16222 14607
rect 16222 14582 16234 14607
rect 16200 14573 16234 14582
rect 16293 14601 16327 14607
rect 16293 14573 16324 14601
rect 16324 14573 16327 14601
rect 4977 14335 5011 14369
rect 5069 14335 5103 14369
rect 5161 14335 5195 14369
rect 5253 14335 5287 14369
rect 5345 14335 5379 14369
rect 5437 14335 5471 14369
rect 5529 14335 5563 14369
rect 5621 14335 5655 14369
rect 5713 14335 5747 14369
rect 5805 14335 5839 14369
rect 5897 14335 5931 14369
rect 5989 14335 6023 14369
rect 6081 14335 6115 14369
rect 6173 14335 6207 14369
rect 6265 14335 6299 14369
rect 6357 14335 6391 14369
rect 6449 14335 6483 14369
rect 6541 14335 6575 14369
rect 6633 14335 6667 14369
rect 6725 14335 6759 14369
rect 6817 14335 6851 14369
rect 6909 14335 6943 14369
rect 7001 14335 7035 14369
rect 7093 14335 7127 14369
rect 7185 14335 7219 14369
rect 7277 14335 7311 14369
rect 7369 14335 7403 14369
rect 7461 14335 7495 14369
rect 7553 14335 7587 14369
rect 7645 14335 7679 14369
rect 7737 14335 7771 14369
rect 7829 14335 7863 14369
rect 7921 14335 7955 14369
rect 8013 14335 8047 14369
rect 8105 14335 8139 14369
rect 8197 14335 8231 14369
rect 8289 14335 8323 14369
rect 8381 14335 8415 14369
rect 8473 14335 8507 14369
rect 8565 14335 8599 14369
rect 8657 14335 8691 14369
rect 8749 14335 8783 14369
rect 8841 14335 8875 14369
rect 8933 14335 8967 14369
rect 9025 14335 9059 14369
rect 9117 14335 9151 14369
rect 9209 14335 9243 14369
rect 9301 14335 9335 14369
rect 9393 14335 9427 14369
rect 9485 14335 9519 14369
rect 9577 14335 9611 14369
rect 9669 14335 9703 14369
rect 9761 14335 9795 14369
rect 9853 14335 9887 14369
rect 9945 14335 9979 14369
rect 10037 14335 10071 14369
rect 10129 14335 10163 14369
rect 10221 14335 10255 14369
rect 10313 14335 10347 14369
rect 10405 14335 10439 14369
rect 10497 14335 10531 14369
rect 10589 14335 10623 14369
rect 10681 14335 10715 14369
rect 10773 14335 10807 14369
rect 10865 14335 10899 14369
rect 10957 14335 10991 14369
rect 11049 14335 11083 14369
rect 11141 14335 11175 14369
rect 11233 14335 11267 14369
rect 11325 14335 11359 14369
rect 11417 14335 11451 14369
rect 11509 14335 11543 14369
rect 11601 14335 11635 14369
rect 11693 14335 11727 14369
rect 11785 14335 11819 14369
rect 11877 14335 11911 14369
rect 11969 14335 12003 14369
rect 12061 14335 12095 14369
rect 12153 14335 12187 14369
rect 12245 14335 12279 14369
rect 12337 14335 12371 14369
rect 12429 14335 12463 14369
rect 12521 14335 12555 14369
rect 12613 14335 12647 14369
rect 12705 14335 12739 14369
rect 12797 14335 12831 14369
rect 12889 14335 12923 14369
rect 12981 14335 13015 14369
rect 13073 14335 13107 14369
rect 13165 14335 13199 14369
rect 13257 14335 13291 14369
rect 13349 14335 13383 14369
rect 13441 14335 13475 14369
rect 13533 14335 13567 14369
rect 13625 14335 13659 14369
rect 13717 14335 13751 14369
rect 13809 14335 13843 14369
rect 13901 14335 13935 14369
rect 13993 14335 14027 14369
rect 14085 14335 14119 14369
rect 14177 14335 14211 14369
rect 14269 14335 14303 14369
rect 14361 14335 14395 14369
rect 14453 14335 14487 14369
rect 14545 14335 14579 14369
rect 14637 14335 14671 14369
rect 14729 14335 14763 14369
rect 14821 14335 14855 14369
rect 14913 14335 14947 14369
rect 15005 14335 15039 14369
rect 15097 14335 15131 14369
rect 15189 14335 15223 14369
rect 15281 14335 15315 14369
rect 15373 14335 15407 14369
rect 15465 14335 15499 14369
rect 15557 14335 15591 14369
rect 15649 14335 15683 14369
rect 15741 14335 15775 14369
rect 15833 14335 15867 14369
rect 15925 14335 15959 14369
rect 16017 14335 16051 14369
rect 16109 14335 16143 14369
rect 16201 14335 16235 14369
rect 16293 14335 16327 14369
rect 16385 14335 16419 14369
rect 16477 14335 16511 14369
rect 16569 14335 16603 14369
rect 16661 14335 16695 14369
rect 16753 14335 16787 14369
rect 16845 14335 16879 14369
rect 16937 14335 16971 14369
rect 17029 14335 17063 14369
rect 17121 14335 17155 14369
rect 17213 14335 17247 14369
rect 17305 14335 17339 14369
rect 17397 14335 17431 14369
rect 17489 14335 17523 14369
rect 17581 14335 17615 14369
rect 17673 14335 17707 14369
rect 17765 14335 17799 14369
rect 17857 14335 17891 14369
rect 17949 14335 17983 14369
rect 18041 14335 18075 14369
rect 18133 14335 18167 14369
rect 18225 14335 18259 14369
rect 18317 14335 18351 14369
rect 18409 14335 18443 14369
rect 18501 14335 18535 14369
rect 18593 14335 18627 14369
rect 18685 14335 18719 14369
rect 18777 14335 18811 14369
rect 18869 14335 18903 14369
rect 18961 14335 18995 14369
rect 19053 14335 19087 14369
rect 19145 14335 19179 14369
rect 19237 14335 19271 14369
rect 19329 14335 19363 14369
rect 19421 14335 19455 14369
rect 19513 14335 19547 14369
rect 19605 14335 19639 14369
rect 19697 14335 19731 14369
rect 19789 14335 19823 14369
rect 19881 14335 19915 14369
rect 19973 14335 20007 14369
rect 20065 14335 20099 14369
rect 20157 14335 20191 14369
rect 10425 14165 10459 14199
rect 10485 14111 10503 14136
rect 10503 14111 10519 14136
rect 10485 14102 10519 14111
rect 10129 13903 10135 13927
rect 10135 13903 10163 13927
rect 10129 13893 10163 13903
rect 10701 14113 10709 14131
rect 10709 14113 10735 14131
rect 10701 14097 10735 14113
rect 11073 14183 11107 14199
rect 11073 14165 11083 14183
rect 11083 14165 11107 14183
rect 11145 14165 11179 14199
rect 10701 13987 10704 13995
rect 10704 13987 10735 13995
rect 10701 13961 10735 13987
rect 11417 14097 11451 14131
rect 11325 13961 11359 13995
rect 11601 14029 11635 14063
rect 11703 13977 11737 13995
rect 11703 13961 11737 13977
rect 11784 14122 11818 14131
rect 11784 14097 11806 14122
rect 11806 14097 11818 14122
rect 11877 14029 11911 14063
rect 12153 14103 12179 14131
rect 12179 14103 12187 14131
rect 12153 14097 12187 14103
rect 13993 14165 14027 14199
rect 11969 13990 12003 13995
rect 11969 13961 11975 13990
rect 11975 13961 12003 13990
rect 12705 13911 12732 13927
rect 12732 13911 12739 13927
rect 12705 13893 12739 13911
rect 14269 14029 14303 14063
rect 15189 14240 15195 14267
rect 15195 14240 15223 14267
rect 15189 14233 15223 14240
rect 14913 14097 14947 14131
rect 15557 14097 15591 14131
rect 15649 14233 15683 14267
rect 16017 14263 16051 14267
rect 16017 14233 16023 14263
rect 16023 14233 16051 14263
rect 15833 14060 15867 14063
rect 15833 14029 15853 14060
rect 15853 14029 15867 14060
rect 16201 14103 16227 14131
rect 16227 14103 16235 14131
rect 16201 14097 16235 14103
rect 16477 14103 16503 14131
rect 16503 14103 16511 14131
rect 16477 14097 16511 14103
rect 16293 13909 16327 13927
rect 16293 13893 16299 13909
rect 16299 13893 16327 13909
rect 4977 13791 5011 13825
rect 5069 13791 5103 13825
rect 5161 13791 5195 13825
rect 5253 13791 5287 13825
rect 5345 13791 5379 13825
rect 5437 13791 5471 13825
rect 5529 13791 5563 13825
rect 5621 13791 5655 13825
rect 5713 13791 5747 13825
rect 5805 13791 5839 13825
rect 5897 13791 5931 13825
rect 5989 13791 6023 13825
rect 6081 13791 6115 13825
rect 6173 13791 6207 13825
rect 6265 13791 6299 13825
rect 6357 13791 6391 13825
rect 6449 13791 6483 13825
rect 6541 13791 6575 13825
rect 6633 13791 6667 13825
rect 6725 13791 6759 13825
rect 6817 13791 6851 13825
rect 6909 13791 6943 13825
rect 7001 13791 7035 13825
rect 7093 13791 7127 13825
rect 7185 13791 7219 13825
rect 7277 13791 7311 13825
rect 7369 13791 7403 13825
rect 7461 13791 7495 13825
rect 7553 13791 7587 13825
rect 7645 13791 7679 13825
rect 7737 13791 7771 13825
rect 7829 13791 7863 13825
rect 7921 13791 7955 13825
rect 8013 13791 8047 13825
rect 8105 13791 8139 13825
rect 8197 13791 8231 13825
rect 8289 13791 8323 13825
rect 8381 13791 8415 13825
rect 8473 13791 8507 13825
rect 8565 13791 8599 13825
rect 8657 13791 8691 13825
rect 8749 13791 8783 13825
rect 8841 13791 8875 13825
rect 8933 13791 8967 13825
rect 9025 13791 9059 13825
rect 9117 13791 9151 13825
rect 9209 13791 9243 13825
rect 9301 13791 9335 13825
rect 9393 13791 9427 13825
rect 9485 13791 9519 13825
rect 9577 13791 9611 13825
rect 9669 13791 9703 13825
rect 9761 13791 9795 13825
rect 9853 13791 9887 13825
rect 9945 13791 9979 13825
rect 10037 13791 10071 13825
rect 10129 13791 10163 13825
rect 10221 13791 10255 13825
rect 10313 13791 10347 13825
rect 10405 13791 10439 13825
rect 10497 13791 10531 13825
rect 10589 13791 10623 13825
rect 10681 13791 10715 13825
rect 10773 13791 10807 13825
rect 10865 13791 10899 13825
rect 10957 13791 10991 13825
rect 11049 13791 11083 13825
rect 11141 13791 11175 13825
rect 11233 13791 11267 13825
rect 11325 13791 11359 13825
rect 11417 13791 11451 13825
rect 11509 13791 11543 13825
rect 11601 13791 11635 13825
rect 11693 13791 11727 13825
rect 11785 13791 11819 13825
rect 11877 13791 11911 13825
rect 11969 13791 12003 13825
rect 12061 13791 12095 13825
rect 12153 13791 12187 13825
rect 12245 13791 12279 13825
rect 12337 13791 12371 13825
rect 12429 13791 12463 13825
rect 12521 13791 12555 13825
rect 12613 13791 12647 13825
rect 12705 13791 12739 13825
rect 12797 13791 12831 13825
rect 12889 13791 12923 13825
rect 12981 13791 13015 13825
rect 13073 13791 13107 13825
rect 13165 13791 13199 13825
rect 13257 13791 13291 13825
rect 13349 13791 13383 13825
rect 13441 13791 13475 13825
rect 13533 13791 13567 13825
rect 13625 13791 13659 13825
rect 13717 13791 13751 13825
rect 13809 13791 13843 13825
rect 13901 13791 13935 13825
rect 13993 13791 14027 13825
rect 14085 13791 14119 13825
rect 14177 13791 14211 13825
rect 14269 13791 14303 13825
rect 14361 13791 14395 13825
rect 14453 13791 14487 13825
rect 14545 13791 14579 13825
rect 14637 13791 14671 13825
rect 14729 13791 14763 13825
rect 14821 13791 14855 13825
rect 14913 13791 14947 13825
rect 15005 13791 15039 13825
rect 15097 13791 15131 13825
rect 15189 13791 15223 13825
rect 15281 13791 15315 13825
rect 15373 13791 15407 13825
rect 15465 13791 15499 13825
rect 15557 13791 15591 13825
rect 15649 13791 15683 13825
rect 15741 13791 15775 13825
rect 15833 13791 15867 13825
rect 15925 13791 15959 13825
rect 16017 13791 16051 13825
rect 16109 13791 16143 13825
rect 16201 13791 16235 13825
rect 16293 13791 16327 13825
rect 16385 13791 16419 13825
rect 16477 13791 16511 13825
rect 16569 13791 16603 13825
rect 16661 13791 16695 13825
rect 16753 13791 16787 13825
rect 16845 13791 16879 13825
rect 16937 13791 16971 13825
rect 17029 13791 17063 13825
rect 17121 13791 17155 13825
rect 17213 13791 17247 13825
rect 17305 13791 17339 13825
rect 17397 13791 17431 13825
rect 17489 13791 17523 13825
rect 17581 13791 17615 13825
rect 17673 13791 17707 13825
rect 17765 13791 17799 13825
rect 17857 13791 17891 13825
rect 17949 13791 17983 13825
rect 18041 13791 18075 13825
rect 18133 13791 18167 13825
rect 18225 13791 18259 13825
rect 18317 13791 18351 13825
rect 18409 13791 18443 13825
rect 18501 13791 18535 13825
rect 18593 13791 18627 13825
rect 18685 13791 18719 13825
rect 18777 13791 18811 13825
rect 18869 13791 18903 13825
rect 18961 13791 18995 13825
rect 19053 13791 19087 13825
rect 19145 13791 19179 13825
rect 19237 13791 19271 13825
rect 19329 13791 19363 13825
rect 19421 13791 19455 13825
rect 19513 13791 19547 13825
rect 19605 13791 19639 13825
rect 19697 13791 19731 13825
rect 19789 13791 19823 13825
rect 19881 13791 19915 13825
rect 19973 13791 20007 13825
rect 20065 13791 20099 13825
rect 20157 13791 20191 13825
rect 9669 13513 9703 13519
rect 9669 13485 9677 13513
rect 9677 13485 9703 13513
rect 10405 13705 10439 13723
rect 10405 13689 10432 13705
rect 10432 13689 10439 13705
rect 9853 13353 9881 13383
rect 9881 13353 9887 13383
rect 9853 13349 9887 13353
rect 11693 13513 11727 13519
rect 11693 13485 11719 13513
rect 11719 13485 11727 13513
rect 12889 13713 12923 13723
rect 12889 13689 12895 13713
rect 12895 13689 12923 13713
rect 12705 13513 12739 13519
rect 12705 13485 12731 13513
rect 12731 13485 12739 13513
rect 12521 13353 12527 13383
rect 12527 13353 12555 13383
rect 12521 13349 12555 13353
rect 13461 13629 13495 13655
rect 13461 13621 13464 13629
rect 13464 13621 13495 13629
rect 13245 13505 13279 13514
rect 13245 13480 13263 13505
rect 13263 13480 13279 13505
rect 13185 13417 13219 13451
rect 13461 13503 13495 13519
rect 13461 13485 13469 13503
rect 13469 13485 13495 13503
rect 14085 13621 14119 13655
rect 13833 13433 13843 13451
rect 13843 13433 13867 13451
rect 13833 13417 13867 13433
rect 13905 13417 13939 13451
rect 14177 13485 14211 13519
rect 14463 13639 14497 13655
rect 14463 13621 14497 13639
rect 14361 13417 14395 13451
rect 14544 13494 14566 13519
rect 14566 13494 14578 13519
rect 14544 13485 14578 13494
rect 14637 13553 14671 13587
rect 16201 13705 16235 13723
rect 16201 13689 16230 13705
rect 16230 13689 16235 13705
rect 16569 13715 16575 13723
rect 16575 13715 16603 13723
rect 16569 13689 16603 13715
rect 14729 13513 14763 13519
rect 14729 13485 14737 13513
rect 14737 13485 14763 13513
rect 16937 13485 16971 13519
rect 17121 13553 17155 13587
rect 17029 13349 17063 13383
rect 4977 13247 5011 13281
rect 5069 13247 5103 13281
rect 5161 13247 5195 13281
rect 5253 13247 5287 13281
rect 5345 13247 5379 13281
rect 5437 13247 5471 13281
rect 5529 13247 5563 13281
rect 5621 13247 5655 13281
rect 5713 13247 5747 13281
rect 5805 13247 5839 13281
rect 5897 13247 5931 13281
rect 5989 13247 6023 13281
rect 6081 13247 6115 13281
rect 6173 13247 6207 13281
rect 6265 13247 6299 13281
rect 6357 13247 6391 13281
rect 6449 13247 6483 13281
rect 6541 13247 6575 13281
rect 6633 13247 6667 13281
rect 6725 13247 6759 13281
rect 6817 13247 6851 13281
rect 6909 13247 6943 13281
rect 7001 13247 7035 13281
rect 7093 13247 7127 13281
rect 7185 13247 7219 13281
rect 7277 13247 7311 13281
rect 7369 13247 7403 13281
rect 7461 13247 7495 13281
rect 7553 13247 7587 13281
rect 7645 13247 7679 13281
rect 7737 13247 7771 13281
rect 7829 13247 7863 13281
rect 7921 13247 7955 13281
rect 8013 13247 8047 13281
rect 8105 13247 8139 13281
rect 8197 13247 8231 13281
rect 8289 13247 8323 13281
rect 8381 13247 8415 13281
rect 8473 13247 8507 13281
rect 8565 13247 8599 13281
rect 8657 13247 8691 13281
rect 8749 13247 8783 13281
rect 8841 13247 8875 13281
rect 8933 13247 8967 13281
rect 9025 13247 9059 13281
rect 9117 13247 9151 13281
rect 9209 13247 9243 13281
rect 9301 13247 9335 13281
rect 9393 13247 9427 13281
rect 9485 13247 9519 13281
rect 9577 13247 9611 13281
rect 9669 13247 9703 13281
rect 9761 13247 9795 13281
rect 9853 13247 9887 13281
rect 9945 13247 9979 13281
rect 10037 13247 10071 13281
rect 10129 13247 10163 13281
rect 10221 13247 10255 13281
rect 10313 13247 10347 13281
rect 10405 13247 10439 13281
rect 10497 13247 10531 13281
rect 10589 13247 10623 13281
rect 10681 13247 10715 13281
rect 10773 13247 10807 13281
rect 10865 13247 10899 13281
rect 10957 13247 10991 13281
rect 11049 13247 11083 13281
rect 11141 13247 11175 13281
rect 11233 13247 11267 13281
rect 11325 13247 11359 13281
rect 11417 13247 11451 13281
rect 11509 13247 11543 13281
rect 11601 13247 11635 13281
rect 11693 13247 11727 13281
rect 11785 13247 11819 13281
rect 11877 13247 11911 13281
rect 11969 13247 12003 13281
rect 12061 13247 12095 13281
rect 12153 13247 12187 13281
rect 12245 13247 12279 13281
rect 12337 13247 12371 13281
rect 12429 13247 12463 13281
rect 12521 13247 12555 13281
rect 12613 13247 12647 13281
rect 12705 13247 12739 13281
rect 12797 13247 12831 13281
rect 12889 13247 12923 13281
rect 12981 13247 13015 13281
rect 13073 13247 13107 13281
rect 13165 13247 13199 13281
rect 13257 13247 13291 13281
rect 13349 13247 13383 13281
rect 13441 13247 13475 13281
rect 13533 13247 13567 13281
rect 13625 13247 13659 13281
rect 13717 13247 13751 13281
rect 13809 13247 13843 13281
rect 13901 13247 13935 13281
rect 13993 13247 14027 13281
rect 14085 13247 14119 13281
rect 14177 13247 14211 13281
rect 14269 13247 14303 13281
rect 14361 13247 14395 13281
rect 14453 13247 14487 13281
rect 14545 13247 14579 13281
rect 14637 13247 14671 13281
rect 14729 13247 14763 13281
rect 14821 13247 14855 13281
rect 14913 13247 14947 13281
rect 15005 13247 15039 13281
rect 15097 13247 15131 13281
rect 15189 13247 15223 13281
rect 15281 13247 15315 13281
rect 15373 13247 15407 13281
rect 15465 13247 15499 13281
rect 15557 13247 15591 13281
rect 15649 13247 15683 13281
rect 15741 13247 15775 13281
rect 15833 13247 15867 13281
rect 15925 13247 15959 13281
rect 16017 13247 16051 13281
rect 16109 13247 16143 13281
rect 16201 13247 16235 13281
rect 16293 13247 16327 13281
rect 16385 13247 16419 13281
rect 16477 13247 16511 13281
rect 16569 13247 16603 13281
rect 16661 13247 16695 13281
rect 16753 13247 16787 13281
rect 16845 13247 16879 13281
rect 16937 13247 16971 13281
rect 17029 13247 17063 13281
rect 17121 13247 17155 13281
rect 17213 13247 17247 13281
rect 17305 13247 17339 13281
rect 17397 13247 17431 13281
rect 17489 13247 17523 13281
rect 17581 13247 17615 13281
rect 17673 13247 17707 13281
rect 17765 13247 17799 13281
rect 17857 13247 17891 13281
rect 17949 13247 17983 13281
rect 18041 13247 18075 13281
rect 18133 13247 18167 13281
rect 18225 13247 18259 13281
rect 18317 13247 18351 13281
rect 18409 13247 18443 13281
rect 18501 13247 18535 13281
rect 18593 13247 18627 13281
rect 18685 13247 18719 13281
rect 18777 13247 18811 13281
rect 18869 13247 18903 13281
rect 18961 13247 18995 13281
rect 19053 13247 19087 13281
rect 19145 13247 19179 13281
rect 19237 13247 19271 13281
rect 19329 13247 19363 13281
rect 19421 13247 19455 13281
rect 19513 13247 19547 13281
rect 19605 13247 19639 13281
rect 19697 13247 19731 13281
rect 19789 13247 19823 13281
rect 19881 13247 19915 13281
rect 19973 13247 20007 13281
rect 20065 13247 20099 13281
rect 20157 13247 20191 13281
rect 9209 12941 9243 12975
rect 9761 12805 9770 12839
rect 9770 12805 9795 12839
rect 10701 13077 10735 13111
rect 10761 13023 10779 13048
rect 10779 13023 10795 13048
rect 10761 13014 10795 13023
rect 10405 12941 10439 12975
rect 10977 13025 10985 13043
rect 10985 13025 11011 13043
rect 10977 13009 11011 13025
rect 11349 13095 11383 13111
rect 11349 13077 11359 13095
rect 11359 13077 11383 13095
rect 11421 13077 11455 13111
rect 10977 12899 10980 12907
rect 10980 12899 11011 12907
rect 10977 12873 11011 12899
rect 11693 13009 11727 13043
rect 11601 12873 11635 12907
rect 11877 12941 11911 12975
rect 11979 12889 12013 12907
rect 11979 12873 12013 12889
rect 12060 13034 12094 13043
rect 12060 13009 12082 13034
rect 12082 13009 12094 13034
rect 12153 13015 12184 13043
rect 12184 13015 12187 13043
rect 12153 13009 12187 13015
rect 12245 13015 12248 13043
rect 12248 13015 12279 13043
rect 12245 13009 12279 13015
rect 12338 13034 12372 13043
rect 12338 13009 12350 13034
rect 12350 13009 12372 13034
rect 12521 12941 12555 12975
rect 12419 12889 12453 12907
rect 12419 12873 12453 12889
rect 12705 13009 12739 13043
rect 12977 13077 13011 13111
rect 13049 13095 13083 13111
rect 13049 13077 13073 13095
rect 13073 13077 13083 13095
rect 12797 12873 12831 12907
rect 13421 13025 13447 13043
rect 13447 13025 13455 13043
rect 13421 13009 13455 13025
rect 13697 13077 13731 13111
rect 13637 13023 13653 13048
rect 13653 13023 13671 13048
rect 13637 13014 13671 13023
rect 13421 12899 13452 12907
rect 13452 12899 13455 12907
rect 13421 12873 13455 12899
rect 13993 12815 14021 12839
rect 14021 12815 14027 12839
rect 13993 12805 14027 12815
rect 14085 12881 14119 12907
rect 14085 12873 14091 12881
rect 14091 12873 14119 12881
rect 14453 13009 14487 13043
rect 14545 13077 14579 13111
rect 14729 12972 14763 12975
rect 14729 12941 14749 12972
rect 14749 12941 14763 12972
rect 15393 13077 15427 13111
rect 15453 13023 15471 13048
rect 15471 13023 15487 13048
rect 15453 13014 15487 13023
rect 15097 12815 15103 12839
rect 15103 12815 15131 12839
rect 15097 12805 15131 12815
rect 15669 13025 15677 13043
rect 15677 13025 15703 13043
rect 15669 13009 15703 13025
rect 16041 13095 16075 13111
rect 16041 13077 16051 13095
rect 16051 13077 16075 13095
rect 16113 13077 16147 13111
rect 15669 12899 15672 12907
rect 15672 12899 15703 12907
rect 15669 12873 15703 12899
rect 16385 13009 16419 13043
rect 16293 12873 16327 12907
rect 16569 12941 16603 12975
rect 16671 12889 16705 12907
rect 16671 12873 16705 12889
rect 16937 13145 16962 13179
rect 16962 13145 16971 13179
rect 16752 13034 16786 13043
rect 16752 13009 16774 13034
rect 16774 13009 16786 13034
rect 16845 13015 16876 13043
rect 16876 13015 16879 13043
rect 16845 13009 16879 13015
rect 17581 12941 17615 12975
rect 4977 12703 5011 12737
rect 5069 12703 5103 12737
rect 5161 12703 5195 12737
rect 5253 12703 5287 12737
rect 5345 12703 5379 12737
rect 5437 12703 5471 12737
rect 5529 12703 5563 12737
rect 5621 12703 5655 12737
rect 5713 12703 5747 12737
rect 5805 12703 5839 12737
rect 5897 12703 5931 12737
rect 5989 12703 6023 12737
rect 6081 12703 6115 12737
rect 6173 12703 6207 12737
rect 6265 12703 6299 12737
rect 6357 12703 6391 12737
rect 6449 12703 6483 12737
rect 6541 12703 6575 12737
rect 6633 12703 6667 12737
rect 6725 12703 6759 12737
rect 6817 12703 6851 12737
rect 6909 12703 6943 12737
rect 7001 12703 7035 12737
rect 7093 12703 7127 12737
rect 7185 12703 7219 12737
rect 7277 12703 7311 12737
rect 7369 12703 7403 12737
rect 7461 12703 7495 12737
rect 7553 12703 7587 12737
rect 7645 12703 7679 12737
rect 7737 12703 7771 12737
rect 7829 12703 7863 12737
rect 7921 12703 7955 12737
rect 8013 12703 8047 12737
rect 8105 12703 8139 12737
rect 8197 12703 8231 12737
rect 8289 12703 8323 12737
rect 8381 12703 8415 12737
rect 8473 12703 8507 12737
rect 8565 12703 8599 12737
rect 8657 12703 8691 12737
rect 8749 12703 8783 12737
rect 8841 12703 8875 12737
rect 8933 12703 8967 12737
rect 9025 12703 9059 12737
rect 9117 12703 9151 12737
rect 9209 12703 9243 12737
rect 9301 12703 9335 12737
rect 9393 12703 9427 12737
rect 9485 12703 9519 12737
rect 9577 12703 9611 12737
rect 9669 12703 9703 12737
rect 9761 12703 9795 12737
rect 9853 12703 9887 12737
rect 9945 12703 9979 12737
rect 10037 12703 10071 12737
rect 10129 12703 10163 12737
rect 10221 12703 10255 12737
rect 10313 12703 10347 12737
rect 10405 12703 10439 12737
rect 10497 12703 10531 12737
rect 10589 12703 10623 12737
rect 10681 12703 10715 12737
rect 10773 12703 10807 12737
rect 10865 12703 10899 12737
rect 10957 12703 10991 12737
rect 11049 12703 11083 12737
rect 11141 12703 11175 12737
rect 11233 12703 11267 12737
rect 11325 12703 11359 12737
rect 11417 12703 11451 12737
rect 11509 12703 11543 12737
rect 11601 12703 11635 12737
rect 11693 12703 11727 12737
rect 11785 12703 11819 12737
rect 11877 12703 11911 12737
rect 11969 12703 12003 12737
rect 12061 12703 12095 12737
rect 12153 12703 12187 12737
rect 12245 12703 12279 12737
rect 12337 12703 12371 12737
rect 12429 12703 12463 12737
rect 12521 12703 12555 12737
rect 12613 12703 12647 12737
rect 12705 12703 12739 12737
rect 12797 12703 12831 12737
rect 12889 12703 12923 12737
rect 12981 12703 13015 12737
rect 13073 12703 13107 12737
rect 13165 12703 13199 12737
rect 13257 12703 13291 12737
rect 13349 12703 13383 12737
rect 13441 12703 13475 12737
rect 13533 12703 13567 12737
rect 13625 12703 13659 12737
rect 13717 12703 13751 12737
rect 13809 12703 13843 12737
rect 13901 12703 13935 12737
rect 13993 12703 14027 12737
rect 14085 12703 14119 12737
rect 14177 12703 14211 12737
rect 14269 12703 14303 12737
rect 14361 12703 14395 12737
rect 14453 12703 14487 12737
rect 14545 12703 14579 12737
rect 14637 12703 14671 12737
rect 14729 12703 14763 12737
rect 14821 12703 14855 12737
rect 14913 12703 14947 12737
rect 15005 12703 15039 12737
rect 15097 12703 15131 12737
rect 15189 12703 15223 12737
rect 15281 12703 15315 12737
rect 15373 12703 15407 12737
rect 15465 12703 15499 12737
rect 15557 12703 15591 12737
rect 15649 12703 15683 12737
rect 15741 12703 15775 12737
rect 15833 12703 15867 12737
rect 15925 12703 15959 12737
rect 16017 12703 16051 12737
rect 16109 12703 16143 12737
rect 16201 12703 16235 12737
rect 16293 12703 16327 12737
rect 16385 12703 16419 12737
rect 16477 12703 16511 12737
rect 16569 12703 16603 12737
rect 16661 12703 16695 12737
rect 16753 12703 16787 12737
rect 16845 12703 16879 12737
rect 16937 12703 16971 12737
rect 17029 12703 17063 12737
rect 17121 12703 17155 12737
rect 17213 12703 17247 12737
rect 17305 12703 17339 12737
rect 17397 12703 17431 12737
rect 17489 12703 17523 12737
rect 17581 12703 17615 12737
rect 17673 12703 17707 12737
rect 17765 12703 17799 12737
rect 17857 12703 17891 12737
rect 17949 12703 17983 12737
rect 18041 12703 18075 12737
rect 18133 12703 18167 12737
rect 18225 12703 18259 12737
rect 18317 12703 18351 12737
rect 18409 12703 18443 12737
rect 18501 12703 18535 12737
rect 18593 12703 18627 12737
rect 18685 12703 18719 12737
rect 18777 12703 18811 12737
rect 18869 12703 18903 12737
rect 18961 12703 18995 12737
rect 19053 12703 19087 12737
rect 19145 12703 19179 12737
rect 19237 12703 19271 12737
rect 19329 12703 19363 12737
rect 19421 12703 19455 12737
rect 19513 12703 19547 12737
rect 19605 12703 19639 12737
rect 19697 12703 19731 12737
rect 19789 12703 19823 12737
rect 19881 12703 19915 12737
rect 19973 12703 20007 12737
rect 20065 12703 20099 12737
rect 20157 12703 20191 12737
rect 5253 12397 5287 12431
rect 7093 12329 7127 12363
rect 7001 12261 7030 12295
rect 7030 12261 7035 12295
rect 9209 12397 9243 12431
rect 9117 12261 9146 12295
rect 9146 12261 9151 12295
rect 10221 12626 10255 12635
rect 10221 12601 10251 12626
rect 10251 12601 10255 12626
rect 10313 12329 10347 12363
rect 10497 12559 10503 12567
rect 10503 12559 10531 12567
rect 10497 12533 10531 12559
rect 10957 12468 10959 12499
rect 10959 12468 10991 12499
rect 10957 12465 10991 12468
rect 10865 12397 10899 12431
rect 11141 12468 11161 12499
rect 11161 12468 11175 12499
rect 11141 12465 11175 12468
rect 11601 12465 11635 12499
rect 11693 12261 11727 12295
rect 11785 12397 11819 12431
rect 12153 12627 12181 12635
rect 12181 12627 12187 12635
rect 12153 12601 12187 12627
rect 13073 12397 13107 12431
rect 12981 12261 13010 12295
rect 13010 12261 13015 12295
rect 13993 12619 14021 12635
rect 14021 12619 14027 12635
rect 13993 12601 14027 12619
rect 13349 12397 13383 12431
rect 13809 12425 13843 12431
rect 13809 12397 13817 12425
rect 13817 12397 13843 12425
rect 13625 12261 13652 12295
rect 13652 12261 13659 12295
rect 14177 12465 14211 12499
rect 14729 12601 14738 12635
rect 14738 12601 14763 12635
rect 15097 12465 15131 12499
rect 15190 12406 15202 12431
rect 15202 12406 15224 12431
rect 15190 12397 15224 12406
rect 15271 12551 15305 12567
rect 15271 12533 15305 12551
rect 15373 12465 15407 12499
rect 15649 12533 15683 12567
rect 15557 12397 15591 12431
rect 16273 12541 16307 12567
rect 16273 12533 16304 12541
rect 16304 12533 16307 12541
rect 15829 12329 15863 12363
rect 15901 12345 15925 12363
rect 15925 12345 15935 12363
rect 15901 12329 15935 12345
rect 16273 12415 16307 12431
rect 16273 12397 16299 12415
rect 16299 12397 16307 12415
rect 16845 12465 16879 12499
rect 16489 12417 16523 12426
rect 16489 12392 16505 12417
rect 16505 12392 16523 12417
rect 16549 12329 16583 12363
rect 17121 12397 17155 12431
rect 17489 12329 17523 12363
rect 19513 12397 19547 12431
rect 19881 12329 19915 12363
rect 4977 12159 5011 12193
rect 5069 12159 5103 12193
rect 5161 12159 5195 12193
rect 5253 12159 5287 12193
rect 5345 12159 5379 12193
rect 5437 12159 5471 12193
rect 5529 12159 5563 12193
rect 5621 12159 5655 12193
rect 5713 12159 5747 12193
rect 5805 12159 5839 12193
rect 5897 12159 5931 12193
rect 5989 12159 6023 12193
rect 6081 12159 6115 12193
rect 6173 12159 6207 12193
rect 6265 12159 6299 12193
rect 6357 12159 6391 12193
rect 6449 12159 6483 12193
rect 6541 12159 6575 12193
rect 6633 12159 6667 12193
rect 6725 12159 6759 12193
rect 6817 12159 6851 12193
rect 6909 12159 6943 12193
rect 7001 12159 7035 12193
rect 7093 12159 7127 12193
rect 7185 12159 7219 12193
rect 7277 12159 7311 12193
rect 7369 12159 7403 12193
rect 7461 12159 7495 12193
rect 7553 12159 7587 12193
rect 7645 12159 7679 12193
rect 7737 12159 7771 12193
rect 7829 12159 7863 12193
rect 7921 12159 7955 12193
rect 8013 12159 8047 12193
rect 8105 12159 8139 12193
rect 8197 12159 8231 12193
rect 8289 12159 8323 12193
rect 8381 12159 8415 12193
rect 8473 12159 8507 12193
rect 8565 12159 8599 12193
rect 8657 12159 8691 12193
rect 8749 12159 8783 12193
rect 8841 12159 8875 12193
rect 8933 12159 8967 12193
rect 9025 12159 9059 12193
rect 9117 12159 9151 12193
rect 9209 12159 9243 12193
rect 9301 12159 9335 12193
rect 9393 12159 9427 12193
rect 9485 12159 9519 12193
rect 9577 12159 9611 12193
rect 9669 12159 9703 12193
rect 9761 12159 9795 12193
rect 9853 12159 9887 12193
rect 9945 12159 9979 12193
rect 10037 12159 10071 12193
rect 10129 12159 10163 12193
rect 10221 12159 10255 12193
rect 10313 12159 10347 12193
rect 10405 12159 10439 12193
rect 10497 12159 10531 12193
rect 10589 12159 10623 12193
rect 10681 12159 10715 12193
rect 10773 12159 10807 12193
rect 10865 12159 10899 12193
rect 10957 12159 10991 12193
rect 11049 12159 11083 12193
rect 11141 12159 11175 12193
rect 11233 12159 11267 12193
rect 11325 12159 11359 12193
rect 11417 12159 11451 12193
rect 11509 12159 11543 12193
rect 11601 12159 11635 12193
rect 11693 12159 11727 12193
rect 11785 12159 11819 12193
rect 11877 12159 11911 12193
rect 11969 12159 12003 12193
rect 12061 12159 12095 12193
rect 12153 12159 12187 12193
rect 12245 12159 12279 12193
rect 12337 12159 12371 12193
rect 12429 12159 12463 12193
rect 12521 12159 12555 12193
rect 12613 12159 12647 12193
rect 12705 12159 12739 12193
rect 12797 12159 12831 12193
rect 12889 12159 12923 12193
rect 12981 12159 13015 12193
rect 13073 12159 13107 12193
rect 13165 12159 13199 12193
rect 13257 12159 13291 12193
rect 13349 12159 13383 12193
rect 13441 12159 13475 12193
rect 13533 12159 13567 12193
rect 13625 12159 13659 12193
rect 13717 12159 13751 12193
rect 13809 12159 13843 12193
rect 13901 12159 13935 12193
rect 13993 12159 14027 12193
rect 14085 12159 14119 12193
rect 14177 12159 14211 12193
rect 14269 12159 14303 12193
rect 14361 12159 14395 12193
rect 14453 12159 14487 12193
rect 14545 12159 14579 12193
rect 14637 12159 14671 12193
rect 14729 12159 14763 12193
rect 14821 12159 14855 12193
rect 14913 12159 14947 12193
rect 15005 12159 15039 12193
rect 15097 12159 15131 12193
rect 15189 12159 15223 12193
rect 15281 12159 15315 12193
rect 15373 12159 15407 12193
rect 15465 12159 15499 12193
rect 15557 12159 15591 12193
rect 15649 12159 15683 12193
rect 15741 12159 15775 12193
rect 15833 12159 15867 12193
rect 15925 12159 15959 12193
rect 16017 12159 16051 12193
rect 16109 12159 16143 12193
rect 16201 12159 16235 12193
rect 16293 12159 16327 12193
rect 16385 12159 16419 12193
rect 16477 12159 16511 12193
rect 16569 12159 16603 12193
rect 16661 12159 16695 12193
rect 16753 12159 16787 12193
rect 16845 12159 16879 12193
rect 16937 12159 16971 12193
rect 17029 12159 17063 12193
rect 17121 12159 17155 12193
rect 17213 12159 17247 12193
rect 17305 12159 17339 12193
rect 17397 12159 17431 12193
rect 17489 12159 17523 12193
rect 17581 12159 17615 12193
rect 17673 12159 17707 12193
rect 17765 12159 17799 12193
rect 17857 12159 17891 12193
rect 17949 12159 17983 12193
rect 18041 12159 18075 12193
rect 18133 12159 18167 12193
rect 18225 12159 18259 12193
rect 18317 12159 18351 12193
rect 18409 12159 18443 12193
rect 18501 12159 18535 12193
rect 18593 12159 18627 12193
rect 18685 12159 18719 12193
rect 18777 12159 18811 12193
rect 18869 12159 18903 12193
rect 18961 12159 18995 12193
rect 19053 12159 19087 12193
rect 19145 12159 19179 12193
rect 19237 12159 19271 12193
rect 19329 12159 19363 12193
rect 19421 12159 19455 12193
rect 19513 12159 19547 12193
rect 19605 12159 19639 12193
rect 19697 12159 19731 12193
rect 19789 12159 19823 12193
rect 19881 12159 19915 12193
rect 19973 12159 20007 12193
rect 20065 12159 20099 12193
rect 20157 12159 20191 12193
rect 25862 8679 25900 9076
rect 26180 8679 26218 9076
rect 26498 8679 26536 9076
rect 26816 8679 26854 9076
rect 27134 8679 27172 9076
rect 27452 8679 27490 9076
rect 27770 8679 27808 9076
rect 28088 8679 28126 9076
rect 25862 7164 25900 7561
rect 26180 7164 26218 7561
rect 26498 7164 26536 7561
rect 26816 7164 26854 7561
rect 27134 7164 27172 7561
rect 27452 7164 27490 7561
rect 27770 7164 27808 7561
rect 28088 7164 28126 7561
rect 29780 7010 30380 7050
rect 3532 5455 3570 5852
rect 3532 4824 3570 5221
rect 6832 5359 6870 5756
rect 6832 4824 6870 5221
rect 10132 5499 10170 5896
rect 10132 4824 10170 5221
rect 13432 5779 13470 6176
rect 13432 4824 13470 5221
rect 17032 6339 17070 6736
rect 17032 4824 17070 5221
rect 20232 6339 20270 6736
rect 20550 6339 20588 6736
rect 20232 4824 20270 5221
rect 20550 4824 20588 5221
rect 23332 6339 23370 6736
rect 23650 6339 23688 6736
rect 23968 6339 24006 6736
rect 24286 6339 24324 6736
rect 23332 4824 23370 5221
rect 23650 4824 23688 5221
rect 23968 4824 24006 5221
rect 24286 4824 24324 5221
rect 25832 6339 25870 6736
rect 26150 6339 26188 6736
rect 26468 6339 26506 6736
rect 26786 6339 26824 6736
rect 27104 6339 27142 6736
rect 27422 6339 27460 6736
rect 27740 6339 27778 6736
rect 28058 6339 28096 6736
rect 25832 4824 25870 5221
rect 26150 4824 26188 5221
rect 26468 4824 26506 5221
rect 26786 4824 26824 5221
rect 27104 4824 27142 5221
rect 27422 4824 27460 5221
rect 27740 4824 27778 5221
rect 28058 4824 28096 5221
rect 29830 6797 29998 6831
rect 30210 6797 30378 6831
rect 30468 6797 30636 6831
rect 30850 6797 31018 6831
rect 31108 6797 31276 6831
rect 31366 6797 31534 6831
rect 31750 6797 31918 6831
rect 32008 6797 32176 6831
rect 32266 6797 32434 6831
rect 32524 6797 32692 6831
rect 32782 6797 32950 6831
rect 33040 6797 33208 6831
rect 33298 6797 33466 6831
rect 33556 6797 33724 6831
rect 33814 6797 33982 6831
rect 34072 6797 34240 6831
rect 34450 6797 34618 6831
rect 29768 6162 29802 6738
rect 30026 6162 30060 6738
rect 30148 6433 30182 6721
rect 30406 6179 30440 6467
rect 30664 6433 30698 6721
rect 30788 6433 30822 6721
rect 31046 6179 31080 6467
rect 31304 6433 31338 6721
rect 31562 6179 31596 6467
rect 31688 6433 31722 6721
rect 31946 6179 31980 6467
rect 32204 6433 32238 6721
rect 32462 6179 32496 6467
rect 32720 6433 32754 6721
rect 32978 6179 33012 6467
rect 33236 6433 33270 6721
rect 33494 6179 33528 6467
rect 33752 6433 33786 6721
rect 34010 6179 34044 6467
rect 34268 6433 34302 6721
rect 34388 6162 34422 6738
rect 34646 6162 34680 6738
rect 29830 6069 29998 6103
rect 30210 6069 30378 6103
rect 30468 6069 30636 6103
rect 30850 6069 31018 6103
rect 31108 6069 31276 6103
rect 31366 6069 31534 6103
rect 31750 6069 31918 6103
rect 32008 6069 32176 6103
rect 32266 6069 32434 6103
rect 32524 6069 32692 6103
rect 32782 6069 32950 6103
rect 33040 6069 33208 6103
rect 33298 6069 33466 6103
rect 33556 6069 33724 6103
rect 33814 6069 33982 6103
rect 34072 6069 34240 6103
rect 34450 6069 34618 6103
rect 30072 5777 30106 5811
rect 30392 5777 30426 5811
rect 30792 5777 30826 5811
rect 31092 5777 31126 5811
rect 30028 5413 30062 5701
rect 30116 5413 30150 5701
rect 30248 5413 30282 5701
rect 30344 5159 30378 5447
rect 30440 5413 30474 5701
rect 30536 5159 30570 5447
rect 30648 5159 30682 5447
rect 30744 5413 30778 5701
rect 30840 5159 30874 5447
rect 30936 5413 30970 5701
rect 31048 5413 31082 5701
rect 31136 5413 31170 5701
rect 30072 5049 30106 5083
rect 30296 5049 30330 5083
rect 30488 5049 30522 5083
rect 30696 5049 30730 5083
rect 30888 5049 30922 5083
rect 31092 5049 31126 5083
rect 1482 4277 1516 4311
rect 1995 4270 2029 4304
rect 2187 4270 2221 4304
rect 2379 4270 2413 4304
rect 2571 4270 2605 4304
rect 2763 4270 2797 4304
rect 2955 4270 2989 4304
rect 3182 4277 3216 4311
rect 1310 3490 1350 3580
rect 1350 3490 1360 3580
rect 1438 3713 1472 4201
rect 1526 3713 1560 4201
rect 1682 3877 1716 3911
rect 1638 3242 1672 3818
rect 1726 3242 1760 3818
rect 1851 3706 1885 4194
rect 1947 3252 1981 3740
rect 2043 3706 2077 4194
rect 2139 3252 2173 3740
rect 2235 3706 2269 4194
rect 2331 3252 2365 3740
rect 2427 3706 2461 4194
rect 2523 3252 2557 3740
rect 2619 3706 2653 4194
rect 2715 3252 2749 3740
rect 2811 3706 2845 4194
rect 2907 3252 2941 3740
rect 3003 3706 3037 4194
rect 3138 3242 3172 4218
rect 3226 3242 3260 4218
rect 1482 3149 1516 3183
rect 1682 3149 1716 3183
rect 1899 3142 1933 3176
rect 2091 3142 2125 3176
rect 2283 3142 2317 3176
rect 2475 3142 2509 3176
rect 2667 3142 2701 3176
rect 2859 3142 2893 3176
rect 3182 3149 3216 3183
rect 4782 4277 4816 4311
rect 5295 4270 5329 4304
rect 5487 4270 5521 4304
rect 5679 4270 5713 4304
rect 5871 4270 5905 4304
rect 6063 4270 6097 4304
rect 6255 4270 6289 4304
rect 6482 4277 6516 4311
rect 4610 3490 4650 3580
rect 4650 3490 4660 3580
rect 4738 3713 4772 4201
rect 4826 3713 4860 4201
rect 4982 3877 5016 3911
rect 4938 3242 4972 3818
rect 5026 3242 5060 3818
rect 5151 3706 5185 4194
rect 5247 3252 5281 3740
rect 5343 3706 5377 4194
rect 5439 3252 5473 3740
rect 5535 3706 5569 4194
rect 5631 3252 5665 3740
rect 5727 3706 5761 4194
rect 5823 3252 5857 3740
rect 5919 3706 5953 4194
rect 6015 3252 6049 3740
rect 6111 3706 6145 4194
rect 6207 3252 6241 3740
rect 6303 3706 6337 4194
rect 6438 3242 6472 4218
rect 6526 3242 6560 4218
rect 4782 3149 4816 3183
rect 4982 3149 5016 3183
rect 5199 3142 5233 3176
rect 5391 3142 5425 3176
rect 5583 3142 5617 3176
rect 5775 3142 5809 3176
rect 5967 3142 6001 3176
rect 6159 3142 6193 3176
rect 6482 3149 6516 3183
rect 8082 4277 8116 4311
rect 8595 4270 8629 4304
rect 8787 4270 8821 4304
rect 8979 4270 9013 4304
rect 9171 4270 9205 4304
rect 9363 4270 9397 4304
rect 9555 4270 9589 4304
rect 9782 4277 9816 4311
rect 7910 3490 7950 3580
rect 7950 3490 7960 3580
rect 8038 3713 8072 4201
rect 8126 3713 8160 4201
rect 8282 3877 8316 3911
rect 8238 3242 8272 3818
rect 8326 3242 8360 3818
rect 8451 3706 8485 4194
rect 8547 3252 8581 3740
rect 8643 3706 8677 4194
rect 8739 3252 8773 3740
rect 8835 3706 8869 4194
rect 8931 3252 8965 3740
rect 9027 3706 9061 4194
rect 9123 3252 9157 3740
rect 9219 3706 9253 4194
rect 9315 3252 9349 3740
rect 9411 3706 9445 4194
rect 9507 3252 9541 3740
rect 9603 3706 9637 4194
rect 9738 3242 9772 4218
rect 9826 3242 9860 4218
rect 8082 3149 8116 3183
rect 8282 3149 8316 3183
rect 8499 3142 8533 3176
rect 8691 3142 8725 3176
rect 8883 3142 8917 3176
rect 9075 3142 9109 3176
rect 9267 3142 9301 3176
rect 9459 3142 9493 3176
rect 9782 3149 9816 3183
rect 11382 4277 11416 4311
rect 11895 4270 11929 4304
rect 12087 4270 12121 4304
rect 12279 4270 12313 4304
rect 12471 4270 12505 4304
rect 12663 4270 12697 4304
rect 12855 4270 12889 4304
rect 13082 4277 13116 4311
rect 11210 3490 11250 3580
rect 11250 3490 11260 3580
rect 11338 3713 11372 4201
rect 11426 3713 11460 4201
rect 11582 3877 11616 3911
rect 11538 3242 11572 3818
rect 11626 3242 11660 3818
rect 11751 3706 11785 4194
rect 11847 3252 11881 3740
rect 11943 3706 11977 4194
rect 12039 3252 12073 3740
rect 12135 3706 12169 4194
rect 12231 3252 12265 3740
rect 12327 3706 12361 4194
rect 12423 3252 12457 3740
rect 12519 3706 12553 4194
rect 12615 3252 12649 3740
rect 12711 3706 12745 4194
rect 12807 3252 12841 3740
rect 12903 3706 12937 4194
rect 13038 3242 13072 4218
rect 13126 3242 13160 4218
rect 11382 3149 11416 3183
rect 11582 3149 11616 3183
rect 11799 3142 11833 3176
rect 11991 3142 12025 3176
rect 12183 3142 12217 3176
rect 12375 3142 12409 3176
rect 12567 3142 12601 3176
rect 12759 3142 12793 3176
rect 13082 3149 13116 3183
rect 14982 4277 15016 4311
rect 15495 4270 15529 4304
rect 15687 4270 15721 4304
rect 15879 4270 15913 4304
rect 16071 4270 16105 4304
rect 16263 4270 16297 4304
rect 16455 4270 16489 4304
rect 16682 4277 16716 4311
rect 14810 3490 14850 3580
rect 14850 3490 14860 3580
rect 14938 3713 14972 4201
rect 15026 3713 15060 4201
rect 15182 3877 15216 3911
rect 15138 3242 15172 3818
rect 15226 3242 15260 3818
rect 15351 3706 15385 4194
rect 15447 3252 15481 3740
rect 15543 3706 15577 4194
rect 15639 3252 15673 3740
rect 15735 3706 15769 4194
rect 15831 3252 15865 3740
rect 15927 3706 15961 4194
rect 16023 3252 16057 3740
rect 16119 3706 16153 4194
rect 16215 3252 16249 3740
rect 16311 3706 16345 4194
rect 16407 3252 16441 3740
rect 16503 3706 16537 4194
rect 16638 3242 16672 4218
rect 16726 3242 16760 4218
rect 14982 3149 15016 3183
rect 15182 3149 15216 3183
rect 15399 3142 15433 3176
rect 15591 3142 15625 3176
rect 15783 3142 15817 3176
rect 15975 3142 16009 3176
rect 16167 3142 16201 3176
rect 16359 3142 16393 3176
rect 16682 3149 16716 3183
rect 18482 4277 18516 4311
rect 18995 4270 19029 4304
rect 19187 4270 19221 4304
rect 19379 4270 19413 4304
rect 19571 4270 19605 4304
rect 19763 4270 19797 4304
rect 19955 4270 19989 4304
rect 20182 4277 20216 4311
rect 18310 3490 18350 3580
rect 18350 3490 18360 3580
rect 18438 3713 18472 4201
rect 18526 3713 18560 4201
rect 18682 3877 18716 3911
rect 18638 3242 18672 3818
rect 18726 3242 18760 3818
rect 18851 3706 18885 4194
rect 18947 3252 18981 3740
rect 19043 3706 19077 4194
rect 19139 3252 19173 3740
rect 19235 3706 19269 4194
rect 19331 3252 19365 3740
rect 19427 3706 19461 4194
rect 19523 3252 19557 3740
rect 19619 3706 19653 4194
rect 19715 3252 19749 3740
rect 19811 3706 19845 4194
rect 19907 3252 19941 3740
rect 20003 3706 20037 4194
rect 20138 3242 20172 4218
rect 20226 3242 20260 4218
rect 18482 3149 18516 3183
rect 18682 3149 18716 3183
rect 18899 3142 18933 3176
rect 19091 3142 19125 3176
rect 19283 3142 19317 3176
rect 19475 3142 19509 3176
rect 19667 3142 19701 3176
rect 19859 3142 19893 3176
rect 20182 3149 20216 3183
rect 22182 4277 22216 4311
rect 22695 4270 22729 4304
rect 22887 4270 22921 4304
rect 23079 4270 23113 4304
rect 23271 4270 23305 4304
rect 23463 4270 23497 4304
rect 23655 4270 23689 4304
rect 23882 4277 23916 4311
rect 22010 3490 22050 3580
rect 22050 3490 22060 3580
rect 22138 3713 22172 4201
rect 22226 3713 22260 4201
rect 22382 3877 22416 3911
rect 22338 3242 22372 3818
rect 22426 3242 22460 3818
rect 22551 3706 22585 4194
rect 22647 3252 22681 3740
rect 22743 3706 22777 4194
rect 22839 3252 22873 3740
rect 22935 3706 22969 4194
rect 23031 3252 23065 3740
rect 23127 3706 23161 4194
rect 23223 3252 23257 3740
rect 23319 3706 23353 4194
rect 23415 3252 23449 3740
rect 23511 3706 23545 4194
rect 23607 3252 23641 3740
rect 23703 3706 23737 4194
rect 23838 3242 23872 4218
rect 23926 3242 23960 4218
rect 22182 3149 22216 3183
rect 22382 3149 22416 3183
rect 22599 3142 22633 3176
rect 22791 3142 22825 3176
rect 22983 3142 23017 3176
rect 23175 3142 23209 3176
rect 23367 3142 23401 3176
rect 23559 3142 23593 3176
rect 23882 3149 23916 3183
rect 25982 4277 26016 4311
rect 26495 4270 26529 4304
rect 26687 4270 26721 4304
rect 26879 4270 26913 4304
rect 27071 4270 27105 4304
rect 27263 4270 27297 4304
rect 27455 4270 27489 4304
rect 27682 4277 27716 4311
rect 25810 3490 25850 3580
rect 25850 3490 25860 3580
rect 25938 3713 25972 4201
rect 26026 3713 26060 4201
rect 26182 3877 26216 3911
rect 26138 3242 26172 3818
rect 26226 3242 26260 3818
rect 26351 3706 26385 4194
rect 26447 3252 26481 3740
rect 26543 3706 26577 4194
rect 26639 3252 26673 3740
rect 26735 3706 26769 4194
rect 26831 3252 26865 3740
rect 26927 3706 26961 4194
rect 27023 3252 27057 3740
rect 27119 3706 27153 4194
rect 27215 3252 27249 3740
rect 27311 3706 27345 4194
rect 27407 3252 27441 3740
rect 27503 3706 27537 4194
rect 27638 3242 27672 4218
rect 27726 3242 27760 4218
rect 25982 3149 26016 3183
rect 26182 3149 26216 3183
rect 26399 3142 26433 3176
rect 26591 3142 26625 3176
rect 26783 3142 26817 3176
rect 26975 3142 27009 3176
rect 27167 3142 27201 3176
rect 27359 3142 27393 3176
rect 27682 3149 27716 3183
rect 29934 4596 30102 4630
rect 30314 4596 30482 4630
rect 30714 4596 30882 4630
rect 31094 4596 31262 4630
rect 31352 4596 31520 4630
rect 31610 4596 31778 4630
rect 31868 4596 32036 4630
rect 32126 4596 32294 4630
rect 32384 4596 32552 4630
rect 32642 4596 32810 4630
rect 32900 4596 33068 4630
rect 33158 4596 33326 4630
rect 33534 4596 33702 4630
rect 29872 4370 29906 4546
rect 30130 4370 30164 4546
rect 30252 4370 30286 4546
rect 30510 4370 30544 4546
rect 30652 4370 30686 4546
rect 30910 4370 30944 4546
rect 31032 4441 31066 4529
rect 31290 4387 31324 4475
rect 31548 4441 31582 4529
rect 31806 4387 31840 4475
rect 32064 4441 32098 4529
rect 32322 4387 32356 4475
rect 32580 4441 32614 4529
rect 32838 4387 32872 4475
rect 33096 4441 33130 4529
rect 33354 4387 33388 4475
rect 33472 4370 33506 4546
rect 33730 4370 33764 4546
rect 29934 4286 30102 4320
rect 30314 4286 30482 4320
rect 30714 4286 30882 4320
rect 31094 4286 31262 4320
rect 31352 4286 31520 4320
rect 31610 4286 31778 4320
rect 31868 4286 32036 4320
rect 32126 4286 32294 4320
rect 32384 4286 32552 4320
rect 32642 4286 32810 4320
rect 32900 4286 33068 4320
rect 33158 4286 33326 4320
rect 33534 4286 33702 4320
rect 29900 4050 30160 4090
rect 440 2510 620 2690
rect 1486 2746 1520 2780
rect 1686 2746 1720 2780
rect 1999 2739 2033 2773
rect 2191 2739 2225 2773
rect 2383 2739 2417 2773
rect 2575 2739 2609 2773
rect 2767 2739 2801 2773
rect 2959 2739 2993 2773
rect 3166 2746 3200 2780
rect 1300 2540 1310 2670
rect 1310 2540 1350 2670
rect 1350 2540 1360 2670
rect 1442 2191 1476 2679
rect 1530 2191 1564 2679
rect 1642 2520 1676 2696
rect 1730 2520 1764 2696
rect 1686 2436 1720 2470
rect 1855 2184 1889 2672
rect 1951 1730 1985 2218
rect 2047 2184 2081 2672
rect 2143 1730 2177 2218
rect 2239 2184 2273 2672
rect 2335 1730 2369 2218
rect 2431 2184 2465 2672
rect 2527 1730 2561 2218
rect 2623 2184 2657 2672
rect 2719 1730 2753 2218
rect 2815 2184 2849 2672
rect 2911 1730 2945 2218
rect 3007 2184 3041 2672
rect 3122 1737 3156 2225
rect 3210 1737 3244 2225
rect 1486 1636 1520 1670
rect 1903 1629 1937 1663
rect 2095 1629 2129 1663
rect 2287 1629 2321 1663
rect 2479 1629 2513 1663
rect 2671 1629 2705 1663
rect 2863 1629 2897 1663
rect 3166 1636 3200 1670
rect 4786 2746 4820 2780
rect 4986 2746 5020 2780
rect 5299 2739 5333 2773
rect 5491 2739 5525 2773
rect 5683 2739 5717 2773
rect 5875 2739 5909 2773
rect 6067 2739 6101 2773
rect 6259 2739 6293 2773
rect 6466 2746 6500 2780
rect 4600 2540 4610 2670
rect 4610 2540 4650 2670
rect 4650 2540 4660 2670
rect 4742 2191 4776 2679
rect 4830 2191 4864 2679
rect 4942 2520 4976 2696
rect 5030 2520 5064 2696
rect 4986 2436 5020 2470
rect 5155 2184 5189 2672
rect 5251 1730 5285 2218
rect 5347 2184 5381 2672
rect 5443 1730 5477 2218
rect 5539 2184 5573 2672
rect 5635 1730 5669 2218
rect 5731 2184 5765 2672
rect 5827 1730 5861 2218
rect 5923 2184 5957 2672
rect 6019 1730 6053 2218
rect 6115 2184 6149 2672
rect 6211 1730 6245 2218
rect 6307 2184 6341 2672
rect 6422 1737 6456 2225
rect 6510 1737 6544 2225
rect 4786 1636 4820 1670
rect 5203 1629 5237 1663
rect 5395 1629 5429 1663
rect 5587 1629 5621 1663
rect 5779 1629 5813 1663
rect 5971 1629 6005 1663
rect 6163 1629 6197 1663
rect 6466 1636 6500 1670
rect 8086 2746 8120 2780
rect 8286 2746 8320 2780
rect 8599 2739 8633 2773
rect 8791 2739 8825 2773
rect 8983 2739 9017 2773
rect 9175 2739 9209 2773
rect 9367 2739 9401 2773
rect 9559 2739 9593 2773
rect 9766 2746 9800 2780
rect 7900 2540 7910 2670
rect 7910 2540 7950 2670
rect 7950 2540 7960 2670
rect 8042 2191 8076 2679
rect 8130 2191 8164 2679
rect 8242 2520 8276 2696
rect 8330 2520 8364 2696
rect 8286 2436 8320 2470
rect 8455 2184 8489 2672
rect 8551 1730 8585 2218
rect 8647 2184 8681 2672
rect 8743 1730 8777 2218
rect 8839 2184 8873 2672
rect 8935 1730 8969 2218
rect 9031 2184 9065 2672
rect 9127 1730 9161 2218
rect 9223 2184 9257 2672
rect 9319 1730 9353 2218
rect 9415 2184 9449 2672
rect 9511 1730 9545 2218
rect 9607 2184 9641 2672
rect 9722 1737 9756 2225
rect 9810 1737 9844 2225
rect 8086 1636 8120 1670
rect 8503 1629 8537 1663
rect 8695 1629 8729 1663
rect 8887 1629 8921 1663
rect 9079 1629 9113 1663
rect 9271 1629 9305 1663
rect 9463 1629 9497 1663
rect 9766 1636 9800 1670
rect 11386 2746 11420 2780
rect 11586 2746 11620 2780
rect 11899 2739 11933 2773
rect 12091 2739 12125 2773
rect 12283 2739 12317 2773
rect 12475 2739 12509 2773
rect 12667 2739 12701 2773
rect 12859 2739 12893 2773
rect 13066 2746 13100 2780
rect 11200 2540 11210 2670
rect 11210 2540 11250 2670
rect 11250 2540 11260 2670
rect 11342 2191 11376 2679
rect 11430 2191 11464 2679
rect 11542 2520 11576 2696
rect 11630 2520 11664 2696
rect 11586 2436 11620 2470
rect 11755 2184 11789 2672
rect 11851 1730 11885 2218
rect 11947 2184 11981 2672
rect 12043 1730 12077 2218
rect 12139 2184 12173 2672
rect 12235 1730 12269 2218
rect 12331 2184 12365 2672
rect 12427 1730 12461 2218
rect 12523 2184 12557 2672
rect 12619 1730 12653 2218
rect 12715 2184 12749 2672
rect 12811 1730 12845 2218
rect 12907 2184 12941 2672
rect 13022 1737 13056 2225
rect 13110 1737 13144 2225
rect 11386 1636 11420 1670
rect 11803 1629 11837 1663
rect 11995 1629 12029 1663
rect 12187 1629 12221 1663
rect 12379 1629 12413 1663
rect 12571 1629 12605 1663
rect 12763 1629 12797 1663
rect 13066 1636 13100 1670
rect 14986 2746 15020 2780
rect 15186 2746 15220 2780
rect 15499 2739 15533 2773
rect 15691 2739 15725 2773
rect 15883 2739 15917 2773
rect 16075 2739 16109 2773
rect 16267 2739 16301 2773
rect 16459 2739 16493 2773
rect 16666 2746 16700 2780
rect 14800 2540 14810 2670
rect 14810 2540 14850 2670
rect 14850 2540 14860 2670
rect 14942 2191 14976 2679
rect 15030 2191 15064 2679
rect 15142 2520 15176 2696
rect 15230 2520 15264 2696
rect 15186 2436 15220 2470
rect 15355 2184 15389 2672
rect 15451 1730 15485 2218
rect 15547 2184 15581 2672
rect 15643 1730 15677 2218
rect 15739 2184 15773 2672
rect 15835 1730 15869 2218
rect 15931 2184 15965 2672
rect 16027 1730 16061 2218
rect 16123 2184 16157 2672
rect 16219 1730 16253 2218
rect 16315 2184 16349 2672
rect 16411 1730 16445 2218
rect 16507 2184 16541 2672
rect 16622 1737 16656 2225
rect 16710 1737 16744 2225
rect 14986 1636 15020 1670
rect 15403 1629 15437 1663
rect 15595 1629 15629 1663
rect 15787 1629 15821 1663
rect 15979 1629 16013 1663
rect 16171 1629 16205 1663
rect 16363 1629 16397 1663
rect 16666 1636 16700 1670
rect 18486 2746 18520 2780
rect 18686 2746 18720 2780
rect 18999 2739 19033 2773
rect 19191 2739 19225 2773
rect 19383 2739 19417 2773
rect 19575 2739 19609 2773
rect 19767 2739 19801 2773
rect 19959 2739 19993 2773
rect 20166 2746 20200 2780
rect 18300 2540 18310 2670
rect 18310 2540 18350 2670
rect 18350 2540 18360 2670
rect 18442 2191 18476 2679
rect 18530 2191 18564 2679
rect 18642 2520 18676 2696
rect 18730 2520 18764 2696
rect 18686 2436 18720 2470
rect 18855 2184 18889 2672
rect 18951 1730 18985 2218
rect 19047 2184 19081 2672
rect 19143 1730 19177 2218
rect 19239 2184 19273 2672
rect 19335 1730 19369 2218
rect 19431 2184 19465 2672
rect 19527 1730 19561 2218
rect 19623 2184 19657 2672
rect 19719 1730 19753 2218
rect 19815 2184 19849 2672
rect 19911 1730 19945 2218
rect 20007 2184 20041 2672
rect 20122 1737 20156 2225
rect 20210 1737 20244 2225
rect 18486 1636 18520 1670
rect 18903 1629 18937 1663
rect 19095 1629 19129 1663
rect 19287 1629 19321 1663
rect 19479 1629 19513 1663
rect 19671 1629 19705 1663
rect 19863 1629 19897 1663
rect 20166 1636 20200 1670
rect 22186 2746 22220 2780
rect 22386 2746 22420 2780
rect 22699 2739 22733 2773
rect 22891 2739 22925 2773
rect 23083 2739 23117 2773
rect 23275 2739 23309 2773
rect 23467 2739 23501 2773
rect 23659 2739 23693 2773
rect 23866 2746 23900 2780
rect 22000 2540 22010 2670
rect 22010 2540 22050 2670
rect 22050 2540 22060 2670
rect 22142 2191 22176 2679
rect 22230 2191 22264 2679
rect 22342 2520 22376 2696
rect 22430 2520 22464 2696
rect 22386 2436 22420 2470
rect 22555 2184 22589 2672
rect 22651 1730 22685 2218
rect 22747 2184 22781 2672
rect 22843 1730 22877 2218
rect 22939 2184 22973 2672
rect 23035 1730 23069 2218
rect 23131 2184 23165 2672
rect 23227 1730 23261 2218
rect 23323 2184 23357 2672
rect 23419 1730 23453 2218
rect 23515 2184 23549 2672
rect 23611 1730 23645 2218
rect 23707 2184 23741 2672
rect 23822 1737 23856 2225
rect 23910 1737 23944 2225
rect 22186 1636 22220 1670
rect 22603 1629 22637 1663
rect 22795 1629 22829 1663
rect 22987 1629 23021 1663
rect 23179 1629 23213 1663
rect 23371 1629 23405 1663
rect 23563 1629 23597 1663
rect 23866 1636 23900 1670
rect 25986 2746 26020 2780
rect 26186 2746 26220 2780
rect 26499 2739 26533 2773
rect 26691 2739 26725 2773
rect 26883 2739 26917 2773
rect 27075 2739 27109 2773
rect 27267 2739 27301 2773
rect 27459 2739 27493 2773
rect 27666 2746 27700 2780
rect 25800 2540 25810 2670
rect 25810 2540 25850 2670
rect 25850 2540 25860 2670
rect 25942 2191 25976 2679
rect 26030 2191 26064 2679
rect 26142 2520 26176 2696
rect 26230 2520 26264 2696
rect 26186 2436 26220 2470
rect 26355 2184 26389 2672
rect 26451 1730 26485 2218
rect 26547 2184 26581 2672
rect 26643 1730 26677 2218
rect 26739 2184 26773 2672
rect 26835 1730 26869 2218
rect 26931 2184 26965 2672
rect 27027 1730 27061 2218
rect 27123 2184 27157 2672
rect 27219 1730 27253 2218
rect 27315 2184 27349 2672
rect 27411 1730 27445 2218
rect 27507 2184 27541 2672
rect 27622 1737 27656 2225
rect 27710 1737 27744 2225
rect 25986 1636 26020 1670
rect 26403 1629 26437 1663
rect 26595 1629 26629 1663
rect 26787 1629 26821 1663
rect 26979 1629 27013 1663
rect 27171 1629 27205 1663
rect 27363 1629 27397 1663
rect 27666 1636 27700 1670
<< metal1 >>
rect 4948 27434 20220 27456
rect 4948 27425 6043 27434
rect 6095 27425 6107 27434
rect 4948 27391 4977 27425
rect 5011 27391 5069 27425
rect 5103 27391 5161 27425
rect 5195 27391 5253 27425
rect 5287 27391 5345 27425
rect 5379 27391 5437 27425
rect 5471 27391 5529 27425
rect 5563 27391 5621 27425
rect 5655 27391 5713 27425
rect 5747 27391 5805 27425
rect 5839 27391 5897 27425
rect 5931 27391 5989 27425
rect 6023 27391 6043 27425
rect 4948 27382 6043 27391
rect 6095 27382 6107 27391
rect 6159 27382 6171 27434
rect 6223 27382 6235 27434
rect 6287 27425 6299 27434
rect 6287 27382 6299 27391
rect 6351 27425 9861 27434
rect 6351 27391 6357 27425
rect 6391 27391 6449 27425
rect 6483 27391 6541 27425
rect 6575 27391 6633 27425
rect 6667 27391 6725 27425
rect 6759 27391 6817 27425
rect 6851 27391 6909 27425
rect 6943 27391 7001 27425
rect 7035 27391 7093 27425
rect 7127 27391 7185 27425
rect 7219 27391 7277 27425
rect 7311 27391 7369 27425
rect 7403 27391 7461 27425
rect 7495 27391 7553 27425
rect 7587 27391 7645 27425
rect 7679 27391 7737 27425
rect 7771 27391 7829 27425
rect 7863 27391 7921 27425
rect 7955 27391 8013 27425
rect 8047 27391 8105 27425
rect 8139 27391 8197 27425
rect 8231 27391 8289 27425
rect 8323 27391 8381 27425
rect 8415 27391 8473 27425
rect 8507 27391 8565 27425
rect 8599 27391 8657 27425
rect 8691 27391 8749 27425
rect 8783 27391 8841 27425
rect 8875 27391 8933 27425
rect 8967 27391 9025 27425
rect 9059 27391 9117 27425
rect 9151 27391 9209 27425
rect 9243 27391 9301 27425
rect 9335 27391 9393 27425
rect 9427 27391 9485 27425
rect 9519 27391 9577 27425
rect 9611 27391 9669 27425
rect 9703 27391 9761 27425
rect 9795 27391 9853 27425
rect 6351 27382 9861 27391
rect 9913 27382 9925 27434
rect 9977 27425 9989 27434
rect 10041 27425 10053 27434
rect 9979 27391 9989 27425
rect 9977 27382 9989 27391
rect 10041 27382 10053 27391
rect 10105 27382 10117 27434
rect 10169 27425 13679 27434
rect 13731 27425 13743 27434
rect 10169 27391 10221 27425
rect 10255 27391 10313 27425
rect 10347 27391 10405 27425
rect 10439 27391 10497 27425
rect 10531 27391 10589 27425
rect 10623 27391 10681 27425
rect 10715 27391 10773 27425
rect 10807 27391 10865 27425
rect 10899 27391 10957 27425
rect 10991 27391 11049 27425
rect 11083 27391 11141 27425
rect 11175 27391 11233 27425
rect 11267 27391 11325 27425
rect 11359 27391 11417 27425
rect 11451 27391 11509 27425
rect 11543 27391 11601 27425
rect 11635 27391 11693 27425
rect 11727 27391 11785 27425
rect 11819 27391 11877 27425
rect 11911 27391 11969 27425
rect 12003 27391 12061 27425
rect 12095 27391 12153 27425
rect 12187 27391 12245 27425
rect 12279 27391 12337 27425
rect 12371 27391 12429 27425
rect 12463 27391 12521 27425
rect 12555 27391 12613 27425
rect 12647 27391 12705 27425
rect 12739 27391 12797 27425
rect 12831 27391 12889 27425
rect 12923 27391 12981 27425
rect 13015 27391 13073 27425
rect 13107 27391 13165 27425
rect 13199 27391 13257 27425
rect 13291 27391 13349 27425
rect 13383 27391 13441 27425
rect 13475 27391 13533 27425
rect 13567 27391 13625 27425
rect 13659 27391 13679 27425
rect 10169 27382 13679 27391
rect 13731 27382 13743 27391
rect 13795 27382 13807 27434
rect 13859 27382 13871 27434
rect 13923 27425 13935 27434
rect 13923 27382 13935 27391
rect 13987 27425 17497 27434
rect 13987 27391 13993 27425
rect 14027 27391 14085 27425
rect 14119 27391 14177 27425
rect 14211 27391 14269 27425
rect 14303 27391 14361 27425
rect 14395 27391 14453 27425
rect 14487 27391 14545 27425
rect 14579 27391 14637 27425
rect 14671 27391 14729 27425
rect 14763 27391 14821 27425
rect 14855 27391 14913 27425
rect 14947 27391 15005 27425
rect 15039 27391 15097 27425
rect 15131 27391 15189 27425
rect 15223 27391 15281 27425
rect 15315 27391 15373 27425
rect 15407 27391 15465 27425
rect 15499 27391 15557 27425
rect 15591 27391 15649 27425
rect 15683 27391 15741 27425
rect 15775 27391 15833 27425
rect 15867 27391 15925 27425
rect 15959 27391 16017 27425
rect 16051 27391 16109 27425
rect 16143 27391 16201 27425
rect 16235 27391 16293 27425
rect 16327 27391 16385 27425
rect 16419 27391 16477 27425
rect 16511 27391 16569 27425
rect 16603 27391 16661 27425
rect 16695 27391 16753 27425
rect 16787 27391 16845 27425
rect 16879 27391 16937 27425
rect 16971 27391 17029 27425
rect 17063 27391 17121 27425
rect 17155 27391 17213 27425
rect 17247 27391 17305 27425
rect 17339 27391 17397 27425
rect 17431 27391 17489 27425
rect 13987 27382 17497 27391
rect 17549 27382 17561 27434
rect 17613 27425 17625 27434
rect 17677 27425 17689 27434
rect 17615 27391 17625 27425
rect 17613 27382 17625 27391
rect 17677 27382 17689 27391
rect 17741 27382 17753 27434
rect 17805 27425 20220 27434
rect 17805 27391 17857 27425
rect 17891 27391 17949 27425
rect 17983 27391 18041 27425
rect 18075 27391 18133 27425
rect 18167 27391 18225 27425
rect 18259 27391 18317 27425
rect 18351 27391 18409 27425
rect 18443 27391 18501 27425
rect 18535 27391 18593 27425
rect 18627 27391 18685 27425
rect 18719 27391 18777 27425
rect 18811 27391 18869 27425
rect 18903 27391 18961 27425
rect 18995 27391 19053 27425
rect 19087 27391 19145 27425
rect 19179 27391 19237 27425
rect 19271 27391 19329 27425
rect 19363 27391 19421 27425
rect 19455 27391 19513 27425
rect 19547 27391 19605 27425
rect 19639 27391 19697 27425
rect 19731 27391 19789 27425
rect 19823 27391 19881 27425
rect 19915 27391 19973 27425
rect 20007 27391 20065 27425
rect 20099 27391 20157 27425
rect 20191 27391 20220 27425
rect 17805 27382 20220 27391
rect 4948 27360 20220 27382
rect 10206 27280 10212 27332
rect 10264 27280 10270 27332
rect 5882 27212 5888 27264
rect 5940 27212 5946 27264
rect 10117 27187 10175 27193
rect 10117 27153 10129 27187
rect 10163 27184 10175 27187
rect 10224 27184 10252 27280
rect 18857 27255 18915 27261
rect 18857 27221 18869 27255
rect 18903 27252 18915 27255
rect 19038 27252 19044 27264
rect 18903 27224 19044 27252
rect 18903 27221 18915 27224
rect 18857 27215 18915 27221
rect 19038 27212 19044 27224
rect 19096 27212 19102 27264
rect 10163 27156 10252 27184
rect 10163 27153 10175 27156
rect 10117 27147 10175 27153
rect 5790 26940 5796 26992
rect 5848 26940 5854 26992
rect 10301 26983 10359 26989
rect 10301 26949 10313 26983
rect 10347 26980 10359 26983
rect 11034 26980 11040 26992
rect 10347 26952 11040 26980
rect 10347 26949 10359 26952
rect 10301 26943 10359 26949
rect 11034 26940 11040 26952
rect 11092 26940 11098 26992
rect 18762 26940 18768 26992
rect 18820 26940 18826 26992
rect 4948 26890 20220 26912
rect 4948 26881 6703 26890
rect 6755 26881 6767 26890
rect 6819 26881 6831 26890
rect 4948 26847 4977 26881
rect 5011 26847 5069 26881
rect 5103 26847 5161 26881
rect 5195 26847 5253 26881
rect 5287 26847 5345 26881
rect 5379 26847 5437 26881
rect 5471 26847 5529 26881
rect 5563 26847 5621 26881
rect 5655 26847 5713 26881
rect 5747 26847 5805 26881
rect 5839 26847 5897 26881
rect 5931 26847 5989 26881
rect 6023 26847 6081 26881
rect 6115 26847 6173 26881
rect 6207 26847 6265 26881
rect 6299 26847 6357 26881
rect 6391 26847 6449 26881
rect 6483 26847 6541 26881
rect 6575 26847 6633 26881
rect 6667 26847 6703 26881
rect 6759 26847 6767 26881
rect 4948 26838 6703 26847
rect 6755 26838 6767 26847
rect 6819 26838 6831 26847
rect 6883 26838 6895 26890
rect 6947 26838 6959 26890
rect 7011 26881 10521 26890
rect 7035 26847 7093 26881
rect 7127 26847 7185 26881
rect 7219 26847 7277 26881
rect 7311 26847 7369 26881
rect 7403 26847 7461 26881
rect 7495 26847 7553 26881
rect 7587 26847 7645 26881
rect 7679 26847 7737 26881
rect 7771 26847 7829 26881
rect 7863 26847 7921 26881
rect 7955 26847 8013 26881
rect 8047 26847 8105 26881
rect 8139 26847 8197 26881
rect 8231 26847 8289 26881
rect 8323 26847 8381 26881
rect 8415 26847 8473 26881
rect 8507 26847 8565 26881
rect 8599 26847 8657 26881
rect 8691 26847 8749 26881
rect 8783 26847 8841 26881
rect 8875 26847 8933 26881
rect 8967 26847 9025 26881
rect 9059 26847 9117 26881
rect 9151 26847 9209 26881
rect 9243 26847 9301 26881
rect 9335 26847 9393 26881
rect 9427 26847 9485 26881
rect 9519 26847 9577 26881
rect 9611 26847 9669 26881
rect 9703 26847 9761 26881
rect 9795 26847 9853 26881
rect 9887 26847 9945 26881
rect 9979 26847 10037 26881
rect 10071 26847 10129 26881
rect 10163 26847 10221 26881
rect 10255 26847 10313 26881
rect 10347 26847 10405 26881
rect 10439 26847 10497 26881
rect 7011 26838 10521 26847
rect 10573 26838 10585 26890
rect 10637 26838 10649 26890
rect 10701 26881 10713 26890
rect 10765 26881 10777 26890
rect 10829 26881 14339 26890
rect 14391 26881 14403 26890
rect 14455 26881 14467 26890
rect 10765 26847 10773 26881
rect 10829 26847 10865 26881
rect 10899 26847 10957 26881
rect 10991 26847 11049 26881
rect 11083 26847 11141 26881
rect 11175 26847 11233 26881
rect 11267 26847 11325 26881
rect 11359 26847 11417 26881
rect 11451 26847 11509 26881
rect 11543 26847 11601 26881
rect 11635 26847 11693 26881
rect 11727 26847 11785 26881
rect 11819 26847 11877 26881
rect 11911 26847 11969 26881
rect 12003 26847 12061 26881
rect 12095 26847 12153 26881
rect 12187 26847 12245 26881
rect 12279 26847 12337 26881
rect 12371 26847 12429 26881
rect 12463 26847 12521 26881
rect 12555 26847 12613 26881
rect 12647 26847 12705 26881
rect 12739 26847 12797 26881
rect 12831 26847 12889 26881
rect 12923 26847 12981 26881
rect 13015 26847 13073 26881
rect 13107 26847 13165 26881
rect 13199 26847 13257 26881
rect 13291 26847 13349 26881
rect 13383 26847 13441 26881
rect 13475 26847 13533 26881
rect 13567 26847 13625 26881
rect 13659 26847 13717 26881
rect 13751 26847 13809 26881
rect 13843 26847 13901 26881
rect 13935 26847 13993 26881
rect 14027 26847 14085 26881
rect 14119 26847 14177 26881
rect 14211 26847 14269 26881
rect 14303 26847 14339 26881
rect 14395 26847 14403 26881
rect 10701 26838 10713 26847
rect 10765 26838 10777 26847
rect 10829 26838 14339 26847
rect 14391 26838 14403 26847
rect 14455 26838 14467 26847
rect 14519 26838 14531 26890
rect 14583 26838 14595 26890
rect 14647 26881 18157 26890
rect 14671 26847 14729 26881
rect 14763 26847 14821 26881
rect 14855 26847 14913 26881
rect 14947 26847 15005 26881
rect 15039 26847 15097 26881
rect 15131 26847 15189 26881
rect 15223 26847 15281 26881
rect 15315 26847 15373 26881
rect 15407 26847 15465 26881
rect 15499 26847 15557 26881
rect 15591 26847 15649 26881
rect 15683 26847 15741 26881
rect 15775 26847 15833 26881
rect 15867 26847 15925 26881
rect 15959 26847 16017 26881
rect 16051 26847 16109 26881
rect 16143 26847 16201 26881
rect 16235 26847 16293 26881
rect 16327 26847 16385 26881
rect 16419 26847 16477 26881
rect 16511 26847 16569 26881
rect 16603 26847 16661 26881
rect 16695 26847 16753 26881
rect 16787 26847 16845 26881
rect 16879 26847 16937 26881
rect 16971 26847 17029 26881
rect 17063 26847 17121 26881
rect 17155 26847 17213 26881
rect 17247 26847 17305 26881
rect 17339 26847 17397 26881
rect 17431 26847 17489 26881
rect 17523 26847 17581 26881
rect 17615 26847 17673 26881
rect 17707 26847 17765 26881
rect 17799 26847 17857 26881
rect 17891 26847 17949 26881
rect 17983 26847 18041 26881
rect 18075 26847 18133 26881
rect 14647 26838 18157 26847
rect 18209 26838 18221 26890
rect 18273 26838 18285 26890
rect 18337 26881 18349 26890
rect 18401 26881 18413 26890
rect 18465 26881 20220 26890
rect 18401 26847 18409 26881
rect 18465 26847 18501 26881
rect 18535 26847 18593 26881
rect 18627 26847 18685 26881
rect 18719 26847 18777 26881
rect 18811 26847 18869 26881
rect 18903 26847 18961 26881
rect 18995 26847 19053 26881
rect 19087 26847 19145 26881
rect 19179 26847 19237 26881
rect 19271 26847 19329 26881
rect 19363 26847 19421 26881
rect 19455 26847 19513 26881
rect 19547 26847 19605 26881
rect 19639 26847 19697 26881
rect 19731 26847 19789 26881
rect 19823 26847 19881 26881
rect 19915 26847 19973 26881
rect 20007 26847 20065 26881
rect 20099 26847 20157 26881
rect 20191 26847 20220 26881
rect 18337 26838 18349 26847
rect 18401 26838 18413 26847
rect 18465 26838 20220 26847
rect 4948 26816 20220 26838
rect 4948 26346 20220 26368
rect 4948 26337 6043 26346
rect 6095 26337 6107 26346
rect 4948 26303 4977 26337
rect 5011 26303 5069 26337
rect 5103 26303 5161 26337
rect 5195 26303 5253 26337
rect 5287 26303 5345 26337
rect 5379 26303 5437 26337
rect 5471 26303 5529 26337
rect 5563 26303 5621 26337
rect 5655 26303 5713 26337
rect 5747 26303 5805 26337
rect 5839 26303 5897 26337
rect 5931 26303 5989 26337
rect 6023 26303 6043 26337
rect 4948 26294 6043 26303
rect 6095 26294 6107 26303
rect 6159 26294 6171 26346
rect 6223 26294 6235 26346
rect 6287 26337 6299 26346
rect 6287 26294 6299 26303
rect 6351 26337 9861 26346
rect 6351 26303 6357 26337
rect 6391 26303 6449 26337
rect 6483 26303 6541 26337
rect 6575 26303 6633 26337
rect 6667 26303 6725 26337
rect 6759 26303 6817 26337
rect 6851 26303 6909 26337
rect 6943 26303 7001 26337
rect 7035 26303 7093 26337
rect 7127 26303 7185 26337
rect 7219 26303 7277 26337
rect 7311 26303 7369 26337
rect 7403 26303 7461 26337
rect 7495 26303 7553 26337
rect 7587 26303 7645 26337
rect 7679 26303 7737 26337
rect 7771 26303 7829 26337
rect 7863 26303 7921 26337
rect 7955 26303 8013 26337
rect 8047 26303 8105 26337
rect 8139 26303 8197 26337
rect 8231 26303 8289 26337
rect 8323 26303 8381 26337
rect 8415 26303 8473 26337
rect 8507 26303 8565 26337
rect 8599 26303 8657 26337
rect 8691 26303 8749 26337
rect 8783 26303 8841 26337
rect 8875 26303 8933 26337
rect 8967 26303 9025 26337
rect 9059 26303 9117 26337
rect 9151 26303 9209 26337
rect 9243 26303 9301 26337
rect 9335 26303 9393 26337
rect 9427 26303 9485 26337
rect 9519 26303 9577 26337
rect 9611 26303 9669 26337
rect 9703 26303 9761 26337
rect 9795 26303 9853 26337
rect 6351 26294 9861 26303
rect 9913 26294 9925 26346
rect 9977 26337 9989 26346
rect 10041 26337 10053 26346
rect 9979 26303 9989 26337
rect 9977 26294 9989 26303
rect 10041 26294 10053 26303
rect 10105 26294 10117 26346
rect 10169 26337 13679 26346
rect 13731 26337 13743 26346
rect 10169 26303 10221 26337
rect 10255 26303 10313 26337
rect 10347 26303 10405 26337
rect 10439 26303 10497 26337
rect 10531 26303 10589 26337
rect 10623 26303 10681 26337
rect 10715 26303 10773 26337
rect 10807 26303 10865 26337
rect 10899 26303 10957 26337
rect 10991 26303 11049 26337
rect 11083 26303 11141 26337
rect 11175 26303 11233 26337
rect 11267 26303 11325 26337
rect 11359 26303 11417 26337
rect 11451 26303 11509 26337
rect 11543 26303 11601 26337
rect 11635 26303 11693 26337
rect 11727 26303 11785 26337
rect 11819 26303 11877 26337
rect 11911 26303 11969 26337
rect 12003 26303 12061 26337
rect 12095 26303 12153 26337
rect 12187 26303 12245 26337
rect 12279 26303 12337 26337
rect 12371 26303 12429 26337
rect 12463 26303 12521 26337
rect 12555 26303 12613 26337
rect 12647 26303 12705 26337
rect 12739 26303 12797 26337
rect 12831 26303 12889 26337
rect 12923 26303 12981 26337
rect 13015 26303 13073 26337
rect 13107 26303 13165 26337
rect 13199 26303 13257 26337
rect 13291 26303 13349 26337
rect 13383 26303 13441 26337
rect 13475 26303 13533 26337
rect 13567 26303 13625 26337
rect 13659 26303 13679 26337
rect 10169 26294 13679 26303
rect 13731 26294 13743 26303
rect 13795 26294 13807 26346
rect 13859 26294 13871 26346
rect 13923 26337 13935 26346
rect 13923 26294 13935 26303
rect 13987 26337 17497 26346
rect 13987 26303 13993 26337
rect 14027 26303 14085 26337
rect 14119 26303 14177 26337
rect 14211 26303 14269 26337
rect 14303 26303 14361 26337
rect 14395 26303 14453 26337
rect 14487 26303 14545 26337
rect 14579 26303 14637 26337
rect 14671 26303 14729 26337
rect 14763 26303 14821 26337
rect 14855 26303 14913 26337
rect 14947 26303 15005 26337
rect 15039 26303 15097 26337
rect 15131 26303 15189 26337
rect 15223 26303 15281 26337
rect 15315 26303 15373 26337
rect 15407 26303 15465 26337
rect 15499 26303 15557 26337
rect 15591 26303 15649 26337
rect 15683 26303 15741 26337
rect 15775 26303 15833 26337
rect 15867 26303 15925 26337
rect 15959 26303 16017 26337
rect 16051 26303 16109 26337
rect 16143 26303 16201 26337
rect 16235 26303 16293 26337
rect 16327 26303 16385 26337
rect 16419 26303 16477 26337
rect 16511 26303 16569 26337
rect 16603 26303 16661 26337
rect 16695 26303 16753 26337
rect 16787 26303 16845 26337
rect 16879 26303 16937 26337
rect 16971 26303 17029 26337
rect 17063 26303 17121 26337
rect 17155 26303 17213 26337
rect 17247 26303 17305 26337
rect 17339 26303 17397 26337
rect 17431 26303 17489 26337
rect 13987 26294 17497 26303
rect 17549 26294 17561 26346
rect 17613 26337 17625 26346
rect 17677 26337 17689 26346
rect 17615 26303 17625 26337
rect 17613 26294 17625 26303
rect 17677 26294 17689 26303
rect 17741 26294 17753 26346
rect 17805 26337 20220 26346
rect 17805 26303 17857 26337
rect 17891 26303 17949 26337
rect 17983 26303 18041 26337
rect 18075 26303 18133 26337
rect 18167 26303 18225 26337
rect 18259 26303 18317 26337
rect 18351 26303 18409 26337
rect 18443 26303 18501 26337
rect 18535 26303 18593 26337
rect 18627 26303 18685 26337
rect 18719 26303 18777 26337
rect 18811 26303 18869 26337
rect 18903 26303 18961 26337
rect 18995 26303 19053 26337
rect 19087 26303 19145 26337
rect 19179 26303 19237 26337
rect 19271 26303 19329 26337
rect 19363 26303 19421 26337
rect 19455 26303 19513 26337
rect 19547 26303 19605 26337
rect 19639 26303 19697 26337
rect 19731 26303 19789 26337
rect 19823 26303 19881 26337
rect 19915 26303 19973 26337
rect 20007 26303 20065 26337
rect 20099 26303 20157 26337
rect 20191 26303 20220 26337
rect 17805 26294 20220 26303
rect 4948 26272 20220 26294
rect 4948 25802 20220 25824
rect 4948 25793 6703 25802
rect 6755 25793 6767 25802
rect 6819 25793 6831 25802
rect 4948 25759 4977 25793
rect 5011 25759 5069 25793
rect 5103 25759 5161 25793
rect 5195 25759 5253 25793
rect 5287 25759 5345 25793
rect 5379 25759 5437 25793
rect 5471 25759 5529 25793
rect 5563 25759 5621 25793
rect 5655 25759 5713 25793
rect 5747 25759 5805 25793
rect 5839 25759 5897 25793
rect 5931 25759 5989 25793
rect 6023 25759 6081 25793
rect 6115 25759 6173 25793
rect 6207 25759 6265 25793
rect 6299 25759 6357 25793
rect 6391 25759 6449 25793
rect 6483 25759 6541 25793
rect 6575 25759 6633 25793
rect 6667 25759 6703 25793
rect 6759 25759 6767 25793
rect 4948 25750 6703 25759
rect 6755 25750 6767 25759
rect 6819 25750 6831 25759
rect 6883 25750 6895 25802
rect 6947 25750 6959 25802
rect 7011 25793 10521 25802
rect 7035 25759 7093 25793
rect 7127 25759 7185 25793
rect 7219 25759 7277 25793
rect 7311 25759 7369 25793
rect 7403 25759 7461 25793
rect 7495 25759 7553 25793
rect 7587 25759 7645 25793
rect 7679 25759 7737 25793
rect 7771 25759 7829 25793
rect 7863 25759 7921 25793
rect 7955 25759 8013 25793
rect 8047 25759 8105 25793
rect 8139 25759 8197 25793
rect 8231 25759 8289 25793
rect 8323 25759 8381 25793
rect 8415 25759 8473 25793
rect 8507 25759 8565 25793
rect 8599 25759 8657 25793
rect 8691 25759 8749 25793
rect 8783 25759 8841 25793
rect 8875 25759 8933 25793
rect 8967 25759 9025 25793
rect 9059 25759 9117 25793
rect 9151 25759 9209 25793
rect 9243 25759 9301 25793
rect 9335 25759 9393 25793
rect 9427 25759 9485 25793
rect 9519 25759 9577 25793
rect 9611 25759 9669 25793
rect 9703 25759 9761 25793
rect 9795 25759 9853 25793
rect 9887 25759 9945 25793
rect 9979 25759 10037 25793
rect 10071 25759 10129 25793
rect 10163 25759 10221 25793
rect 10255 25759 10313 25793
rect 10347 25759 10405 25793
rect 10439 25759 10497 25793
rect 7011 25750 10521 25759
rect 10573 25750 10585 25802
rect 10637 25750 10649 25802
rect 10701 25793 10713 25802
rect 10765 25793 10777 25802
rect 10829 25793 14339 25802
rect 14391 25793 14403 25802
rect 14455 25793 14467 25802
rect 10765 25759 10773 25793
rect 10829 25759 10865 25793
rect 10899 25759 10957 25793
rect 10991 25759 11049 25793
rect 11083 25759 11141 25793
rect 11175 25759 11233 25793
rect 11267 25759 11325 25793
rect 11359 25759 11417 25793
rect 11451 25759 11509 25793
rect 11543 25759 11601 25793
rect 11635 25759 11693 25793
rect 11727 25759 11785 25793
rect 11819 25759 11877 25793
rect 11911 25759 11969 25793
rect 12003 25759 12061 25793
rect 12095 25759 12153 25793
rect 12187 25759 12245 25793
rect 12279 25759 12337 25793
rect 12371 25759 12429 25793
rect 12463 25759 12521 25793
rect 12555 25759 12613 25793
rect 12647 25759 12705 25793
rect 12739 25759 12797 25793
rect 12831 25759 12889 25793
rect 12923 25759 12981 25793
rect 13015 25759 13073 25793
rect 13107 25759 13165 25793
rect 13199 25759 13257 25793
rect 13291 25759 13349 25793
rect 13383 25759 13441 25793
rect 13475 25759 13533 25793
rect 13567 25759 13625 25793
rect 13659 25759 13717 25793
rect 13751 25759 13809 25793
rect 13843 25759 13901 25793
rect 13935 25759 13993 25793
rect 14027 25759 14085 25793
rect 14119 25759 14177 25793
rect 14211 25759 14269 25793
rect 14303 25759 14339 25793
rect 14395 25759 14403 25793
rect 10701 25750 10713 25759
rect 10765 25750 10777 25759
rect 10829 25750 14339 25759
rect 14391 25750 14403 25759
rect 14455 25750 14467 25759
rect 14519 25750 14531 25802
rect 14583 25750 14595 25802
rect 14647 25793 18157 25802
rect 14671 25759 14729 25793
rect 14763 25759 14821 25793
rect 14855 25759 14913 25793
rect 14947 25759 15005 25793
rect 15039 25759 15097 25793
rect 15131 25759 15189 25793
rect 15223 25759 15281 25793
rect 15315 25759 15373 25793
rect 15407 25759 15465 25793
rect 15499 25759 15557 25793
rect 15591 25759 15649 25793
rect 15683 25759 15741 25793
rect 15775 25759 15833 25793
rect 15867 25759 15925 25793
rect 15959 25759 16017 25793
rect 16051 25759 16109 25793
rect 16143 25759 16201 25793
rect 16235 25759 16293 25793
rect 16327 25759 16385 25793
rect 16419 25759 16477 25793
rect 16511 25759 16569 25793
rect 16603 25759 16661 25793
rect 16695 25759 16753 25793
rect 16787 25759 16845 25793
rect 16879 25759 16937 25793
rect 16971 25759 17029 25793
rect 17063 25759 17121 25793
rect 17155 25759 17213 25793
rect 17247 25759 17305 25793
rect 17339 25759 17397 25793
rect 17431 25759 17489 25793
rect 17523 25759 17581 25793
rect 17615 25759 17673 25793
rect 17707 25759 17765 25793
rect 17799 25759 17857 25793
rect 17891 25759 17949 25793
rect 17983 25759 18041 25793
rect 18075 25759 18133 25793
rect 14647 25750 18157 25759
rect 18209 25750 18221 25802
rect 18273 25750 18285 25802
rect 18337 25793 18349 25802
rect 18401 25793 18413 25802
rect 18465 25793 20220 25802
rect 18401 25759 18409 25793
rect 18465 25759 18501 25793
rect 18535 25759 18593 25793
rect 18627 25759 18685 25793
rect 18719 25759 18777 25793
rect 18811 25759 18869 25793
rect 18903 25759 18961 25793
rect 18995 25759 19053 25793
rect 19087 25759 19145 25793
rect 19179 25759 19237 25793
rect 19271 25759 19329 25793
rect 19363 25759 19421 25793
rect 19455 25759 19513 25793
rect 19547 25759 19605 25793
rect 19639 25759 19697 25793
rect 19731 25759 19789 25793
rect 19823 25759 19881 25793
rect 19915 25759 19973 25793
rect 20007 25759 20065 25793
rect 20099 25759 20157 25793
rect 20191 25759 20220 25793
rect 18337 25750 18349 25759
rect 18401 25750 18413 25759
rect 18465 25750 20220 25759
rect 4948 25728 20220 25750
rect 14070 25308 14076 25360
rect 14128 25348 14134 25360
rect 14714 25348 14720 25360
rect 14128 25320 14720 25348
rect 14128 25308 14134 25320
rect 14714 25308 14720 25320
rect 14772 25308 14778 25360
rect 4948 25258 20220 25280
rect 4948 25249 6043 25258
rect 6095 25249 6107 25258
rect 4948 25215 4977 25249
rect 5011 25215 5069 25249
rect 5103 25215 5161 25249
rect 5195 25215 5253 25249
rect 5287 25215 5345 25249
rect 5379 25215 5437 25249
rect 5471 25215 5529 25249
rect 5563 25215 5621 25249
rect 5655 25215 5713 25249
rect 5747 25215 5805 25249
rect 5839 25215 5897 25249
rect 5931 25215 5989 25249
rect 6023 25215 6043 25249
rect 4948 25206 6043 25215
rect 6095 25206 6107 25215
rect 6159 25206 6171 25258
rect 6223 25206 6235 25258
rect 6287 25249 6299 25258
rect 6287 25206 6299 25215
rect 6351 25249 9861 25258
rect 6351 25215 6357 25249
rect 6391 25215 6449 25249
rect 6483 25215 6541 25249
rect 6575 25215 6633 25249
rect 6667 25215 6725 25249
rect 6759 25215 6817 25249
rect 6851 25215 6909 25249
rect 6943 25215 7001 25249
rect 7035 25215 7093 25249
rect 7127 25215 7185 25249
rect 7219 25215 7277 25249
rect 7311 25215 7369 25249
rect 7403 25215 7461 25249
rect 7495 25215 7553 25249
rect 7587 25215 7645 25249
rect 7679 25215 7737 25249
rect 7771 25215 7829 25249
rect 7863 25215 7921 25249
rect 7955 25215 8013 25249
rect 8047 25215 8105 25249
rect 8139 25215 8197 25249
rect 8231 25215 8289 25249
rect 8323 25215 8381 25249
rect 8415 25215 8473 25249
rect 8507 25215 8565 25249
rect 8599 25215 8657 25249
rect 8691 25215 8749 25249
rect 8783 25215 8841 25249
rect 8875 25215 8933 25249
rect 8967 25215 9025 25249
rect 9059 25215 9117 25249
rect 9151 25215 9209 25249
rect 9243 25215 9301 25249
rect 9335 25215 9393 25249
rect 9427 25215 9485 25249
rect 9519 25215 9577 25249
rect 9611 25215 9669 25249
rect 9703 25215 9761 25249
rect 9795 25215 9853 25249
rect 6351 25206 9861 25215
rect 9913 25206 9925 25258
rect 9977 25249 9989 25258
rect 10041 25249 10053 25258
rect 9979 25215 9989 25249
rect 9977 25206 9989 25215
rect 10041 25206 10053 25215
rect 10105 25206 10117 25258
rect 10169 25249 13679 25258
rect 13731 25249 13743 25258
rect 10169 25215 10221 25249
rect 10255 25215 10313 25249
rect 10347 25215 10405 25249
rect 10439 25215 10497 25249
rect 10531 25215 10589 25249
rect 10623 25215 10681 25249
rect 10715 25215 10773 25249
rect 10807 25215 10865 25249
rect 10899 25215 10957 25249
rect 10991 25215 11049 25249
rect 11083 25215 11141 25249
rect 11175 25215 11233 25249
rect 11267 25215 11325 25249
rect 11359 25215 11417 25249
rect 11451 25215 11509 25249
rect 11543 25215 11601 25249
rect 11635 25215 11693 25249
rect 11727 25215 11785 25249
rect 11819 25215 11877 25249
rect 11911 25215 11969 25249
rect 12003 25215 12061 25249
rect 12095 25215 12153 25249
rect 12187 25215 12245 25249
rect 12279 25215 12337 25249
rect 12371 25215 12429 25249
rect 12463 25215 12521 25249
rect 12555 25215 12613 25249
rect 12647 25215 12705 25249
rect 12739 25215 12797 25249
rect 12831 25215 12889 25249
rect 12923 25215 12981 25249
rect 13015 25215 13073 25249
rect 13107 25215 13165 25249
rect 13199 25215 13257 25249
rect 13291 25215 13349 25249
rect 13383 25215 13441 25249
rect 13475 25215 13533 25249
rect 13567 25215 13625 25249
rect 13659 25215 13679 25249
rect 10169 25206 13679 25215
rect 13731 25206 13743 25215
rect 13795 25206 13807 25258
rect 13859 25206 13871 25258
rect 13923 25249 13935 25258
rect 13923 25206 13935 25215
rect 13987 25249 17497 25258
rect 13987 25215 13993 25249
rect 14027 25215 14085 25249
rect 14119 25215 14177 25249
rect 14211 25215 14269 25249
rect 14303 25215 14361 25249
rect 14395 25215 14453 25249
rect 14487 25215 14545 25249
rect 14579 25215 14637 25249
rect 14671 25215 14729 25249
rect 14763 25215 14821 25249
rect 14855 25215 14913 25249
rect 14947 25215 15005 25249
rect 15039 25215 15097 25249
rect 15131 25215 15189 25249
rect 15223 25215 15281 25249
rect 15315 25215 15373 25249
rect 15407 25215 15465 25249
rect 15499 25215 15557 25249
rect 15591 25215 15649 25249
rect 15683 25215 15741 25249
rect 15775 25215 15833 25249
rect 15867 25215 15925 25249
rect 15959 25215 16017 25249
rect 16051 25215 16109 25249
rect 16143 25215 16201 25249
rect 16235 25215 16293 25249
rect 16327 25215 16385 25249
rect 16419 25215 16477 25249
rect 16511 25215 16569 25249
rect 16603 25215 16661 25249
rect 16695 25215 16753 25249
rect 16787 25215 16845 25249
rect 16879 25215 16937 25249
rect 16971 25215 17029 25249
rect 17063 25215 17121 25249
rect 17155 25215 17213 25249
rect 17247 25215 17305 25249
rect 17339 25215 17397 25249
rect 17431 25215 17489 25249
rect 13987 25206 17497 25215
rect 17549 25206 17561 25258
rect 17613 25249 17625 25258
rect 17677 25249 17689 25258
rect 17615 25215 17625 25249
rect 17613 25206 17625 25215
rect 17677 25206 17689 25215
rect 17741 25206 17753 25258
rect 17805 25249 20220 25258
rect 17805 25215 17857 25249
rect 17891 25215 17949 25249
rect 17983 25215 18041 25249
rect 18075 25215 18133 25249
rect 18167 25215 18225 25249
rect 18259 25215 18317 25249
rect 18351 25215 18409 25249
rect 18443 25215 18501 25249
rect 18535 25215 18593 25249
rect 18627 25215 18685 25249
rect 18719 25215 18777 25249
rect 18811 25215 18869 25249
rect 18903 25215 18961 25249
rect 18995 25215 19053 25249
rect 19087 25215 19145 25249
rect 19179 25215 19237 25249
rect 19271 25215 19329 25249
rect 19363 25215 19421 25249
rect 19455 25215 19513 25249
rect 19547 25215 19605 25249
rect 19639 25215 19697 25249
rect 19731 25215 19789 25249
rect 19823 25215 19881 25249
rect 19915 25215 19973 25249
rect 20007 25215 20065 25249
rect 20099 25215 20157 25249
rect 20191 25215 20220 25249
rect 17805 25206 20220 25215
rect 4948 25184 20220 25206
rect 4948 24714 20220 24736
rect 4948 24705 6703 24714
rect 6755 24705 6767 24714
rect 6819 24705 6831 24714
rect 4948 24671 4977 24705
rect 5011 24671 5069 24705
rect 5103 24671 5161 24705
rect 5195 24671 5253 24705
rect 5287 24671 5345 24705
rect 5379 24671 5437 24705
rect 5471 24671 5529 24705
rect 5563 24671 5621 24705
rect 5655 24671 5713 24705
rect 5747 24671 5805 24705
rect 5839 24671 5897 24705
rect 5931 24671 5989 24705
rect 6023 24671 6081 24705
rect 6115 24671 6173 24705
rect 6207 24671 6265 24705
rect 6299 24671 6357 24705
rect 6391 24671 6449 24705
rect 6483 24671 6541 24705
rect 6575 24671 6633 24705
rect 6667 24671 6703 24705
rect 6759 24671 6767 24705
rect 4948 24662 6703 24671
rect 6755 24662 6767 24671
rect 6819 24662 6831 24671
rect 6883 24662 6895 24714
rect 6947 24662 6959 24714
rect 7011 24705 10521 24714
rect 7035 24671 7093 24705
rect 7127 24671 7185 24705
rect 7219 24671 7277 24705
rect 7311 24671 7369 24705
rect 7403 24671 7461 24705
rect 7495 24671 7553 24705
rect 7587 24671 7645 24705
rect 7679 24671 7737 24705
rect 7771 24671 7829 24705
rect 7863 24671 7921 24705
rect 7955 24671 8013 24705
rect 8047 24671 8105 24705
rect 8139 24671 8197 24705
rect 8231 24671 8289 24705
rect 8323 24671 8381 24705
rect 8415 24671 8473 24705
rect 8507 24671 8565 24705
rect 8599 24671 8657 24705
rect 8691 24671 8749 24705
rect 8783 24671 8841 24705
rect 8875 24671 8933 24705
rect 8967 24671 9025 24705
rect 9059 24671 9117 24705
rect 9151 24671 9209 24705
rect 9243 24671 9301 24705
rect 9335 24671 9393 24705
rect 9427 24671 9485 24705
rect 9519 24671 9577 24705
rect 9611 24671 9669 24705
rect 9703 24671 9761 24705
rect 9795 24671 9853 24705
rect 9887 24671 9945 24705
rect 9979 24671 10037 24705
rect 10071 24671 10129 24705
rect 10163 24671 10221 24705
rect 10255 24671 10313 24705
rect 10347 24671 10405 24705
rect 10439 24671 10497 24705
rect 7011 24662 10521 24671
rect 10573 24662 10585 24714
rect 10637 24662 10649 24714
rect 10701 24705 10713 24714
rect 10765 24705 10777 24714
rect 10829 24705 14339 24714
rect 14391 24705 14403 24714
rect 14455 24705 14467 24714
rect 10765 24671 10773 24705
rect 10829 24671 10865 24705
rect 10899 24671 10957 24705
rect 10991 24671 11049 24705
rect 11083 24671 11141 24705
rect 11175 24671 11233 24705
rect 11267 24671 11325 24705
rect 11359 24671 11417 24705
rect 11451 24671 11509 24705
rect 11543 24671 11601 24705
rect 11635 24671 11693 24705
rect 11727 24671 11785 24705
rect 11819 24671 11877 24705
rect 11911 24671 11969 24705
rect 12003 24671 12061 24705
rect 12095 24671 12153 24705
rect 12187 24671 12245 24705
rect 12279 24671 12337 24705
rect 12371 24671 12429 24705
rect 12463 24671 12521 24705
rect 12555 24671 12613 24705
rect 12647 24671 12705 24705
rect 12739 24671 12797 24705
rect 12831 24671 12889 24705
rect 12923 24671 12981 24705
rect 13015 24671 13073 24705
rect 13107 24671 13165 24705
rect 13199 24671 13257 24705
rect 13291 24671 13349 24705
rect 13383 24671 13441 24705
rect 13475 24671 13533 24705
rect 13567 24671 13625 24705
rect 13659 24671 13717 24705
rect 13751 24671 13809 24705
rect 13843 24671 13901 24705
rect 13935 24671 13993 24705
rect 14027 24671 14085 24705
rect 14119 24671 14177 24705
rect 14211 24671 14269 24705
rect 14303 24671 14339 24705
rect 14395 24671 14403 24705
rect 10701 24662 10713 24671
rect 10765 24662 10777 24671
rect 10829 24662 14339 24671
rect 14391 24662 14403 24671
rect 14455 24662 14467 24671
rect 14519 24662 14531 24714
rect 14583 24662 14595 24714
rect 14647 24705 18157 24714
rect 14671 24671 14729 24705
rect 14763 24671 14821 24705
rect 14855 24671 14913 24705
rect 14947 24671 15005 24705
rect 15039 24671 15097 24705
rect 15131 24671 15189 24705
rect 15223 24671 15281 24705
rect 15315 24671 15373 24705
rect 15407 24671 15465 24705
rect 15499 24671 15557 24705
rect 15591 24671 15649 24705
rect 15683 24671 15741 24705
rect 15775 24671 15833 24705
rect 15867 24671 15925 24705
rect 15959 24671 16017 24705
rect 16051 24671 16109 24705
rect 16143 24671 16201 24705
rect 16235 24671 16293 24705
rect 16327 24671 16385 24705
rect 16419 24671 16477 24705
rect 16511 24671 16569 24705
rect 16603 24671 16661 24705
rect 16695 24671 16753 24705
rect 16787 24671 16845 24705
rect 16879 24671 16937 24705
rect 16971 24671 17029 24705
rect 17063 24671 17121 24705
rect 17155 24671 17213 24705
rect 17247 24671 17305 24705
rect 17339 24671 17397 24705
rect 17431 24671 17489 24705
rect 17523 24671 17581 24705
rect 17615 24671 17673 24705
rect 17707 24671 17765 24705
rect 17799 24671 17857 24705
rect 17891 24671 17949 24705
rect 17983 24671 18041 24705
rect 18075 24671 18133 24705
rect 14647 24662 18157 24671
rect 18209 24662 18221 24714
rect 18273 24662 18285 24714
rect 18337 24705 18349 24714
rect 18401 24705 18413 24714
rect 18465 24705 20220 24714
rect 18401 24671 18409 24705
rect 18465 24671 18501 24705
rect 18535 24671 18593 24705
rect 18627 24671 18685 24705
rect 18719 24671 18777 24705
rect 18811 24671 18869 24705
rect 18903 24671 18961 24705
rect 18995 24671 19053 24705
rect 19087 24671 19145 24705
rect 19179 24671 19237 24705
rect 19271 24671 19329 24705
rect 19363 24671 19421 24705
rect 19455 24671 19513 24705
rect 19547 24671 19605 24705
rect 19639 24671 19697 24705
rect 19731 24671 19789 24705
rect 19823 24671 19881 24705
rect 19915 24671 19973 24705
rect 20007 24671 20065 24705
rect 20099 24671 20157 24705
rect 20191 24671 20220 24705
rect 18337 24662 18349 24671
rect 18401 24662 18413 24671
rect 18465 24662 20220 24671
rect 4948 24640 20220 24662
rect 4948 24170 20220 24192
rect 4948 24161 6043 24170
rect 6095 24161 6107 24170
rect 4948 24127 4977 24161
rect 5011 24127 5069 24161
rect 5103 24127 5161 24161
rect 5195 24127 5253 24161
rect 5287 24127 5345 24161
rect 5379 24127 5437 24161
rect 5471 24127 5529 24161
rect 5563 24127 5621 24161
rect 5655 24127 5713 24161
rect 5747 24127 5805 24161
rect 5839 24127 5897 24161
rect 5931 24127 5989 24161
rect 6023 24127 6043 24161
rect 4948 24118 6043 24127
rect 6095 24118 6107 24127
rect 6159 24118 6171 24170
rect 6223 24118 6235 24170
rect 6287 24161 6299 24170
rect 6287 24118 6299 24127
rect 6351 24161 9861 24170
rect 6351 24127 6357 24161
rect 6391 24127 6449 24161
rect 6483 24127 6541 24161
rect 6575 24127 6633 24161
rect 6667 24127 6725 24161
rect 6759 24127 6817 24161
rect 6851 24127 6909 24161
rect 6943 24127 7001 24161
rect 7035 24127 7093 24161
rect 7127 24127 7185 24161
rect 7219 24127 7277 24161
rect 7311 24127 7369 24161
rect 7403 24127 7461 24161
rect 7495 24127 7553 24161
rect 7587 24127 7645 24161
rect 7679 24127 7737 24161
rect 7771 24127 7829 24161
rect 7863 24127 7921 24161
rect 7955 24127 8013 24161
rect 8047 24127 8105 24161
rect 8139 24127 8197 24161
rect 8231 24127 8289 24161
rect 8323 24127 8381 24161
rect 8415 24127 8473 24161
rect 8507 24127 8565 24161
rect 8599 24127 8657 24161
rect 8691 24127 8749 24161
rect 8783 24127 8841 24161
rect 8875 24127 8933 24161
rect 8967 24127 9025 24161
rect 9059 24127 9117 24161
rect 9151 24127 9209 24161
rect 9243 24127 9301 24161
rect 9335 24127 9393 24161
rect 9427 24127 9485 24161
rect 9519 24127 9577 24161
rect 9611 24127 9669 24161
rect 9703 24127 9761 24161
rect 9795 24127 9853 24161
rect 6351 24118 9861 24127
rect 9913 24118 9925 24170
rect 9977 24161 9989 24170
rect 10041 24161 10053 24170
rect 9979 24127 9989 24161
rect 9977 24118 9989 24127
rect 10041 24118 10053 24127
rect 10105 24118 10117 24170
rect 10169 24161 13679 24170
rect 13731 24161 13743 24170
rect 10169 24127 10221 24161
rect 10255 24127 10313 24161
rect 10347 24127 10405 24161
rect 10439 24127 10497 24161
rect 10531 24127 10589 24161
rect 10623 24127 10681 24161
rect 10715 24127 10773 24161
rect 10807 24127 10865 24161
rect 10899 24127 10957 24161
rect 10991 24127 11049 24161
rect 11083 24127 11141 24161
rect 11175 24127 11233 24161
rect 11267 24127 11325 24161
rect 11359 24127 11417 24161
rect 11451 24127 11509 24161
rect 11543 24127 11601 24161
rect 11635 24127 11693 24161
rect 11727 24127 11785 24161
rect 11819 24127 11877 24161
rect 11911 24127 11969 24161
rect 12003 24127 12061 24161
rect 12095 24127 12153 24161
rect 12187 24127 12245 24161
rect 12279 24127 12337 24161
rect 12371 24127 12429 24161
rect 12463 24127 12521 24161
rect 12555 24127 12613 24161
rect 12647 24127 12705 24161
rect 12739 24127 12797 24161
rect 12831 24127 12889 24161
rect 12923 24127 12981 24161
rect 13015 24127 13073 24161
rect 13107 24127 13165 24161
rect 13199 24127 13257 24161
rect 13291 24127 13349 24161
rect 13383 24127 13441 24161
rect 13475 24127 13533 24161
rect 13567 24127 13625 24161
rect 13659 24127 13679 24161
rect 10169 24118 13679 24127
rect 13731 24118 13743 24127
rect 13795 24118 13807 24170
rect 13859 24118 13871 24170
rect 13923 24161 13935 24170
rect 13923 24118 13935 24127
rect 13987 24161 17497 24170
rect 13987 24127 13993 24161
rect 14027 24127 14085 24161
rect 14119 24127 14177 24161
rect 14211 24127 14269 24161
rect 14303 24127 14361 24161
rect 14395 24127 14453 24161
rect 14487 24127 14545 24161
rect 14579 24127 14637 24161
rect 14671 24127 14729 24161
rect 14763 24127 14821 24161
rect 14855 24127 14913 24161
rect 14947 24127 15005 24161
rect 15039 24127 15097 24161
rect 15131 24127 15189 24161
rect 15223 24127 15281 24161
rect 15315 24127 15373 24161
rect 15407 24127 15465 24161
rect 15499 24127 15557 24161
rect 15591 24127 15649 24161
rect 15683 24127 15741 24161
rect 15775 24127 15833 24161
rect 15867 24127 15925 24161
rect 15959 24127 16017 24161
rect 16051 24127 16109 24161
rect 16143 24127 16201 24161
rect 16235 24127 16293 24161
rect 16327 24127 16385 24161
rect 16419 24127 16477 24161
rect 16511 24127 16569 24161
rect 16603 24127 16661 24161
rect 16695 24127 16753 24161
rect 16787 24127 16845 24161
rect 16879 24127 16937 24161
rect 16971 24127 17029 24161
rect 17063 24127 17121 24161
rect 17155 24127 17213 24161
rect 17247 24127 17305 24161
rect 17339 24127 17397 24161
rect 17431 24127 17489 24161
rect 13987 24118 17497 24127
rect 17549 24118 17561 24170
rect 17613 24161 17625 24170
rect 17677 24161 17689 24170
rect 17615 24127 17625 24161
rect 17613 24118 17625 24127
rect 17677 24118 17689 24127
rect 17741 24118 17753 24170
rect 17805 24161 20220 24170
rect 17805 24127 17857 24161
rect 17891 24127 17949 24161
rect 17983 24127 18041 24161
rect 18075 24127 18133 24161
rect 18167 24127 18225 24161
rect 18259 24127 18317 24161
rect 18351 24127 18409 24161
rect 18443 24127 18501 24161
rect 18535 24127 18593 24161
rect 18627 24127 18685 24161
rect 18719 24127 18777 24161
rect 18811 24127 18869 24161
rect 18903 24127 18961 24161
rect 18995 24127 19053 24161
rect 19087 24127 19145 24161
rect 19179 24127 19237 24161
rect 19271 24127 19329 24161
rect 19363 24127 19421 24161
rect 19455 24127 19513 24161
rect 19547 24127 19605 24161
rect 19639 24127 19697 24161
rect 19731 24127 19789 24161
rect 19823 24127 19881 24161
rect 19915 24127 19973 24161
rect 20007 24127 20065 24161
rect 20099 24127 20157 24161
rect 20191 24127 20220 24161
rect 17805 24118 20220 24127
rect 4948 24096 20220 24118
rect 4948 23626 20220 23648
rect 4948 23617 6703 23626
rect 6755 23617 6767 23626
rect 6819 23617 6831 23626
rect 4948 23583 4977 23617
rect 5011 23583 5069 23617
rect 5103 23583 5161 23617
rect 5195 23583 5253 23617
rect 5287 23583 5345 23617
rect 5379 23583 5437 23617
rect 5471 23583 5529 23617
rect 5563 23583 5621 23617
rect 5655 23583 5713 23617
rect 5747 23583 5805 23617
rect 5839 23583 5897 23617
rect 5931 23583 5989 23617
rect 6023 23583 6081 23617
rect 6115 23583 6173 23617
rect 6207 23583 6265 23617
rect 6299 23583 6357 23617
rect 6391 23583 6449 23617
rect 6483 23583 6541 23617
rect 6575 23583 6633 23617
rect 6667 23583 6703 23617
rect 6759 23583 6767 23617
rect 4948 23574 6703 23583
rect 6755 23574 6767 23583
rect 6819 23574 6831 23583
rect 6883 23574 6895 23626
rect 6947 23574 6959 23626
rect 7011 23617 10521 23626
rect 7035 23583 7093 23617
rect 7127 23583 7185 23617
rect 7219 23583 7277 23617
rect 7311 23583 7369 23617
rect 7403 23583 7461 23617
rect 7495 23583 7553 23617
rect 7587 23583 7645 23617
rect 7679 23583 7737 23617
rect 7771 23583 7829 23617
rect 7863 23583 7921 23617
rect 7955 23583 8013 23617
rect 8047 23583 8105 23617
rect 8139 23583 8197 23617
rect 8231 23583 8289 23617
rect 8323 23583 8381 23617
rect 8415 23583 8473 23617
rect 8507 23583 8565 23617
rect 8599 23583 8657 23617
rect 8691 23583 8749 23617
rect 8783 23583 8841 23617
rect 8875 23583 8933 23617
rect 8967 23583 9025 23617
rect 9059 23583 9117 23617
rect 9151 23583 9209 23617
rect 9243 23583 9301 23617
rect 9335 23583 9393 23617
rect 9427 23583 9485 23617
rect 9519 23583 9577 23617
rect 9611 23583 9669 23617
rect 9703 23583 9761 23617
rect 9795 23583 9853 23617
rect 9887 23583 9945 23617
rect 9979 23583 10037 23617
rect 10071 23583 10129 23617
rect 10163 23583 10221 23617
rect 10255 23583 10313 23617
rect 10347 23583 10405 23617
rect 10439 23583 10497 23617
rect 7011 23574 10521 23583
rect 10573 23574 10585 23626
rect 10637 23574 10649 23626
rect 10701 23617 10713 23626
rect 10765 23617 10777 23626
rect 10829 23617 14339 23626
rect 14391 23617 14403 23626
rect 14455 23617 14467 23626
rect 10765 23583 10773 23617
rect 10829 23583 10865 23617
rect 10899 23583 10957 23617
rect 10991 23583 11049 23617
rect 11083 23583 11141 23617
rect 11175 23583 11233 23617
rect 11267 23583 11325 23617
rect 11359 23583 11417 23617
rect 11451 23583 11509 23617
rect 11543 23583 11601 23617
rect 11635 23583 11693 23617
rect 11727 23583 11785 23617
rect 11819 23583 11877 23617
rect 11911 23583 11969 23617
rect 12003 23583 12061 23617
rect 12095 23583 12153 23617
rect 12187 23583 12245 23617
rect 12279 23583 12337 23617
rect 12371 23583 12429 23617
rect 12463 23583 12521 23617
rect 12555 23583 12613 23617
rect 12647 23583 12705 23617
rect 12739 23583 12797 23617
rect 12831 23583 12889 23617
rect 12923 23583 12981 23617
rect 13015 23583 13073 23617
rect 13107 23583 13165 23617
rect 13199 23583 13257 23617
rect 13291 23583 13349 23617
rect 13383 23583 13441 23617
rect 13475 23583 13533 23617
rect 13567 23583 13625 23617
rect 13659 23583 13717 23617
rect 13751 23583 13809 23617
rect 13843 23583 13901 23617
rect 13935 23583 13993 23617
rect 14027 23583 14085 23617
rect 14119 23583 14177 23617
rect 14211 23583 14269 23617
rect 14303 23583 14339 23617
rect 14395 23583 14403 23617
rect 10701 23574 10713 23583
rect 10765 23574 10777 23583
rect 10829 23574 14339 23583
rect 14391 23574 14403 23583
rect 14455 23574 14467 23583
rect 14519 23574 14531 23626
rect 14583 23574 14595 23626
rect 14647 23617 18157 23626
rect 14671 23583 14729 23617
rect 14763 23583 14821 23617
rect 14855 23583 14913 23617
rect 14947 23583 15005 23617
rect 15039 23583 15097 23617
rect 15131 23583 15189 23617
rect 15223 23583 15281 23617
rect 15315 23583 15373 23617
rect 15407 23583 15465 23617
rect 15499 23583 15557 23617
rect 15591 23583 15649 23617
rect 15683 23583 15741 23617
rect 15775 23583 15833 23617
rect 15867 23583 15925 23617
rect 15959 23583 16017 23617
rect 16051 23583 16109 23617
rect 16143 23583 16201 23617
rect 16235 23583 16293 23617
rect 16327 23583 16385 23617
rect 16419 23583 16477 23617
rect 16511 23583 16569 23617
rect 16603 23583 16661 23617
rect 16695 23583 16753 23617
rect 16787 23583 16845 23617
rect 16879 23583 16937 23617
rect 16971 23583 17029 23617
rect 17063 23583 17121 23617
rect 17155 23583 17213 23617
rect 17247 23583 17305 23617
rect 17339 23583 17397 23617
rect 17431 23583 17489 23617
rect 17523 23583 17581 23617
rect 17615 23583 17673 23617
rect 17707 23583 17765 23617
rect 17799 23583 17857 23617
rect 17891 23583 17949 23617
rect 17983 23583 18041 23617
rect 18075 23583 18133 23617
rect 14647 23574 18157 23583
rect 18209 23574 18221 23626
rect 18273 23574 18285 23626
rect 18337 23617 18349 23626
rect 18401 23617 18413 23626
rect 18465 23617 20220 23626
rect 18401 23583 18409 23617
rect 18465 23583 18501 23617
rect 18535 23583 18593 23617
rect 18627 23583 18685 23617
rect 18719 23583 18777 23617
rect 18811 23583 18869 23617
rect 18903 23583 18961 23617
rect 18995 23583 19053 23617
rect 19087 23583 19145 23617
rect 19179 23583 19237 23617
rect 19271 23583 19329 23617
rect 19363 23583 19421 23617
rect 19455 23583 19513 23617
rect 19547 23583 19605 23617
rect 19639 23583 19697 23617
rect 19731 23583 19789 23617
rect 19823 23583 19881 23617
rect 19915 23583 19973 23617
rect 20007 23583 20065 23617
rect 20099 23583 20157 23617
rect 20191 23583 20220 23617
rect 18337 23574 18349 23583
rect 18401 23574 18413 23583
rect 18465 23574 20220 23583
rect 4948 23552 20220 23574
rect 4948 23082 20220 23104
rect 4948 23073 6043 23082
rect 6095 23073 6107 23082
rect 4948 23039 4977 23073
rect 5011 23039 5069 23073
rect 5103 23039 5161 23073
rect 5195 23039 5253 23073
rect 5287 23039 5345 23073
rect 5379 23039 5437 23073
rect 5471 23039 5529 23073
rect 5563 23039 5621 23073
rect 5655 23039 5713 23073
rect 5747 23039 5805 23073
rect 5839 23039 5897 23073
rect 5931 23039 5989 23073
rect 6023 23039 6043 23073
rect 4948 23030 6043 23039
rect 6095 23030 6107 23039
rect 6159 23030 6171 23082
rect 6223 23030 6235 23082
rect 6287 23073 6299 23082
rect 6287 23030 6299 23039
rect 6351 23073 9861 23082
rect 6351 23039 6357 23073
rect 6391 23039 6449 23073
rect 6483 23039 6541 23073
rect 6575 23039 6633 23073
rect 6667 23039 6725 23073
rect 6759 23039 6817 23073
rect 6851 23039 6909 23073
rect 6943 23039 7001 23073
rect 7035 23039 7093 23073
rect 7127 23039 7185 23073
rect 7219 23039 7277 23073
rect 7311 23039 7369 23073
rect 7403 23039 7461 23073
rect 7495 23039 7553 23073
rect 7587 23039 7645 23073
rect 7679 23039 7737 23073
rect 7771 23039 7829 23073
rect 7863 23039 7921 23073
rect 7955 23039 8013 23073
rect 8047 23039 8105 23073
rect 8139 23039 8197 23073
rect 8231 23039 8289 23073
rect 8323 23039 8381 23073
rect 8415 23039 8473 23073
rect 8507 23039 8565 23073
rect 8599 23039 8657 23073
rect 8691 23039 8749 23073
rect 8783 23039 8841 23073
rect 8875 23039 8933 23073
rect 8967 23039 9025 23073
rect 9059 23039 9117 23073
rect 9151 23039 9209 23073
rect 9243 23039 9301 23073
rect 9335 23039 9393 23073
rect 9427 23039 9485 23073
rect 9519 23039 9577 23073
rect 9611 23039 9669 23073
rect 9703 23039 9761 23073
rect 9795 23039 9853 23073
rect 6351 23030 9861 23039
rect 9913 23030 9925 23082
rect 9977 23073 9989 23082
rect 10041 23073 10053 23082
rect 9979 23039 9989 23073
rect 9977 23030 9989 23039
rect 10041 23030 10053 23039
rect 10105 23030 10117 23082
rect 10169 23073 13679 23082
rect 13731 23073 13743 23082
rect 10169 23039 10221 23073
rect 10255 23039 10313 23073
rect 10347 23039 10405 23073
rect 10439 23039 10497 23073
rect 10531 23039 10589 23073
rect 10623 23039 10681 23073
rect 10715 23039 10773 23073
rect 10807 23039 10865 23073
rect 10899 23039 10957 23073
rect 10991 23039 11049 23073
rect 11083 23039 11141 23073
rect 11175 23039 11233 23073
rect 11267 23039 11325 23073
rect 11359 23039 11417 23073
rect 11451 23039 11509 23073
rect 11543 23039 11601 23073
rect 11635 23039 11693 23073
rect 11727 23039 11785 23073
rect 11819 23039 11877 23073
rect 11911 23039 11969 23073
rect 12003 23039 12061 23073
rect 12095 23039 12153 23073
rect 12187 23039 12245 23073
rect 12279 23039 12337 23073
rect 12371 23039 12429 23073
rect 12463 23039 12521 23073
rect 12555 23039 12613 23073
rect 12647 23039 12705 23073
rect 12739 23039 12797 23073
rect 12831 23039 12889 23073
rect 12923 23039 12981 23073
rect 13015 23039 13073 23073
rect 13107 23039 13165 23073
rect 13199 23039 13257 23073
rect 13291 23039 13349 23073
rect 13383 23039 13441 23073
rect 13475 23039 13533 23073
rect 13567 23039 13625 23073
rect 13659 23039 13679 23073
rect 10169 23030 13679 23039
rect 13731 23030 13743 23039
rect 13795 23030 13807 23082
rect 13859 23030 13871 23082
rect 13923 23073 13935 23082
rect 13923 23030 13935 23039
rect 13987 23073 17497 23082
rect 13987 23039 13993 23073
rect 14027 23039 14085 23073
rect 14119 23039 14177 23073
rect 14211 23039 14269 23073
rect 14303 23039 14361 23073
rect 14395 23039 14453 23073
rect 14487 23039 14545 23073
rect 14579 23039 14637 23073
rect 14671 23039 14729 23073
rect 14763 23039 14821 23073
rect 14855 23039 14913 23073
rect 14947 23039 15005 23073
rect 15039 23039 15097 23073
rect 15131 23039 15189 23073
rect 15223 23039 15281 23073
rect 15315 23039 15373 23073
rect 15407 23039 15465 23073
rect 15499 23039 15557 23073
rect 15591 23039 15649 23073
rect 15683 23039 15741 23073
rect 15775 23039 15833 23073
rect 15867 23039 15925 23073
rect 15959 23039 16017 23073
rect 16051 23039 16109 23073
rect 16143 23039 16201 23073
rect 16235 23039 16293 23073
rect 16327 23039 16385 23073
rect 16419 23039 16477 23073
rect 16511 23039 16569 23073
rect 16603 23039 16661 23073
rect 16695 23039 16753 23073
rect 16787 23039 16845 23073
rect 16879 23039 16937 23073
rect 16971 23039 17029 23073
rect 17063 23039 17121 23073
rect 17155 23039 17213 23073
rect 17247 23039 17305 23073
rect 17339 23039 17397 23073
rect 17431 23039 17489 23073
rect 13987 23030 17497 23039
rect 17549 23030 17561 23082
rect 17613 23073 17625 23082
rect 17677 23073 17689 23082
rect 17615 23039 17625 23073
rect 17613 23030 17625 23039
rect 17677 23030 17689 23039
rect 17741 23030 17753 23082
rect 17805 23073 20220 23082
rect 17805 23039 17857 23073
rect 17891 23039 17949 23073
rect 17983 23039 18041 23073
rect 18075 23039 18133 23073
rect 18167 23039 18225 23073
rect 18259 23039 18317 23073
rect 18351 23039 18409 23073
rect 18443 23039 18501 23073
rect 18535 23039 18593 23073
rect 18627 23039 18685 23073
rect 18719 23039 18777 23073
rect 18811 23039 18869 23073
rect 18903 23039 18961 23073
rect 18995 23039 19053 23073
rect 19087 23039 19145 23073
rect 19179 23039 19237 23073
rect 19271 23039 19329 23073
rect 19363 23039 19421 23073
rect 19455 23039 19513 23073
rect 19547 23039 19605 23073
rect 19639 23039 19697 23073
rect 19731 23039 19789 23073
rect 19823 23039 19881 23073
rect 19915 23039 19973 23073
rect 20007 23039 20065 23073
rect 20099 23039 20157 23073
rect 20191 23039 20220 23073
rect 17805 23030 20220 23039
rect 4948 23008 20220 23030
rect 4948 22538 20220 22560
rect 4948 22529 6703 22538
rect 6755 22529 6767 22538
rect 6819 22529 6831 22538
rect 4948 22495 4977 22529
rect 5011 22495 5069 22529
rect 5103 22495 5161 22529
rect 5195 22495 5253 22529
rect 5287 22495 5345 22529
rect 5379 22495 5437 22529
rect 5471 22495 5529 22529
rect 5563 22495 5621 22529
rect 5655 22495 5713 22529
rect 5747 22495 5805 22529
rect 5839 22495 5897 22529
rect 5931 22495 5989 22529
rect 6023 22495 6081 22529
rect 6115 22495 6173 22529
rect 6207 22495 6265 22529
rect 6299 22495 6357 22529
rect 6391 22495 6449 22529
rect 6483 22495 6541 22529
rect 6575 22495 6633 22529
rect 6667 22495 6703 22529
rect 6759 22495 6767 22529
rect 4948 22486 6703 22495
rect 6755 22486 6767 22495
rect 6819 22486 6831 22495
rect 6883 22486 6895 22538
rect 6947 22486 6959 22538
rect 7011 22529 10521 22538
rect 7035 22495 7093 22529
rect 7127 22495 7185 22529
rect 7219 22495 7277 22529
rect 7311 22495 7369 22529
rect 7403 22495 7461 22529
rect 7495 22495 7553 22529
rect 7587 22495 7645 22529
rect 7679 22495 7737 22529
rect 7771 22495 7829 22529
rect 7863 22495 7921 22529
rect 7955 22495 8013 22529
rect 8047 22495 8105 22529
rect 8139 22495 8197 22529
rect 8231 22495 8289 22529
rect 8323 22495 8381 22529
rect 8415 22495 8473 22529
rect 8507 22495 8565 22529
rect 8599 22495 8657 22529
rect 8691 22495 8749 22529
rect 8783 22495 8841 22529
rect 8875 22495 8933 22529
rect 8967 22495 9025 22529
rect 9059 22495 9117 22529
rect 9151 22495 9209 22529
rect 9243 22495 9301 22529
rect 9335 22495 9393 22529
rect 9427 22495 9485 22529
rect 9519 22495 9577 22529
rect 9611 22495 9669 22529
rect 9703 22495 9761 22529
rect 9795 22495 9853 22529
rect 9887 22495 9945 22529
rect 9979 22495 10037 22529
rect 10071 22495 10129 22529
rect 10163 22495 10221 22529
rect 10255 22495 10313 22529
rect 10347 22495 10405 22529
rect 10439 22495 10497 22529
rect 7011 22486 10521 22495
rect 10573 22486 10585 22538
rect 10637 22486 10649 22538
rect 10701 22529 10713 22538
rect 10765 22529 10777 22538
rect 10829 22529 14339 22538
rect 14391 22529 14403 22538
rect 14455 22529 14467 22538
rect 10765 22495 10773 22529
rect 10829 22495 10865 22529
rect 10899 22495 10957 22529
rect 10991 22495 11049 22529
rect 11083 22495 11141 22529
rect 11175 22495 11233 22529
rect 11267 22495 11325 22529
rect 11359 22495 11417 22529
rect 11451 22495 11509 22529
rect 11543 22495 11601 22529
rect 11635 22495 11693 22529
rect 11727 22495 11785 22529
rect 11819 22495 11877 22529
rect 11911 22495 11969 22529
rect 12003 22495 12061 22529
rect 12095 22495 12153 22529
rect 12187 22495 12245 22529
rect 12279 22495 12337 22529
rect 12371 22495 12429 22529
rect 12463 22495 12521 22529
rect 12555 22495 12613 22529
rect 12647 22495 12705 22529
rect 12739 22495 12797 22529
rect 12831 22495 12889 22529
rect 12923 22495 12981 22529
rect 13015 22495 13073 22529
rect 13107 22495 13165 22529
rect 13199 22495 13257 22529
rect 13291 22495 13349 22529
rect 13383 22495 13441 22529
rect 13475 22495 13533 22529
rect 13567 22495 13625 22529
rect 13659 22495 13717 22529
rect 13751 22495 13809 22529
rect 13843 22495 13901 22529
rect 13935 22495 13993 22529
rect 14027 22495 14085 22529
rect 14119 22495 14177 22529
rect 14211 22495 14269 22529
rect 14303 22495 14339 22529
rect 14395 22495 14403 22529
rect 10701 22486 10713 22495
rect 10765 22486 10777 22495
rect 10829 22486 14339 22495
rect 14391 22486 14403 22495
rect 14455 22486 14467 22495
rect 14519 22486 14531 22538
rect 14583 22486 14595 22538
rect 14647 22529 18157 22538
rect 14671 22495 14729 22529
rect 14763 22495 14821 22529
rect 14855 22495 14913 22529
rect 14947 22495 15005 22529
rect 15039 22495 15097 22529
rect 15131 22495 15189 22529
rect 15223 22495 15281 22529
rect 15315 22495 15373 22529
rect 15407 22495 15465 22529
rect 15499 22495 15557 22529
rect 15591 22495 15649 22529
rect 15683 22495 15741 22529
rect 15775 22495 15833 22529
rect 15867 22495 15925 22529
rect 15959 22495 16017 22529
rect 16051 22495 16109 22529
rect 16143 22495 16201 22529
rect 16235 22495 16293 22529
rect 16327 22495 16385 22529
rect 16419 22495 16477 22529
rect 16511 22495 16569 22529
rect 16603 22495 16661 22529
rect 16695 22495 16753 22529
rect 16787 22495 16845 22529
rect 16879 22495 16937 22529
rect 16971 22495 17029 22529
rect 17063 22495 17121 22529
rect 17155 22495 17213 22529
rect 17247 22495 17305 22529
rect 17339 22495 17397 22529
rect 17431 22495 17489 22529
rect 17523 22495 17581 22529
rect 17615 22495 17673 22529
rect 17707 22495 17765 22529
rect 17799 22495 17857 22529
rect 17891 22495 17949 22529
rect 17983 22495 18041 22529
rect 18075 22495 18133 22529
rect 14647 22486 18157 22495
rect 18209 22486 18221 22538
rect 18273 22486 18285 22538
rect 18337 22529 18349 22538
rect 18401 22529 18413 22538
rect 18465 22529 20220 22538
rect 18401 22495 18409 22529
rect 18465 22495 18501 22529
rect 18535 22495 18593 22529
rect 18627 22495 18685 22529
rect 18719 22495 18777 22529
rect 18811 22495 18869 22529
rect 18903 22495 18961 22529
rect 18995 22495 19053 22529
rect 19087 22495 19145 22529
rect 19179 22495 19237 22529
rect 19271 22495 19329 22529
rect 19363 22495 19421 22529
rect 19455 22495 19513 22529
rect 19547 22495 19605 22529
rect 19639 22495 19697 22529
rect 19731 22495 19789 22529
rect 19823 22495 19881 22529
rect 19915 22495 19973 22529
rect 20007 22495 20065 22529
rect 20099 22495 20157 22529
rect 20191 22495 20220 22529
rect 18337 22486 18349 22495
rect 18401 22486 18413 22495
rect 18465 22486 20220 22495
rect 4948 22464 20220 22486
rect 4948 21994 20220 22016
rect 4948 21985 6043 21994
rect 6095 21985 6107 21994
rect 4948 21951 4977 21985
rect 5011 21951 5069 21985
rect 5103 21951 5161 21985
rect 5195 21951 5253 21985
rect 5287 21951 5345 21985
rect 5379 21951 5437 21985
rect 5471 21951 5529 21985
rect 5563 21951 5621 21985
rect 5655 21951 5713 21985
rect 5747 21951 5805 21985
rect 5839 21951 5897 21985
rect 5931 21951 5989 21985
rect 6023 21951 6043 21985
rect 4948 21942 6043 21951
rect 6095 21942 6107 21951
rect 6159 21942 6171 21994
rect 6223 21942 6235 21994
rect 6287 21985 6299 21994
rect 6287 21942 6299 21951
rect 6351 21985 9861 21994
rect 6351 21951 6357 21985
rect 6391 21951 6449 21985
rect 6483 21951 6541 21985
rect 6575 21951 6633 21985
rect 6667 21951 6725 21985
rect 6759 21951 6817 21985
rect 6851 21951 6909 21985
rect 6943 21951 7001 21985
rect 7035 21951 7093 21985
rect 7127 21951 7185 21985
rect 7219 21951 7277 21985
rect 7311 21951 7369 21985
rect 7403 21951 7461 21985
rect 7495 21951 7553 21985
rect 7587 21951 7645 21985
rect 7679 21951 7737 21985
rect 7771 21951 7829 21985
rect 7863 21951 7921 21985
rect 7955 21951 8013 21985
rect 8047 21951 8105 21985
rect 8139 21951 8197 21985
rect 8231 21951 8289 21985
rect 8323 21951 8381 21985
rect 8415 21951 8473 21985
rect 8507 21951 8565 21985
rect 8599 21951 8657 21985
rect 8691 21951 8749 21985
rect 8783 21951 8841 21985
rect 8875 21951 8933 21985
rect 8967 21951 9025 21985
rect 9059 21951 9117 21985
rect 9151 21951 9209 21985
rect 9243 21951 9301 21985
rect 9335 21951 9393 21985
rect 9427 21951 9485 21985
rect 9519 21951 9577 21985
rect 9611 21951 9669 21985
rect 9703 21951 9761 21985
rect 9795 21951 9853 21985
rect 6351 21942 9861 21951
rect 9913 21942 9925 21994
rect 9977 21985 9989 21994
rect 10041 21985 10053 21994
rect 9979 21951 9989 21985
rect 9977 21942 9989 21951
rect 10041 21942 10053 21951
rect 10105 21942 10117 21994
rect 10169 21985 13679 21994
rect 13731 21985 13743 21994
rect 10169 21951 10221 21985
rect 10255 21951 10313 21985
rect 10347 21951 10405 21985
rect 10439 21951 10497 21985
rect 10531 21951 10589 21985
rect 10623 21951 10681 21985
rect 10715 21951 10773 21985
rect 10807 21951 10865 21985
rect 10899 21951 10957 21985
rect 10991 21951 11049 21985
rect 11083 21951 11141 21985
rect 11175 21951 11233 21985
rect 11267 21951 11325 21985
rect 11359 21951 11417 21985
rect 11451 21951 11509 21985
rect 11543 21951 11601 21985
rect 11635 21951 11693 21985
rect 11727 21951 11785 21985
rect 11819 21951 11877 21985
rect 11911 21951 11969 21985
rect 12003 21951 12061 21985
rect 12095 21951 12153 21985
rect 12187 21951 12245 21985
rect 12279 21951 12337 21985
rect 12371 21951 12429 21985
rect 12463 21951 12521 21985
rect 12555 21951 12613 21985
rect 12647 21951 12705 21985
rect 12739 21951 12797 21985
rect 12831 21951 12889 21985
rect 12923 21951 12981 21985
rect 13015 21951 13073 21985
rect 13107 21951 13165 21985
rect 13199 21951 13257 21985
rect 13291 21951 13349 21985
rect 13383 21951 13441 21985
rect 13475 21951 13533 21985
rect 13567 21951 13625 21985
rect 13659 21951 13679 21985
rect 10169 21942 13679 21951
rect 13731 21942 13743 21951
rect 13795 21942 13807 21994
rect 13859 21942 13871 21994
rect 13923 21985 13935 21994
rect 13923 21942 13935 21951
rect 13987 21985 17497 21994
rect 13987 21951 13993 21985
rect 14027 21951 14085 21985
rect 14119 21951 14177 21985
rect 14211 21951 14269 21985
rect 14303 21951 14361 21985
rect 14395 21951 14453 21985
rect 14487 21951 14545 21985
rect 14579 21951 14637 21985
rect 14671 21951 14729 21985
rect 14763 21951 14821 21985
rect 14855 21951 14913 21985
rect 14947 21951 15005 21985
rect 15039 21951 15097 21985
rect 15131 21951 15189 21985
rect 15223 21951 15281 21985
rect 15315 21951 15373 21985
rect 15407 21951 15465 21985
rect 15499 21951 15557 21985
rect 15591 21951 15649 21985
rect 15683 21951 15741 21985
rect 15775 21951 15833 21985
rect 15867 21951 15925 21985
rect 15959 21951 16017 21985
rect 16051 21951 16109 21985
rect 16143 21951 16201 21985
rect 16235 21951 16293 21985
rect 16327 21951 16385 21985
rect 16419 21951 16477 21985
rect 16511 21951 16569 21985
rect 16603 21951 16661 21985
rect 16695 21951 16753 21985
rect 16787 21951 16845 21985
rect 16879 21951 16937 21985
rect 16971 21951 17029 21985
rect 17063 21951 17121 21985
rect 17155 21951 17213 21985
rect 17247 21951 17305 21985
rect 17339 21951 17397 21985
rect 17431 21951 17489 21985
rect 13987 21942 17497 21951
rect 17549 21942 17561 21994
rect 17613 21985 17625 21994
rect 17677 21985 17689 21994
rect 17615 21951 17625 21985
rect 17613 21942 17625 21951
rect 17677 21942 17689 21951
rect 17741 21942 17753 21994
rect 17805 21985 20220 21994
rect 17805 21951 17857 21985
rect 17891 21951 17949 21985
rect 17983 21951 18041 21985
rect 18075 21951 18133 21985
rect 18167 21951 18225 21985
rect 18259 21951 18317 21985
rect 18351 21951 18409 21985
rect 18443 21951 18501 21985
rect 18535 21951 18593 21985
rect 18627 21951 18685 21985
rect 18719 21951 18777 21985
rect 18811 21951 18869 21985
rect 18903 21951 18961 21985
rect 18995 21951 19053 21985
rect 19087 21951 19145 21985
rect 19179 21951 19237 21985
rect 19271 21951 19329 21985
rect 19363 21951 19421 21985
rect 19455 21951 19513 21985
rect 19547 21951 19605 21985
rect 19639 21951 19697 21985
rect 19731 21951 19789 21985
rect 19823 21951 19881 21985
rect 19915 21951 19973 21985
rect 20007 21951 20065 21985
rect 20099 21951 20157 21985
rect 20191 21951 20220 21985
rect 17805 21942 20220 21951
rect 4948 21920 20220 21942
rect 4948 21450 20220 21472
rect 4948 21441 6703 21450
rect 6755 21441 6767 21450
rect 6819 21441 6831 21450
rect 4948 21407 4977 21441
rect 5011 21407 5069 21441
rect 5103 21407 5161 21441
rect 5195 21407 5253 21441
rect 5287 21407 5345 21441
rect 5379 21407 5437 21441
rect 5471 21407 5529 21441
rect 5563 21407 5621 21441
rect 5655 21407 5713 21441
rect 5747 21407 5805 21441
rect 5839 21407 5897 21441
rect 5931 21407 5989 21441
rect 6023 21407 6081 21441
rect 6115 21407 6173 21441
rect 6207 21407 6265 21441
rect 6299 21407 6357 21441
rect 6391 21407 6449 21441
rect 6483 21407 6541 21441
rect 6575 21407 6633 21441
rect 6667 21407 6703 21441
rect 6759 21407 6767 21441
rect 4948 21398 6703 21407
rect 6755 21398 6767 21407
rect 6819 21398 6831 21407
rect 6883 21398 6895 21450
rect 6947 21398 6959 21450
rect 7011 21441 10521 21450
rect 7035 21407 7093 21441
rect 7127 21407 7185 21441
rect 7219 21407 7277 21441
rect 7311 21407 7369 21441
rect 7403 21407 7461 21441
rect 7495 21407 7553 21441
rect 7587 21407 7645 21441
rect 7679 21407 7737 21441
rect 7771 21407 7829 21441
rect 7863 21407 7921 21441
rect 7955 21407 8013 21441
rect 8047 21407 8105 21441
rect 8139 21407 8197 21441
rect 8231 21407 8289 21441
rect 8323 21407 8381 21441
rect 8415 21407 8473 21441
rect 8507 21407 8565 21441
rect 8599 21407 8657 21441
rect 8691 21407 8749 21441
rect 8783 21407 8841 21441
rect 8875 21407 8933 21441
rect 8967 21407 9025 21441
rect 9059 21407 9117 21441
rect 9151 21407 9209 21441
rect 9243 21407 9301 21441
rect 9335 21407 9393 21441
rect 9427 21407 9485 21441
rect 9519 21407 9577 21441
rect 9611 21407 9669 21441
rect 9703 21407 9761 21441
rect 9795 21407 9853 21441
rect 9887 21407 9945 21441
rect 9979 21407 10037 21441
rect 10071 21407 10129 21441
rect 10163 21407 10221 21441
rect 10255 21407 10313 21441
rect 10347 21407 10405 21441
rect 10439 21407 10497 21441
rect 7011 21398 10521 21407
rect 10573 21398 10585 21450
rect 10637 21398 10649 21450
rect 10701 21441 10713 21450
rect 10765 21441 10777 21450
rect 10829 21441 14339 21450
rect 14391 21441 14403 21450
rect 14455 21441 14467 21450
rect 10765 21407 10773 21441
rect 10829 21407 10865 21441
rect 10899 21407 10957 21441
rect 10991 21407 11049 21441
rect 11083 21407 11141 21441
rect 11175 21407 11233 21441
rect 11267 21407 11325 21441
rect 11359 21407 11417 21441
rect 11451 21407 11509 21441
rect 11543 21407 11601 21441
rect 11635 21407 11693 21441
rect 11727 21407 11785 21441
rect 11819 21407 11877 21441
rect 11911 21407 11969 21441
rect 12003 21407 12061 21441
rect 12095 21407 12153 21441
rect 12187 21407 12245 21441
rect 12279 21407 12337 21441
rect 12371 21407 12429 21441
rect 12463 21407 12521 21441
rect 12555 21407 12613 21441
rect 12647 21407 12705 21441
rect 12739 21407 12797 21441
rect 12831 21407 12889 21441
rect 12923 21407 12981 21441
rect 13015 21407 13073 21441
rect 13107 21407 13165 21441
rect 13199 21407 13257 21441
rect 13291 21407 13349 21441
rect 13383 21407 13441 21441
rect 13475 21407 13533 21441
rect 13567 21407 13625 21441
rect 13659 21407 13717 21441
rect 13751 21407 13809 21441
rect 13843 21407 13901 21441
rect 13935 21407 13993 21441
rect 14027 21407 14085 21441
rect 14119 21407 14177 21441
rect 14211 21407 14269 21441
rect 14303 21407 14339 21441
rect 14395 21407 14403 21441
rect 10701 21398 10713 21407
rect 10765 21398 10777 21407
rect 10829 21398 14339 21407
rect 14391 21398 14403 21407
rect 14455 21398 14467 21407
rect 14519 21398 14531 21450
rect 14583 21398 14595 21450
rect 14647 21441 18157 21450
rect 14671 21407 14729 21441
rect 14763 21407 14821 21441
rect 14855 21407 14913 21441
rect 14947 21407 15005 21441
rect 15039 21407 15097 21441
rect 15131 21407 15189 21441
rect 15223 21407 15281 21441
rect 15315 21407 15373 21441
rect 15407 21407 15465 21441
rect 15499 21407 15557 21441
rect 15591 21407 15649 21441
rect 15683 21407 15741 21441
rect 15775 21407 15833 21441
rect 15867 21407 15925 21441
rect 15959 21407 16017 21441
rect 16051 21407 16109 21441
rect 16143 21407 16201 21441
rect 16235 21407 16293 21441
rect 16327 21407 16385 21441
rect 16419 21407 16477 21441
rect 16511 21407 16569 21441
rect 16603 21407 16661 21441
rect 16695 21407 16753 21441
rect 16787 21407 16845 21441
rect 16879 21407 16937 21441
rect 16971 21407 17029 21441
rect 17063 21407 17121 21441
rect 17155 21407 17213 21441
rect 17247 21407 17305 21441
rect 17339 21407 17397 21441
rect 17431 21407 17489 21441
rect 17523 21407 17581 21441
rect 17615 21407 17673 21441
rect 17707 21407 17765 21441
rect 17799 21407 17857 21441
rect 17891 21407 17949 21441
rect 17983 21407 18041 21441
rect 18075 21407 18133 21441
rect 14647 21398 18157 21407
rect 18209 21398 18221 21450
rect 18273 21398 18285 21450
rect 18337 21441 18349 21450
rect 18401 21441 18413 21450
rect 18465 21441 20220 21450
rect 18401 21407 18409 21441
rect 18465 21407 18501 21441
rect 18535 21407 18593 21441
rect 18627 21407 18685 21441
rect 18719 21407 18777 21441
rect 18811 21407 18869 21441
rect 18903 21407 18961 21441
rect 18995 21407 19053 21441
rect 19087 21407 19145 21441
rect 19179 21407 19237 21441
rect 19271 21407 19329 21441
rect 19363 21407 19421 21441
rect 19455 21407 19513 21441
rect 19547 21407 19605 21441
rect 19639 21407 19697 21441
rect 19731 21407 19789 21441
rect 19823 21407 19881 21441
rect 19915 21407 19973 21441
rect 20007 21407 20065 21441
rect 20099 21407 20157 21441
rect 20191 21407 20220 21441
rect 18337 21398 18349 21407
rect 18401 21398 18413 21407
rect 18465 21398 20220 21407
rect 4948 21376 20220 21398
rect 4948 20906 20220 20928
rect 4948 20897 6043 20906
rect 6095 20897 6107 20906
rect 4948 20863 4977 20897
rect 5011 20863 5069 20897
rect 5103 20863 5161 20897
rect 5195 20863 5253 20897
rect 5287 20863 5345 20897
rect 5379 20863 5437 20897
rect 5471 20863 5529 20897
rect 5563 20863 5621 20897
rect 5655 20863 5713 20897
rect 5747 20863 5805 20897
rect 5839 20863 5897 20897
rect 5931 20863 5989 20897
rect 6023 20863 6043 20897
rect 4948 20854 6043 20863
rect 6095 20854 6107 20863
rect 6159 20854 6171 20906
rect 6223 20854 6235 20906
rect 6287 20897 6299 20906
rect 6287 20854 6299 20863
rect 6351 20897 9861 20906
rect 6351 20863 6357 20897
rect 6391 20863 6449 20897
rect 6483 20863 6541 20897
rect 6575 20863 6633 20897
rect 6667 20863 6725 20897
rect 6759 20863 6817 20897
rect 6851 20863 6909 20897
rect 6943 20863 7001 20897
rect 7035 20863 7093 20897
rect 7127 20863 7185 20897
rect 7219 20863 7277 20897
rect 7311 20863 7369 20897
rect 7403 20863 7461 20897
rect 7495 20863 7553 20897
rect 7587 20863 7645 20897
rect 7679 20863 7737 20897
rect 7771 20863 7829 20897
rect 7863 20863 7921 20897
rect 7955 20863 8013 20897
rect 8047 20863 8105 20897
rect 8139 20863 8197 20897
rect 8231 20863 8289 20897
rect 8323 20863 8381 20897
rect 8415 20863 8473 20897
rect 8507 20863 8565 20897
rect 8599 20863 8657 20897
rect 8691 20863 8749 20897
rect 8783 20863 8841 20897
rect 8875 20863 8933 20897
rect 8967 20863 9025 20897
rect 9059 20863 9117 20897
rect 9151 20863 9209 20897
rect 9243 20863 9301 20897
rect 9335 20863 9393 20897
rect 9427 20863 9485 20897
rect 9519 20863 9577 20897
rect 9611 20863 9669 20897
rect 9703 20863 9761 20897
rect 9795 20863 9853 20897
rect 6351 20854 9861 20863
rect 9913 20854 9925 20906
rect 9977 20897 9989 20906
rect 10041 20897 10053 20906
rect 9979 20863 9989 20897
rect 9977 20854 9989 20863
rect 10041 20854 10053 20863
rect 10105 20854 10117 20906
rect 10169 20897 13679 20906
rect 13731 20897 13743 20906
rect 10169 20863 10221 20897
rect 10255 20863 10313 20897
rect 10347 20863 10405 20897
rect 10439 20863 10497 20897
rect 10531 20863 10589 20897
rect 10623 20863 10681 20897
rect 10715 20863 10773 20897
rect 10807 20863 10865 20897
rect 10899 20863 10957 20897
rect 10991 20863 11049 20897
rect 11083 20863 11141 20897
rect 11175 20863 11233 20897
rect 11267 20863 11325 20897
rect 11359 20863 11417 20897
rect 11451 20863 11509 20897
rect 11543 20863 11601 20897
rect 11635 20863 11693 20897
rect 11727 20863 11785 20897
rect 11819 20863 11877 20897
rect 11911 20863 11969 20897
rect 12003 20863 12061 20897
rect 12095 20863 12153 20897
rect 12187 20863 12245 20897
rect 12279 20863 12337 20897
rect 12371 20863 12429 20897
rect 12463 20863 12521 20897
rect 12555 20863 12613 20897
rect 12647 20863 12705 20897
rect 12739 20863 12797 20897
rect 12831 20863 12889 20897
rect 12923 20863 12981 20897
rect 13015 20863 13073 20897
rect 13107 20863 13165 20897
rect 13199 20863 13257 20897
rect 13291 20863 13349 20897
rect 13383 20863 13441 20897
rect 13475 20863 13533 20897
rect 13567 20863 13625 20897
rect 13659 20863 13679 20897
rect 10169 20854 13679 20863
rect 13731 20854 13743 20863
rect 13795 20854 13807 20906
rect 13859 20854 13871 20906
rect 13923 20897 13935 20906
rect 13923 20854 13935 20863
rect 13987 20897 17497 20906
rect 13987 20863 13993 20897
rect 14027 20863 14085 20897
rect 14119 20863 14177 20897
rect 14211 20863 14269 20897
rect 14303 20863 14361 20897
rect 14395 20863 14453 20897
rect 14487 20863 14545 20897
rect 14579 20863 14637 20897
rect 14671 20863 14729 20897
rect 14763 20863 14821 20897
rect 14855 20863 14913 20897
rect 14947 20863 15005 20897
rect 15039 20863 15097 20897
rect 15131 20863 15189 20897
rect 15223 20863 15281 20897
rect 15315 20863 15373 20897
rect 15407 20863 15465 20897
rect 15499 20863 15557 20897
rect 15591 20863 15649 20897
rect 15683 20863 15741 20897
rect 15775 20863 15833 20897
rect 15867 20863 15925 20897
rect 15959 20863 16017 20897
rect 16051 20863 16109 20897
rect 16143 20863 16201 20897
rect 16235 20863 16293 20897
rect 16327 20863 16385 20897
rect 16419 20863 16477 20897
rect 16511 20863 16569 20897
rect 16603 20863 16661 20897
rect 16695 20863 16753 20897
rect 16787 20863 16845 20897
rect 16879 20863 16937 20897
rect 16971 20863 17029 20897
rect 17063 20863 17121 20897
rect 17155 20863 17213 20897
rect 17247 20863 17305 20897
rect 17339 20863 17397 20897
rect 17431 20863 17489 20897
rect 13987 20854 17497 20863
rect 17549 20854 17561 20906
rect 17613 20897 17625 20906
rect 17677 20897 17689 20906
rect 17615 20863 17625 20897
rect 17613 20854 17625 20863
rect 17677 20854 17689 20863
rect 17741 20854 17753 20906
rect 17805 20897 20220 20906
rect 17805 20863 17857 20897
rect 17891 20863 17949 20897
rect 17983 20863 18041 20897
rect 18075 20863 18133 20897
rect 18167 20863 18225 20897
rect 18259 20863 18317 20897
rect 18351 20863 18409 20897
rect 18443 20863 18501 20897
rect 18535 20863 18593 20897
rect 18627 20863 18685 20897
rect 18719 20863 18777 20897
rect 18811 20863 18869 20897
rect 18903 20863 18961 20897
rect 18995 20863 19053 20897
rect 19087 20863 19145 20897
rect 19179 20863 19237 20897
rect 19271 20863 19329 20897
rect 19363 20863 19421 20897
rect 19455 20863 19513 20897
rect 19547 20863 19605 20897
rect 19639 20863 19697 20897
rect 19731 20863 19789 20897
rect 19823 20863 19881 20897
rect 19915 20863 19973 20897
rect 20007 20863 20065 20897
rect 20099 20863 20157 20897
rect 20191 20863 20220 20897
rect 17805 20854 20220 20863
rect 4948 20832 20220 20854
rect 4948 20362 20220 20384
rect 4948 20353 6703 20362
rect 6755 20353 6767 20362
rect 6819 20353 6831 20362
rect 4948 20319 4977 20353
rect 5011 20319 5069 20353
rect 5103 20319 5161 20353
rect 5195 20319 5253 20353
rect 5287 20319 5345 20353
rect 5379 20319 5437 20353
rect 5471 20319 5529 20353
rect 5563 20319 5621 20353
rect 5655 20319 5713 20353
rect 5747 20319 5805 20353
rect 5839 20319 5897 20353
rect 5931 20319 5989 20353
rect 6023 20319 6081 20353
rect 6115 20319 6173 20353
rect 6207 20319 6265 20353
rect 6299 20319 6357 20353
rect 6391 20319 6449 20353
rect 6483 20319 6541 20353
rect 6575 20319 6633 20353
rect 6667 20319 6703 20353
rect 6759 20319 6767 20353
rect 4948 20310 6703 20319
rect 6755 20310 6767 20319
rect 6819 20310 6831 20319
rect 6883 20310 6895 20362
rect 6947 20310 6959 20362
rect 7011 20353 10521 20362
rect 7035 20319 7093 20353
rect 7127 20319 7185 20353
rect 7219 20319 7277 20353
rect 7311 20319 7369 20353
rect 7403 20319 7461 20353
rect 7495 20319 7553 20353
rect 7587 20319 7645 20353
rect 7679 20319 7737 20353
rect 7771 20319 7829 20353
rect 7863 20319 7921 20353
rect 7955 20319 8013 20353
rect 8047 20319 8105 20353
rect 8139 20319 8197 20353
rect 8231 20319 8289 20353
rect 8323 20319 8381 20353
rect 8415 20319 8473 20353
rect 8507 20319 8565 20353
rect 8599 20319 8657 20353
rect 8691 20319 8749 20353
rect 8783 20319 8841 20353
rect 8875 20319 8933 20353
rect 8967 20319 9025 20353
rect 9059 20319 9117 20353
rect 9151 20319 9209 20353
rect 9243 20319 9301 20353
rect 9335 20319 9393 20353
rect 9427 20319 9485 20353
rect 9519 20319 9577 20353
rect 9611 20319 9669 20353
rect 9703 20319 9761 20353
rect 9795 20319 9853 20353
rect 9887 20319 9945 20353
rect 9979 20319 10037 20353
rect 10071 20319 10129 20353
rect 10163 20319 10221 20353
rect 10255 20319 10313 20353
rect 10347 20319 10405 20353
rect 10439 20319 10497 20353
rect 7011 20310 10521 20319
rect 10573 20310 10585 20362
rect 10637 20310 10649 20362
rect 10701 20353 10713 20362
rect 10765 20353 10777 20362
rect 10829 20353 14339 20362
rect 14391 20353 14403 20362
rect 14455 20353 14467 20362
rect 10765 20319 10773 20353
rect 10829 20319 10865 20353
rect 10899 20319 10957 20353
rect 10991 20319 11049 20353
rect 11083 20319 11141 20353
rect 11175 20319 11233 20353
rect 11267 20319 11325 20353
rect 11359 20319 11417 20353
rect 11451 20319 11509 20353
rect 11543 20319 11601 20353
rect 11635 20319 11693 20353
rect 11727 20319 11785 20353
rect 11819 20319 11877 20353
rect 11911 20319 11969 20353
rect 12003 20319 12061 20353
rect 12095 20319 12153 20353
rect 12187 20319 12245 20353
rect 12279 20319 12337 20353
rect 12371 20319 12429 20353
rect 12463 20319 12521 20353
rect 12555 20319 12613 20353
rect 12647 20319 12705 20353
rect 12739 20319 12797 20353
rect 12831 20319 12889 20353
rect 12923 20319 12981 20353
rect 13015 20319 13073 20353
rect 13107 20319 13165 20353
rect 13199 20319 13257 20353
rect 13291 20319 13349 20353
rect 13383 20319 13441 20353
rect 13475 20319 13533 20353
rect 13567 20319 13625 20353
rect 13659 20319 13717 20353
rect 13751 20319 13809 20353
rect 13843 20319 13901 20353
rect 13935 20319 13993 20353
rect 14027 20319 14085 20353
rect 14119 20319 14177 20353
rect 14211 20319 14269 20353
rect 14303 20319 14339 20353
rect 14395 20319 14403 20353
rect 10701 20310 10713 20319
rect 10765 20310 10777 20319
rect 10829 20310 14339 20319
rect 14391 20310 14403 20319
rect 14455 20310 14467 20319
rect 14519 20310 14531 20362
rect 14583 20310 14595 20362
rect 14647 20353 18157 20362
rect 14671 20319 14729 20353
rect 14763 20319 14821 20353
rect 14855 20319 14913 20353
rect 14947 20319 15005 20353
rect 15039 20319 15097 20353
rect 15131 20319 15189 20353
rect 15223 20319 15281 20353
rect 15315 20319 15373 20353
rect 15407 20319 15465 20353
rect 15499 20319 15557 20353
rect 15591 20319 15649 20353
rect 15683 20319 15741 20353
rect 15775 20319 15833 20353
rect 15867 20319 15925 20353
rect 15959 20319 16017 20353
rect 16051 20319 16109 20353
rect 16143 20319 16201 20353
rect 16235 20319 16293 20353
rect 16327 20319 16385 20353
rect 16419 20319 16477 20353
rect 16511 20319 16569 20353
rect 16603 20319 16661 20353
rect 16695 20319 16753 20353
rect 16787 20319 16845 20353
rect 16879 20319 16937 20353
rect 16971 20319 17029 20353
rect 17063 20319 17121 20353
rect 17155 20319 17213 20353
rect 17247 20319 17305 20353
rect 17339 20319 17397 20353
rect 17431 20319 17489 20353
rect 17523 20319 17581 20353
rect 17615 20319 17673 20353
rect 17707 20319 17765 20353
rect 17799 20319 17857 20353
rect 17891 20319 17949 20353
rect 17983 20319 18041 20353
rect 18075 20319 18133 20353
rect 14647 20310 18157 20319
rect 18209 20310 18221 20362
rect 18273 20310 18285 20362
rect 18337 20353 18349 20362
rect 18401 20353 18413 20362
rect 18465 20353 20220 20362
rect 18401 20319 18409 20353
rect 18465 20319 18501 20353
rect 18535 20319 18593 20353
rect 18627 20319 18685 20353
rect 18719 20319 18777 20353
rect 18811 20319 18869 20353
rect 18903 20319 18961 20353
rect 18995 20319 19053 20353
rect 19087 20319 19145 20353
rect 19179 20319 19237 20353
rect 19271 20319 19329 20353
rect 19363 20319 19421 20353
rect 19455 20319 19513 20353
rect 19547 20319 19605 20353
rect 19639 20319 19697 20353
rect 19731 20319 19789 20353
rect 19823 20319 19881 20353
rect 19915 20319 19973 20353
rect 20007 20319 20065 20353
rect 20099 20319 20157 20353
rect 20191 20319 20220 20353
rect 18337 20310 18349 20319
rect 18401 20310 18413 20319
rect 18465 20310 20220 20319
rect 4948 20288 20220 20310
rect -200 19840 0 19880
rect -200 19750 290 19840
rect 320 19818 20220 19840
rect 320 19809 6043 19818
rect 6095 19809 6107 19818
rect 320 19775 4977 19809
rect 5011 19775 5069 19809
rect 5103 19775 5161 19809
rect 5195 19775 5253 19809
rect 5287 19775 5345 19809
rect 5379 19775 5437 19809
rect 5471 19775 5529 19809
rect 5563 19775 5621 19809
rect 5655 19775 5713 19809
rect 5747 19775 5805 19809
rect 5839 19775 5897 19809
rect 5931 19775 5989 19809
rect 6023 19775 6043 19809
rect 320 19766 6043 19775
rect 6095 19766 6107 19775
rect 6159 19766 6171 19818
rect 6223 19766 6235 19818
rect 6287 19809 6299 19818
rect 6287 19766 6299 19775
rect 6351 19809 9861 19818
rect 6351 19775 6357 19809
rect 6391 19775 6449 19809
rect 6483 19775 6541 19809
rect 6575 19775 6633 19809
rect 6667 19775 6725 19809
rect 6759 19775 6817 19809
rect 6851 19775 6909 19809
rect 6943 19775 7001 19809
rect 7035 19775 7093 19809
rect 7127 19775 7185 19809
rect 7219 19775 7277 19809
rect 7311 19775 7369 19809
rect 7403 19775 7461 19809
rect 7495 19775 7553 19809
rect 7587 19775 7645 19809
rect 7679 19775 7737 19809
rect 7771 19775 7829 19809
rect 7863 19775 7921 19809
rect 7955 19775 8013 19809
rect 8047 19775 8105 19809
rect 8139 19775 8197 19809
rect 8231 19775 8289 19809
rect 8323 19775 8381 19809
rect 8415 19775 8473 19809
rect 8507 19775 8565 19809
rect 8599 19775 8657 19809
rect 8691 19775 8749 19809
rect 8783 19775 8841 19809
rect 8875 19775 8933 19809
rect 8967 19775 9025 19809
rect 9059 19775 9117 19809
rect 9151 19775 9209 19809
rect 9243 19775 9301 19809
rect 9335 19775 9393 19809
rect 9427 19775 9485 19809
rect 9519 19775 9577 19809
rect 9611 19775 9669 19809
rect 9703 19775 9761 19809
rect 9795 19775 9853 19809
rect 6351 19766 9861 19775
rect 9913 19766 9925 19818
rect 9977 19809 9989 19818
rect 10041 19809 10053 19818
rect 9979 19775 9989 19809
rect 9977 19766 9989 19775
rect 10041 19766 10053 19775
rect 10105 19766 10117 19818
rect 10169 19809 13679 19818
rect 13731 19809 13743 19818
rect 10169 19775 10221 19809
rect 10255 19775 10313 19809
rect 10347 19775 10405 19809
rect 10439 19775 10497 19809
rect 10531 19775 10589 19809
rect 10623 19775 10681 19809
rect 10715 19775 10773 19809
rect 10807 19775 10865 19809
rect 10899 19775 10957 19809
rect 10991 19775 11049 19809
rect 11083 19775 11141 19809
rect 11175 19775 11233 19809
rect 11267 19775 11325 19809
rect 11359 19775 11417 19809
rect 11451 19775 11509 19809
rect 11543 19775 11601 19809
rect 11635 19775 11693 19809
rect 11727 19775 11785 19809
rect 11819 19775 11877 19809
rect 11911 19775 11969 19809
rect 12003 19775 12061 19809
rect 12095 19775 12153 19809
rect 12187 19775 12245 19809
rect 12279 19775 12337 19809
rect 12371 19775 12429 19809
rect 12463 19775 12521 19809
rect 12555 19775 12613 19809
rect 12647 19775 12705 19809
rect 12739 19775 12797 19809
rect 12831 19775 12889 19809
rect 12923 19775 12981 19809
rect 13015 19775 13073 19809
rect 13107 19775 13165 19809
rect 13199 19775 13257 19809
rect 13291 19775 13349 19809
rect 13383 19775 13441 19809
rect 13475 19775 13533 19809
rect 13567 19775 13625 19809
rect 13659 19775 13679 19809
rect 10169 19766 13679 19775
rect 13731 19766 13743 19775
rect 13795 19766 13807 19818
rect 13859 19766 13871 19818
rect 13923 19809 13935 19818
rect 13923 19766 13935 19775
rect 13987 19809 17497 19818
rect 13987 19775 13993 19809
rect 14027 19775 14085 19809
rect 14119 19775 14177 19809
rect 14211 19775 14269 19809
rect 14303 19775 14361 19809
rect 14395 19775 14453 19809
rect 14487 19775 14545 19809
rect 14579 19775 14637 19809
rect 14671 19775 14729 19809
rect 14763 19775 14821 19809
rect 14855 19775 14913 19809
rect 14947 19775 15005 19809
rect 15039 19775 15097 19809
rect 15131 19775 15189 19809
rect 15223 19775 15281 19809
rect 15315 19775 15373 19809
rect 15407 19775 15465 19809
rect 15499 19775 15557 19809
rect 15591 19775 15649 19809
rect 15683 19775 15741 19809
rect 15775 19775 15833 19809
rect 15867 19775 15925 19809
rect 15959 19775 16017 19809
rect 16051 19775 16109 19809
rect 16143 19775 16201 19809
rect 16235 19775 16293 19809
rect 16327 19775 16385 19809
rect 16419 19775 16477 19809
rect 16511 19775 16569 19809
rect 16603 19775 16661 19809
rect 16695 19775 16753 19809
rect 16787 19775 16845 19809
rect 16879 19775 16937 19809
rect 16971 19775 17029 19809
rect 17063 19775 17121 19809
rect 17155 19775 17213 19809
rect 17247 19775 17305 19809
rect 17339 19775 17397 19809
rect 17431 19775 17489 19809
rect 13987 19766 17497 19775
rect 17549 19766 17561 19818
rect 17613 19809 17625 19818
rect 17677 19809 17689 19818
rect 17615 19775 17625 19809
rect 17613 19766 17625 19775
rect 17677 19766 17689 19775
rect 17741 19766 17753 19818
rect 17805 19809 20220 19818
rect 17805 19775 17857 19809
rect 17891 19775 17949 19809
rect 17983 19775 18041 19809
rect 18075 19775 18133 19809
rect 18167 19775 18225 19809
rect 18259 19775 18317 19809
rect 18351 19775 18409 19809
rect 18443 19775 18501 19809
rect 18535 19775 18593 19809
rect 18627 19775 18685 19809
rect 18719 19775 18777 19809
rect 18811 19775 18869 19809
rect 18903 19775 18961 19809
rect 18995 19775 19053 19809
rect 19087 19775 19145 19809
rect 19179 19775 19237 19809
rect 19271 19775 19329 19809
rect 19363 19775 19421 19809
rect 19455 19775 19513 19809
rect 19547 19775 19605 19809
rect 19639 19775 19697 19809
rect 19731 19775 19789 19809
rect 19823 19775 19881 19809
rect 19915 19775 19973 19809
rect 20007 19775 20065 19809
rect 20099 19775 20157 19809
rect 20191 19775 20220 19809
rect 17805 19766 20220 19775
rect 320 19750 20220 19766
rect -200 19690 0 19750
rect 4948 19744 20220 19750
rect -200 19300 0 19360
rect -200 19296 4960 19300
rect -200 19274 20220 19296
rect -200 19265 6703 19274
rect 6755 19265 6767 19274
rect 6819 19265 6831 19274
rect -200 19231 4977 19265
rect 5011 19231 5069 19265
rect 5103 19231 5161 19265
rect 5195 19231 5253 19265
rect 5287 19231 5345 19265
rect 5379 19231 5437 19265
rect 5471 19231 5529 19265
rect 5563 19231 5621 19265
rect 5655 19231 5713 19265
rect 5747 19231 5805 19265
rect 5839 19231 5897 19265
rect 5931 19231 5989 19265
rect 6023 19231 6081 19265
rect 6115 19231 6173 19265
rect 6207 19231 6265 19265
rect 6299 19231 6357 19265
rect 6391 19231 6449 19265
rect 6483 19231 6541 19265
rect 6575 19231 6633 19265
rect 6667 19231 6703 19265
rect 6759 19231 6767 19265
rect -200 19222 6703 19231
rect 6755 19222 6767 19231
rect 6819 19222 6831 19231
rect 6883 19222 6895 19274
rect 6947 19222 6959 19274
rect 7011 19265 10521 19274
rect 7035 19231 7093 19265
rect 7127 19231 7185 19265
rect 7219 19231 7277 19265
rect 7311 19231 7369 19265
rect 7403 19231 7461 19265
rect 7495 19231 7553 19265
rect 7587 19231 7645 19265
rect 7679 19231 7737 19265
rect 7771 19231 7829 19265
rect 7863 19231 7921 19265
rect 7955 19231 8013 19265
rect 8047 19231 8105 19265
rect 8139 19231 8197 19265
rect 8231 19231 8289 19265
rect 8323 19231 8381 19265
rect 8415 19231 8473 19265
rect 8507 19231 8565 19265
rect 8599 19231 8657 19265
rect 8691 19231 8749 19265
rect 8783 19231 8841 19265
rect 8875 19231 8933 19265
rect 8967 19231 9025 19265
rect 9059 19231 9117 19265
rect 9151 19231 9209 19265
rect 9243 19231 9301 19265
rect 9335 19231 9393 19265
rect 9427 19231 9485 19265
rect 9519 19231 9577 19265
rect 9611 19231 9669 19265
rect 9703 19231 9761 19265
rect 9795 19231 9853 19265
rect 9887 19231 9945 19265
rect 9979 19231 10037 19265
rect 10071 19231 10129 19265
rect 10163 19231 10221 19265
rect 10255 19231 10313 19265
rect 10347 19231 10405 19265
rect 10439 19231 10497 19265
rect 7011 19222 10521 19231
rect 10573 19222 10585 19274
rect 10637 19222 10649 19274
rect 10701 19265 10713 19274
rect 10765 19265 10777 19274
rect 10829 19265 14339 19274
rect 14391 19265 14403 19274
rect 14455 19265 14467 19274
rect 10765 19231 10773 19265
rect 10829 19231 10865 19265
rect 10899 19231 10957 19265
rect 10991 19231 11049 19265
rect 11083 19231 11141 19265
rect 11175 19231 11233 19265
rect 11267 19231 11325 19265
rect 11359 19231 11417 19265
rect 11451 19231 11509 19265
rect 11543 19231 11601 19265
rect 11635 19231 11693 19265
rect 11727 19231 11785 19265
rect 11819 19231 11877 19265
rect 11911 19231 11969 19265
rect 12003 19231 12061 19265
rect 12095 19231 12153 19265
rect 12187 19231 12245 19265
rect 12279 19231 12337 19265
rect 12371 19231 12429 19265
rect 12463 19231 12521 19265
rect 12555 19231 12613 19265
rect 12647 19231 12705 19265
rect 12739 19231 12797 19265
rect 12831 19231 12889 19265
rect 12923 19231 12981 19265
rect 13015 19231 13073 19265
rect 13107 19231 13165 19265
rect 13199 19231 13257 19265
rect 13291 19231 13349 19265
rect 13383 19231 13441 19265
rect 13475 19231 13533 19265
rect 13567 19231 13625 19265
rect 13659 19231 13717 19265
rect 13751 19231 13809 19265
rect 13843 19231 13901 19265
rect 13935 19231 13993 19265
rect 14027 19231 14085 19265
rect 14119 19231 14177 19265
rect 14211 19231 14269 19265
rect 14303 19231 14339 19265
rect 14395 19231 14403 19265
rect 10701 19222 10713 19231
rect 10765 19222 10777 19231
rect 10829 19222 14339 19231
rect 14391 19222 14403 19231
rect 14455 19222 14467 19231
rect 14519 19222 14531 19274
rect 14583 19222 14595 19274
rect 14647 19265 18157 19274
rect 14671 19231 14729 19265
rect 14763 19231 14821 19265
rect 14855 19231 14913 19265
rect 14947 19231 15005 19265
rect 15039 19231 15097 19265
rect 15131 19231 15189 19265
rect 15223 19231 15281 19265
rect 15315 19231 15373 19265
rect 15407 19231 15465 19265
rect 15499 19231 15557 19265
rect 15591 19231 15649 19265
rect 15683 19231 15741 19265
rect 15775 19231 15833 19265
rect 15867 19231 15925 19265
rect 15959 19231 16017 19265
rect 16051 19231 16109 19265
rect 16143 19231 16201 19265
rect 16235 19231 16293 19265
rect 16327 19231 16385 19265
rect 16419 19231 16477 19265
rect 16511 19231 16569 19265
rect 16603 19231 16661 19265
rect 16695 19231 16753 19265
rect 16787 19231 16845 19265
rect 16879 19231 16937 19265
rect 16971 19231 17029 19265
rect 17063 19231 17121 19265
rect 17155 19231 17213 19265
rect 17247 19231 17305 19265
rect 17339 19231 17397 19265
rect 17431 19231 17489 19265
rect 17523 19231 17581 19265
rect 17615 19231 17673 19265
rect 17707 19231 17765 19265
rect 17799 19231 17857 19265
rect 17891 19231 17949 19265
rect 17983 19231 18041 19265
rect 18075 19231 18133 19265
rect 14647 19222 18157 19231
rect 18209 19222 18221 19274
rect 18273 19222 18285 19274
rect 18337 19265 18349 19274
rect 18401 19265 18413 19274
rect 18465 19265 20220 19274
rect 18401 19231 18409 19265
rect 18465 19231 18501 19265
rect 18535 19231 18593 19265
rect 18627 19231 18685 19265
rect 18719 19231 18777 19265
rect 18811 19231 18869 19265
rect 18903 19231 18961 19265
rect 18995 19231 19053 19265
rect 19087 19231 19145 19265
rect 19179 19231 19237 19265
rect 19271 19231 19329 19265
rect 19363 19231 19421 19265
rect 19455 19231 19513 19265
rect 19547 19231 19605 19265
rect 19639 19231 19697 19265
rect 19731 19231 19789 19265
rect 19823 19231 19881 19265
rect 19915 19231 19973 19265
rect 20007 19231 20065 19265
rect 20099 19231 20157 19265
rect 20191 19231 20220 19265
rect 18337 19222 18349 19231
rect 18401 19222 18413 19231
rect 18465 19222 20220 19231
rect -200 19200 20220 19222
rect -200 19170 0 19200
rect 4948 18730 20220 18752
rect 4948 18721 6043 18730
rect 6095 18721 6107 18730
rect 4948 18687 4977 18721
rect 5011 18687 5069 18721
rect 5103 18687 5161 18721
rect 5195 18687 5253 18721
rect 5287 18687 5345 18721
rect 5379 18687 5437 18721
rect 5471 18687 5529 18721
rect 5563 18687 5621 18721
rect 5655 18687 5713 18721
rect 5747 18687 5805 18721
rect 5839 18687 5897 18721
rect 5931 18687 5989 18721
rect 6023 18687 6043 18721
rect 4948 18678 6043 18687
rect 6095 18678 6107 18687
rect 6159 18678 6171 18730
rect 6223 18678 6235 18730
rect 6287 18721 6299 18730
rect 6287 18678 6299 18687
rect 6351 18721 9861 18730
rect 6351 18687 6357 18721
rect 6391 18687 6449 18721
rect 6483 18687 6541 18721
rect 6575 18687 6633 18721
rect 6667 18687 6725 18721
rect 6759 18687 6817 18721
rect 6851 18687 6909 18721
rect 6943 18687 7001 18721
rect 7035 18687 7093 18721
rect 7127 18687 7185 18721
rect 7219 18687 7277 18721
rect 7311 18687 7369 18721
rect 7403 18687 7461 18721
rect 7495 18687 7553 18721
rect 7587 18687 7645 18721
rect 7679 18687 7737 18721
rect 7771 18687 7829 18721
rect 7863 18687 7921 18721
rect 7955 18687 8013 18721
rect 8047 18687 8105 18721
rect 8139 18687 8197 18721
rect 8231 18687 8289 18721
rect 8323 18687 8381 18721
rect 8415 18687 8473 18721
rect 8507 18687 8565 18721
rect 8599 18687 8657 18721
rect 8691 18687 8749 18721
rect 8783 18687 8841 18721
rect 8875 18687 8933 18721
rect 8967 18687 9025 18721
rect 9059 18687 9117 18721
rect 9151 18687 9209 18721
rect 9243 18687 9301 18721
rect 9335 18687 9393 18721
rect 9427 18687 9485 18721
rect 9519 18687 9577 18721
rect 9611 18687 9669 18721
rect 9703 18687 9761 18721
rect 9795 18687 9853 18721
rect 6351 18678 9861 18687
rect 9913 18678 9925 18730
rect 9977 18721 9989 18730
rect 10041 18721 10053 18730
rect 9979 18687 9989 18721
rect 9977 18678 9989 18687
rect 10041 18678 10053 18687
rect 10105 18678 10117 18730
rect 10169 18721 13679 18730
rect 13731 18721 13743 18730
rect 10169 18687 10221 18721
rect 10255 18687 10313 18721
rect 10347 18687 10405 18721
rect 10439 18687 10497 18721
rect 10531 18687 10589 18721
rect 10623 18687 10681 18721
rect 10715 18687 10773 18721
rect 10807 18687 10865 18721
rect 10899 18687 10957 18721
rect 10991 18687 11049 18721
rect 11083 18687 11141 18721
rect 11175 18687 11233 18721
rect 11267 18687 11325 18721
rect 11359 18687 11417 18721
rect 11451 18687 11509 18721
rect 11543 18687 11601 18721
rect 11635 18687 11693 18721
rect 11727 18687 11785 18721
rect 11819 18687 11877 18721
rect 11911 18687 11969 18721
rect 12003 18687 12061 18721
rect 12095 18687 12153 18721
rect 12187 18687 12245 18721
rect 12279 18687 12337 18721
rect 12371 18687 12429 18721
rect 12463 18687 12521 18721
rect 12555 18687 12613 18721
rect 12647 18687 12705 18721
rect 12739 18687 12797 18721
rect 12831 18687 12889 18721
rect 12923 18687 12981 18721
rect 13015 18687 13073 18721
rect 13107 18687 13165 18721
rect 13199 18687 13257 18721
rect 13291 18687 13349 18721
rect 13383 18687 13441 18721
rect 13475 18687 13533 18721
rect 13567 18687 13625 18721
rect 13659 18687 13679 18721
rect 10169 18678 13679 18687
rect 13731 18678 13743 18687
rect 13795 18678 13807 18730
rect 13859 18678 13871 18730
rect 13923 18721 13935 18730
rect 13923 18678 13935 18687
rect 13987 18721 17497 18730
rect 13987 18687 13993 18721
rect 14027 18687 14085 18721
rect 14119 18687 14177 18721
rect 14211 18687 14269 18721
rect 14303 18687 14361 18721
rect 14395 18687 14453 18721
rect 14487 18687 14545 18721
rect 14579 18687 14637 18721
rect 14671 18687 14729 18721
rect 14763 18687 14821 18721
rect 14855 18687 14913 18721
rect 14947 18687 15005 18721
rect 15039 18687 15097 18721
rect 15131 18687 15189 18721
rect 15223 18687 15281 18721
rect 15315 18687 15373 18721
rect 15407 18687 15465 18721
rect 15499 18687 15557 18721
rect 15591 18687 15649 18721
rect 15683 18687 15741 18721
rect 15775 18687 15833 18721
rect 15867 18687 15925 18721
rect 15959 18687 16017 18721
rect 16051 18687 16109 18721
rect 16143 18687 16201 18721
rect 16235 18687 16293 18721
rect 16327 18687 16385 18721
rect 16419 18687 16477 18721
rect 16511 18687 16569 18721
rect 16603 18687 16661 18721
rect 16695 18687 16753 18721
rect 16787 18687 16845 18721
rect 16879 18687 16937 18721
rect 16971 18687 17029 18721
rect 17063 18687 17121 18721
rect 17155 18687 17213 18721
rect 17247 18687 17305 18721
rect 17339 18687 17397 18721
rect 17431 18687 17489 18721
rect 13987 18678 17497 18687
rect 17549 18678 17561 18730
rect 17613 18721 17625 18730
rect 17677 18721 17689 18730
rect 17615 18687 17625 18721
rect 17613 18678 17625 18687
rect 17677 18678 17689 18687
rect 17741 18678 17753 18730
rect 17805 18721 20220 18730
rect 17805 18687 17857 18721
rect 17891 18687 17949 18721
rect 17983 18687 18041 18721
rect 18075 18687 18133 18721
rect 18167 18687 18225 18721
rect 18259 18687 18317 18721
rect 18351 18687 18409 18721
rect 18443 18687 18501 18721
rect 18535 18687 18593 18721
rect 18627 18687 18685 18721
rect 18719 18687 18777 18721
rect 18811 18687 18869 18721
rect 18903 18687 18961 18721
rect 18995 18687 19053 18721
rect 19087 18687 19145 18721
rect 19179 18687 19237 18721
rect 19271 18687 19329 18721
rect 19363 18687 19421 18721
rect 19455 18687 19513 18721
rect 19547 18687 19605 18721
rect 19639 18687 19697 18721
rect 19731 18687 19789 18721
rect 19823 18687 19881 18721
rect 19915 18687 19973 18721
rect 20007 18687 20065 18721
rect 20099 18687 20157 18721
rect 20191 18687 20220 18721
rect 17805 18678 20220 18687
rect 4948 18656 20220 18678
rect 4948 18186 20220 18208
rect 4948 18177 6703 18186
rect 6755 18177 6767 18186
rect 6819 18177 6831 18186
rect 4948 18143 4977 18177
rect 5011 18143 5069 18177
rect 5103 18143 5161 18177
rect 5195 18143 5253 18177
rect 5287 18143 5345 18177
rect 5379 18143 5437 18177
rect 5471 18143 5529 18177
rect 5563 18143 5621 18177
rect 5655 18143 5713 18177
rect 5747 18143 5805 18177
rect 5839 18143 5897 18177
rect 5931 18143 5989 18177
rect 6023 18143 6081 18177
rect 6115 18143 6173 18177
rect 6207 18143 6265 18177
rect 6299 18143 6357 18177
rect 6391 18143 6449 18177
rect 6483 18143 6541 18177
rect 6575 18143 6633 18177
rect 6667 18143 6703 18177
rect 6759 18143 6767 18177
rect 4948 18134 6703 18143
rect 6755 18134 6767 18143
rect 6819 18134 6831 18143
rect 6883 18134 6895 18186
rect 6947 18134 6959 18186
rect 7011 18177 10521 18186
rect 7035 18143 7093 18177
rect 7127 18143 7185 18177
rect 7219 18143 7277 18177
rect 7311 18143 7369 18177
rect 7403 18143 7461 18177
rect 7495 18143 7553 18177
rect 7587 18143 7645 18177
rect 7679 18143 7737 18177
rect 7771 18143 7829 18177
rect 7863 18143 7921 18177
rect 7955 18143 8013 18177
rect 8047 18143 8105 18177
rect 8139 18143 8197 18177
rect 8231 18143 8289 18177
rect 8323 18143 8381 18177
rect 8415 18143 8473 18177
rect 8507 18143 8565 18177
rect 8599 18143 8657 18177
rect 8691 18143 8749 18177
rect 8783 18143 8841 18177
rect 8875 18143 8933 18177
rect 8967 18143 9025 18177
rect 9059 18143 9117 18177
rect 9151 18143 9209 18177
rect 9243 18143 9301 18177
rect 9335 18143 9393 18177
rect 9427 18143 9485 18177
rect 9519 18143 9577 18177
rect 9611 18143 9669 18177
rect 9703 18143 9761 18177
rect 9795 18143 9853 18177
rect 9887 18143 9945 18177
rect 9979 18143 10037 18177
rect 10071 18143 10129 18177
rect 10163 18143 10221 18177
rect 10255 18143 10313 18177
rect 10347 18143 10405 18177
rect 10439 18143 10497 18177
rect 7011 18134 10521 18143
rect 10573 18134 10585 18186
rect 10637 18134 10649 18186
rect 10701 18177 10713 18186
rect 10765 18177 10777 18186
rect 10829 18177 14339 18186
rect 14391 18177 14403 18186
rect 14455 18177 14467 18186
rect 10765 18143 10773 18177
rect 10829 18143 10865 18177
rect 10899 18143 10957 18177
rect 10991 18143 11049 18177
rect 11083 18143 11141 18177
rect 11175 18143 11233 18177
rect 11267 18143 11325 18177
rect 11359 18143 11417 18177
rect 11451 18143 11509 18177
rect 11543 18143 11601 18177
rect 11635 18143 11693 18177
rect 11727 18143 11785 18177
rect 11819 18143 11877 18177
rect 11911 18143 11969 18177
rect 12003 18143 12061 18177
rect 12095 18143 12153 18177
rect 12187 18143 12245 18177
rect 12279 18143 12337 18177
rect 12371 18143 12429 18177
rect 12463 18143 12521 18177
rect 12555 18143 12613 18177
rect 12647 18143 12705 18177
rect 12739 18143 12797 18177
rect 12831 18143 12889 18177
rect 12923 18143 12981 18177
rect 13015 18143 13073 18177
rect 13107 18143 13165 18177
rect 13199 18143 13257 18177
rect 13291 18143 13349 18177
rect 13383 18143 13441 18177
rect 13475 18143 13533 18177
rect 13567 18143 13625 18177
rect 13659 18143 13717 18177
rect 13751 18143 13809 18177
rect 13843 18143 13901 18177
rect 13935 18143 13993 18177
rect 14027 18143 14085 18177
rect 14119 18143 14177 18177
rect 14211 18143 14269 18177
rect 14303 18143 14339 18177
rect 14395 18143 14403 18177
rect 10701 18134 10713 18143
rect 10765 18134 10777 18143
rect 10829 18134 14339 18143
rect 14391 18134 14403 18143
rect 14455 18134 14467 18143
rect 14519 18134 14531 18186
rect 14583 18134 14595 18186
rect 14647 18177 18157 18186
rect 14671 18143 14729 18177
rect 14763 18143 14821 18177
rect 14855 18143 14913 18177
rect 14947 18143 15005 18177
rect 15039 18143 15097 18177
rect 15131 18143 15189 18177
rect 15223 18143 15281 18177
rect 15315 18143 15373 18177
rect 15407 18143 15465 18177
rect 15499 18143 15557 18177
rect 15591 18143 15649 18177
rect 15683 18143 15741 18177
rect 15775 18143 15833 18177
rect 15867 18143 15925 18177
rect 15959 18143 16017 18177
rect 16051 18143 16109 18177
rect 16143 18143 16201 18177
rect 16235 18143 16293 18177
rect 16327 18143 16385 18177
rect 16419 18143 16477 18177
rect 16511 18143 16569 18177
rect 16603 18143 16661 18177
rect 16695 18143 16753 18177
rect 16787 18143 16845 18177
rect 16879 18143 16937 18177
rect 16971 18143 17029 18177
rect 17063 18143 17121 18177
rect 17155 18143 17213 18177
rect 17247 18143 17305 18177
rect 17339 18143 17397 18177
rect 17431 18143 17489 18177
rect 17523 18143 17581 18177
rect 17615 18143 17673 18177
rect 17707 18143 17765 18177
rect 17799 18143 17857 18177
rect 17891 18143 17949 18177
rect 17983 18143 18041 18177
rect 18075 18143 18133 18177
rect 14647 18134 18157 18143
rect 18209 18134 18221 18186
rect 18273 18134 18285 18186
rect 18337 18177 18349 18186
rect 18401 18177 18413 18186
rect 18465 18177 20220 18186
rect 18401 18143 18409 18177
rect 18465 18143 18501 18177
rect 18535 18143 18593 18177
rect 18627 18143 18685 18177
rect 18719 18143 18777 18177
rect 18811 18143 18869 18177
rect 18903 18143 18961 18177
rect 18995 18143 19053 18177
rect 19087 18143 19145 18177
rect 19179 18143 19237 18177
rect 19271 18143 19329 18177
rect 19363 18143 19421 18177
rect 19455 18143 19513 18177
rect 19547 18143 19605 18177
rect 19639 18143 19697 18177
rect 19731 18143 19789 18177
rect 19823 18143 19881 18177
rect 19915 18143 19973 18177
rect 20007 18143 20065 18177
rect 20099 18143 20157 18177
rect 20191 18143 20220 18177
rect 18337 18134 18349 18143
rect 18401 18134 18413 18143
rect 18465 18134 20220 18143
rect 4948 18112 20220 18134
rect 4948 17642 20220 17664
rect 4948 17633 6043 17642
rect 6095 17633 6107 17642
rect 4948 17599 4977 17633
rect 5011 17599 5069 17633
rect 5103 17599 5161 17633
rect 5195 17599 5253 17633
rect 5287 17599 5345 17633
rect 5379 17599 5437 17633
rect 5471 17599 5529 17633
rect 5563 17599 5621 17633
rect 5655 17599 5713 17633
rect 5747 17599 5805 17633
rect 5839 17599 5897 17633
rect 5931 17599 5989 17633
rect 6023 17599 6043 17633
rect 4948 17590 6043 17599
rect 6095 17590 6107 17599
rect 6159 17590 6171 17642
rect 6223 17590 6235 17642
rect 6287 17633 6299 17642
rect 6287 17590 6299 17599
rect 6351 17633 9861 17642
rect 6351 17599 6357 17633
rect 6391 17599 6449 17633
rect 6483 17599 6541 17633
rect 6575 17599 6633 17633
rect 6667 17599 6725 17633
rect 6759 17599 6817 17633
rect 6851 17599 6909 17633
rect 6943 17599 7001 17633
rect 7035 17599 7093 17633
rect 7127 17599 7185 17633
rect 7219 17599 7277 17633
rect 7311 17599 7369 17633
rect 7403 17599 7461 17633
rect 7495 17599 7553 17633
rect 7587 17599 7645 17633
rect 7679 17599 7737 17633
rect 7771 17599 7829 17633
rect 7863 17599 7921 17633
rect 7955 17599 8013 17633
rect 8047 17599 8105 17633
rect 8139 17599 8197 17633
rect 8231 17599 8289 17633
rect 8323 17599 8381 17633
rect 8415 17599 8473 17633
rect 8507 17599 8565 17633
rect 8599 17599 8657 17633
rect 8691 17599 8749 17633
rect 8783 17599 8841 17633
rect 8875 17599 8933 17633
rect 8967 17599 9025 17633
rect 9059 17599 9117 17633
rect 9151 17599 9209 17633
rect 9243 17599 9301 17633
rect 9335 17599 9393 17633
rect 9427 17599 9485 17633
rect 9519 17599 9577 17633
rect 9611 17599 9669 17633
rect 9703 17599 9761 17633
rect 9795 17599 9853 17633
rect 6351 17590 9861 17599
rect 9913 17590 9925 17642
rect 9977 17633 9989 17642
rect 10041 17633 10053 17642
rect 9979 17599 9989 17633
rect 9977 17590 9989 17599
rect 10041 17590 10053 17599
rect 10105 17590 10117 17642
rect 10169 17633 13679 17642
rect 13731 17633 13743 17642
rect 10169 17599 10221 17633
rect 10255 17599 10313 17633
rect 10347 17599 10405 17633
rect 10439 17599 10497 17633
rect 10531 17599 10589 17633
rect 10623 17599 10681 17633
rect 10715 17599 10773 17633
rect 10807 17599 10865 17633
rect 10899 17599 10957 17633
rect 10991 17599 11049 17633
rect 11083 17599 11141 17633
rect 11175 17599 11233 17633
rect 11267 17599 11325 17633
rect 11359 17599 11417 17633
rect 11451 17599 11509 17633
rect 11543 17599 11601 17633
rect 11635 17599 11693 17633
rect 11727 17599 11785 17633
rect 11819 17599 11877 17633
rect 11911 17599 11969 17633
rect 12003 17599 12061 17633
rect 12095 17599 12153 17633
rect 12187 17599 12245 17633
rect 12279 17599 12337 17633
rect 12371 17599 12429 17633
rect 12463 17599 12521 17633
rect 12555 17599 12613 17633
rect 12647 17599 12705 17633
rect 12739 17599 12797 17633
rect 12831 17599 12889 17633
rect 12923 17599 12981 17633
rect 13015 17599 13073 17633
rect 13107 17599 13165 17633
rect 13199 17599 13257 17633
rect 13291 17599 13349 17633
rect 13383 17599 13441 17633
rect 13475 17599 13533 17633
rect 13567 17599 13625 17633
rect 13659 17599 13679 17633
rect 10169 17590 13679 17599
rect 13731 17590 13743 17599
rect 13795 17590 13807 17642
rect 13859 17590 13871 17642
rect 13923 17633 13935 17642
rect 13923 17590 13935 17599
rect 13987 17633 17497 17642
rect 13987 17599 13993 17633
rect 14027 17599 14085 17633
rect 14119 17599 14177 17633
rect 14211 17599 14269 17633
rect 14303 17599 14361 17633
rect 14395 17599 14453 17633
rect 14487 17599 14545 17633
rect 14579 17599 14637 17633
rect 14671 17599 14729 17633
rect 14763 17599 14821 17633
rect 14855 17599 14913 17633
rect 14947 17599 15005 17633
rect 15039 17599 15097 17633
rect 15131 17599 15189 17633
rect 15223 17599 15281 17633
rect 15315 17599 15373 17633
rect 15407 17599 15465 17633
rect 15499 17599 15557 17633
rect 15591 17599 15649 17633
rect 15683 17599 15741 17633
rect 15775 17599 15833 17633
rect 15867 17599 15925 17633
rect 15959 17599 16017 17633
rect 16051 17599 16109 17633
rect 16143 17599 16201 17633
rect 16235 17599 16293 17633
rect 16327 17599 16385 17633
rect 16419 17599 16477 17633
rect 16511 17599 16569 17633
rect 16603 17599 16661 17633
rect 16695 17599 16753 17633
rect 16787 17599 16845 17633
rect 16879 17599 16937 17633
rect 16971 17599 17029 17633
rect 17063 17599 17121 17633
rect 17155 17599 17213 17633
rect 17247 17599 17305 17633
rect 17339 17599 17397 17633
rect 17431 17599 17489 17633
rect 13987 17590 17497 17599
rect 17549 17590 17561 17642
rect 17613 17633 17625 17642
rect 17677 17633 17689 17642
rect 17615 17599 17625 17633
rect 17613 17590 17625 17599
rect 17677 17590 17689 17599
rect 17741 17590 17753 17642
rect 17805 17633 20220 17642
rect 17805 17599 17857 17633
rect 17891 17599 17949 17633
rect 17983 17599 18041 17633
rect 18075 17599 18133 17633
rect 18167 17599 18225 17633
rect 18259 17599 18317 17633
rect 18351 17599 18409 17633
rect 18443 17599 18501 17633
rect 18535 17599 18593 17633
rect 18627 17599 18685 17633
rect 18719 17599 18777 17633
rect 18811 17599 18869 17633
rect 18903 17599 18961 17633
rect 18995 17599 19053 17633
rect 19087 17599 19145 17633
rect 19179 17599 19237 17633
rect 19271 17599 19329 17633
rect 19363 17599 19421 17633
rect 19455 17599 19513 17633
rect 19547 17599 19605 17633
rect 19639 17599 19697 17633
rect 19731 17599 19789 17633
rect 19823 17599 19881 17633
rect 19915 17599 19973 17633
rect 20007 17599 20065 17633
rect 20099 17599 20157 17633
rect 20191 17599 20220 17633
rect 17805 17590 20220 17599
rect 4948 17568 20220 17590
rect 4948 17098 20220 17120
rect 4948 17089 6703 17098
rect 6755 17089 6767 17098
rect 6819 17089 6831 17098
rect 4948 17055 4977 17089
rect 5011 17055 5069 17089
rect 5103 17055 5161 17089
rect 5195 17055 5253 17089
rect 5287 17055 5345 17089
rect 5379 17055 5437 17089
rect 5471 17055 5529 17089
rect 5563 17055 5621 17089
rect 5655 17055 5713 17089
rect 5747 17055 5805 17089
rect 5839 17055 5897 17089
rect 5931 17055 5989 17089
rect 6023 17055 6081 17089
rect 6115 17055 6173 17089
rect 6207 17055 6265 17089
rect 6299 17055 6357 17089
rect 6391 17055 6449 17089
rect 6483 17055 6541 17089
rect 6575 17055 6633 17089
rect 6667 17055 6703 17089
rect 6759 17055 6767 17089
rect 4948 17046 6703 17055
rect 6755 17046 6767 17055
rect 6819 17046 6831 17055
rect 6883 17046 6895 17098
rect 6947 17046 6959 17098
rect 7011 17089 10521 17098
rect 7035 17055 7093 17089
rect 7127 17055 7185 17089
rect 7219 17055 7277 17089
rect 7311 17055 7369 17089
rect 7403 17055 7461 17089
rect 7495 17055 7553 17089
rect 7587 17055 7645 17089
rect 7679 17055 7737 17089
rect 7771 17055 7829 17089
rect 7863 17055 7921 17089
rect 7955 17055 8013 17089
rect 8047 17055 8105 17089
rect 8139 17055 8197 17089
rect 8231 17055 8289 17089
rect 8323 17055 8381 17089
rect 8415 17055 8473 17089
rect 8507 17055 8565 17089
rect 8599 17055 8657 17089
rect 8691 17055 8749 17089
rect 8783 17055 8841 17089
rect 8875 17055 8933 17089
rect 8967 17055 9025 17089
rect 9059 17055 9117 17089
rect 9151 17055 9209 17089
rect 9243 17055 9301 17089
rect 9335 17055 9393 17089
rect 9427 17055 9485 17089
rect 9519 17055 9577 17089
rect 9611 17055 9669 17089
rect 9703 17055 9761 17089
rect 9795 17055 9853 17089
rect 9887 17055 9945 17089
rect 9979 17055 10037 17089
rect 10071 17055 10129 17089
rect 10163 17055 10221 17089
rect 10255 17055 10313 17089
rect 10347 17055 10405 17089
rect 10439 17055 10497 17089
rect 7011 17046 10521 17055
rect 10573 17046 10585 17098
rect 10637 17046 10649 17098
rect 10701 17089 10713 17098
rect 10765 17089 10777 17098
rect 10829 17089 14339 17098
rect 14391 17089 14403 17098
rect 14455 17089 14467 17098
rect 10765 17055 10773 17089
rect 10829 17055 10865 17089
rect 10899 17055 10957 17089
rect 10991 17055 11049 17089
rect 11083 17055 11141 17089
rect 11175 17055 11233 17089
rect 11267 17055 11325 17089
rect 11359 17055 11417 17089
rect 11451 17055 11509 17089
rect 11543 17055 11601 17089
rect 11635 17055 11693 17089
rect 11727 17055 11785 17089
rect 11819 17055 11877 17089
rect 11911 17055 11969 17089
rect 12003 17055 12061 17089
rect 12095 17055 12153 17089
rect 12187 17055 12245 17089
rect 12279 17055 12337 17089
rect 12371 17055 12429 17089
rect 12463 17055 12521 17089
rect 12555 17055 12613 17089
rect 12647 17055 12705 17089
rect 12739 17055 12797 17089
rect 12831 17055 12889 17089
rect 12923 17055 12981 17089
rect 13015 17055 13073 17089
rect 13107 17055 13165 17089
rect 13199 17055 13257 17089
rect 13291 17055 13349 17089
rect 13383 17055 13441 17089
rect 13475 17055 13533 17089
rect 13567 17055 13625 17089
rect 13659 17055 13717 17089
rect 13751 17055 13809 17089
rect 13843 17055 13901 17089
rect 13935 17055 13993 17089
rect 14027 17055 14085 17089
rect 14119 17055 14177 17089
rect 14211 17055 14269 17089
rect 14303 17055 14339 17089
rect 14395 17055 14403 17089
rect 10701 17046 10713 17055
rect 10765 17046 10777 17055
rect 10829 17046 14339 17055
rect 14391 17046 14403 17055
rect 14455 17046 14467 17055
rect 14519 17046 14531 17098
rect 14583 17046 14595 17098
rect 14647 17089 18157 17098
rect 14671 17055 14729 17089
rect 14763 17055 14821 17089
rect 14855 17055 14913 17089
rect 14947 17055 15005 17089
rect 15039 17055 15097 17089
rect 15131 17055 15189 17089
rect 15223 17055 15281 17089
rect 15315 17055 15373 17089
rect 15407 17055 15465 17089
rect 15499 17055 15557 17089
rect 15591 17055 15649 17089
rect 15683 17055 15741 17089
rect 15775 17055 15833 17089
rect 15867 17055 15925 17089
rect 15959 17055 16017 17089
rect 16051 17055 16109 17089
rect 16143 17055 16201 17089
rect 16235 17055 16293 17089
rect 16327 17055 16385 17089
rect 16419 17055 16477 17089
rect 16511 17055 16569 17089
rect 16603 17055 16661 17089
rect 16695 17055 16753 17089
rect 16787 17055 16845 17089
rect 16879 17055 16937 17089
rect 16971 17055 17029 17089
rect 17063 17055 17121 17089
rect 17155 17055 17213 17089
rect 17247 17055 17305 17089
rect 17339 17055 17397 17089
rect 17431 17055 17489 17089
rect 17523 17055 17581 17089
rect 17615 17055 17673 17089
rect 17707 17055 17765 17089
rect 17799 17055 17857 17089
rect 17891 17055 17949 17089
rect 17983 17055 18041 17089
rect 18075 17055 18133 17089
rect 14647 17046 18157 17055
rect 18209 17046 18221 17098
rect 18273 17046 18285 17098
rect 18337 17089 18349 17098
rect 18401 17089 18413 17098
rect 18465 17089 20220 17098
rect 18401 17055 18409 17089
rect 18465 17055 18501 17089
rect 18535 17055 18593 17089
rect 18627 17055 18685 17089
rect 18719 17055 18777 17089
rect 18811 17055 18869 17089
rect 18903 17055 18961 17089
rect 18995 17055 19053 17089
rect 19087 17055 19145 17089
rect 19179 17055 19237 17089
rect 19271 17055 19329 17089
rect 19363 17055 19421 17089
rect 19455 17055 19513 17089
rect 19547 17055 19605 17089
rect 19639 17055 19697 17089
rect 19731 17055 19789 17089
rect 19823 17055 19881 17089
rect 19915 17055 19973 17089
rect 20007 17055 20065 17089
rect 20099 17055 20157 17089
rect 20191 17055 20220 17089
rect 18337 17046 18349 17055
rect 18401 17046 18413 17055
rect 18465 17046 20220 17055
rect 4948 17024 20220 17046
rect 4948 16554 20220 16576
rect 4948 16545 6043 16554
rect 6095 16545 6107 16554
rect 4948 16511 4977 16545
rect 5011 16511 5069 16545
rect 5103 16511 5161 16545
rect 5195 16511 5253 16545
rect 5287 16511 5345 16545
rect 5379 16511 5437 16545
rect 5471 16511 5529 16545
rect 5563 16511 5621 16545
rect 5655 16511 5713 16545
rect 5747 16511 5805 16545
rect 5839 16511 5897 16545
rect 5931 16511 5989 16545
rect 6023 16511 6043 16545
rect 4948 16502 6043 16511
rect 6095 16502 6107 16511
rect 6159 16502 6171 16554
rect 6223 16502 6235 16554
rect 6287 16545 6299 16554
rect 6287 16502 6299 16511
rect 6351 16545 9861 16554
rect 6351 16511 6357 16545
rect 6391 16511 6449 16545
rect 6483 16511 6541 16545
rect 6575 16511 6633 16545
rect 6667 16511 6725 16545
rect 6759 16511 6817 16545
rect 6851 16511 6909 16545
rect 6943 16511 7001 16545
rect 7035 16511 7093 16545
rect 7127 16511 7185 16545
rect 7219 16511 7277 16545
rect 7311 16511 7369 16545
rect 7403 16511 7461 16545
rect 7495 16511 7553 16545
rect 7587 16511 7645 16545
rect 7679 16511 7737 16545
rect 7771 16511 7829 16545
rect 7863 16511 7921 16545
rect 7955 16511 8013 16545
rect 8047 16511 8105 16545
rect 8139 16511 8197 16545
rect 8231 16511 8289 16545
rect 8323 16511 8381 16545
rect 8415 16511 8473 16545
rect 8507 16511 8565 16545
rect 8599 16511 8657 16545
rect 8691 16511 8749 16545
rect 8783 16511 8841 16545
rect 8875 16511 8933 16545
rect 8967 16511 9025 16545
rect 9059 16511 9117 16545
rect 9151 16511 9209 16545
rect 9243 16511 9301 16545
rect 9335 16511 9393 16545
rect 9427 16511 9485 16545
rect 9519 16511 9577 16545
rect 9611 16511 9669 16545
rect 9703 16511 9761 16545
rect 9795 16511 9853 16545
rect 6351 16502 9861 16511
rect 9913 16502 9925 16554
rect 9977 16545 9989 16554
rect 10041 16545 10053 16554
rect 9979 16511 9989 16545
rect 9977 16502 9989 16511
rect 10041 16502 10053 16511
rect 10105 16502 10117 16554
rect 10169 16545 13679 16554
rect 13731 16545 13743 16554
rect 10169 16511 10221 16545
rect 10255 16511 10313 16545
rect 10347 16511 10405 16545
rect 10439 16511 10497 16545
rect 10531 16511 10589 16545
rect 10623 16511 10681 16545
rect 10715 16511 10773 16545
rect 10807 16511 10865 16545
rect 10899 16511 10957 16545
rect 10991 16511 11049 16545
rect 11083 16511 11141 16545
rect 11175 16511 11233 16545
rect 11267 16511 11325 16545
rect 11359 16511 11417 16545
rect 11451 16511 11509 16545
rect 11543 16511 11601 16545
rect 11635 16511 11693 16545
rect 11727 16511 11785 16545
rect 11819 16511 11877 16545
rect 11911 16511 11969 16545
rect 12003 16511 12061 16545
rect 12095 16511 12153 16545
rect 12187 16511 12245 16545
rect 12279 16511 12337 16545
rect 12371 16511 12429 16545
rect 12463 16511 12521 16545
rect 12555 16511 12613 16545
rect 12647 16511 12705 16545
rect 12739 16511 12797 16545
rect 12831 16511 12889 16545
rect 12923 16511 12981 16545
rect 13015 16511 13073 16545
rect 13107 16511 13165 16545
rect 13199 16511 13257 16545
rect 13291 16511 13349 16545
rect 13383 16511 13441 16545
rect 13475 16511 13533 16545
rect 13567 16511 13625 16545
rect 13659 16511 13679 16545
rect 10169 16502 13679 16511
rect 13731 16502 13743 16511
rect 13795 16502 13807 16554
rect 13859 16502 13871 16554
rect 13923 16545 13935 16554
rect 13923 16502 13935 16511
rect 13987 16545 17497 16554
rect 13987 16511 13993 16545
rect 14027 16511 14085 16545
rect 14119 16511 14177 16545
rect 14211 16511 14269 16545
rect 14303 16511 14361 16545
rect 14395 16511 14453 16545
rect 14487 16511 14545 16545
rect 14579 16511 14637 16545
rect 14671 16511 14729 16545
rect 14763 16511 14821 16545
rect 14855 16511 14913 16545
rect 14947 16511 15005 16545
rect 15039 16511 15097 16545
rect 15131 16511 15189 16545
rect 15223 16511 15281 16545
rect 15315 16511 15373 16545
rect 15407 16511 15465 16545
rect 15499 16511 15557 16545
rect 15591 16511 15649 16545
rect 15683 16511 15741 16545
rect 15775 16511 15833 16545
rect 15867 16511 15925 16545
rect 15959 16511 16017 16545
rect 16051 16511 16109 16545
rect 16143 16511 16201 16545
rect 16235 16511 16293 16545
rect 16327 16511 16385 16545
rect 16419 16511 16477 16545
rect 16511 16511 16569 16545
rect 16603 16511 16661 16545
rect 16695 16511 16753 16545
rect 16787 16511 16845 16545
rect 16879 16511 16937 16545
rect 16971 16511 17029 16545
rect 17063 16511 17121 16545
rect 17155 16511 17213 16545
rect 17247 16511 17305 16545
rect 17339 16511 17397 16545
rect 17431 16511 17489 16545
rect 13987 16502 17497 16511
rect 17549 16502 17561 16554
rect 17613 16545 17625 16554
rect 17677 16545 17689 16554
rect 17615 16511 17625 16545
rect 17613 16502 17625 16511
rect 17677 16502 17689 16511
rect 17741 16502 17753 16554
rect 17805 16545 20220 16554
rect 17805 16511 17857 16545
rect 17891 16511 17949 16545
rect 17983 16511 18041 16545
rect 18075 16511 18133 16545
rect 18167 16511 18225 16545
rect 18259 16511 18317 16545
rect 18351 16511 18409 16545
rect 18443 16511 18501 16545
rect 18535 16511 18593 16545
rect 18627 16511 18685 16545
rect 18719 16511 18777 16545
rect 18811 16511 18869 16545
rect 18903 16511 18961 16545
rect 18995 16511 19053 16545
rect 19087 16511 19145 16545
rect 19179 16511 19237 16545
rect 19271 16511 19329 16545
rect 19363 16511 19421 16545
rect 19455 16511 19513 16545
rect 19547 16511 19605 16545
rect 19639 16511 19697 16545
rect 19731 16511 19789 16545
rect 19823 16511 19881 16545
rect 19915 16511 19973 16545
rect 20007 16511 20065 16545
rect 20099 16511 20157 16545
rect 20191 16511 20220 16545
rect 17805 16502 20220 16511
rect 4948 16480 20220 16502
rect 4948 16010 20220 16032
rect 4948 16001 6703 16010
rect 6755 16001 6767 16010
rect 6819 16001 6831 16010
rect 4948 15967 4977 16001
rect 5011 15967 5069 16001
rect 5103 15967 5161 16001
rect 5195 15967 5253 16001
rect 5287 15967 5345 16001
rect 5379 15967 5437 16001
rect 5471 15967 5529 16001
rect 5563 15967 5621 16001
rect 5655 15967 5713 16001
rect 5747 15967 5805 16001
rect 5839 15967 5897 16001
rect 5931 15967 5989 16001
rect 6023 15967 6081 16001
rect 6115 15967 6173 16001
rect 6207 15967 6265 16001
rect 6299 15967 6357 16001
rect 6391 15967 6449 16001
rect 6483 15967 6541 16001
rect 6575 15967 6633 16001
rect 6667 15967 6703 16001
rect 6759 15967 6767 16001
rect 4948 15958 6703 15967
rect 6755 15958 6767 15967
rect 6819 15958 6831 15967
rect 6883 15958 6895 16010
rect 6947 15958 6959 16010
rect 7011 16001 10521 16010
rect 7035 15967 7093 16001
rect 7127 15967 7185 16001
rect 7219 15967 7277 16001
rect 7311 15967 7369 16001
rect 7403 15967 7461 16001
rect 7495 15967 7553 16001
rect 7587 15967 7645 16001
rect 7679 15967 7737 16001
rect 7771 15967 7829 16001
rect 7863 15967 7921 16001
rect 7955 15967 8013 16001
rect 8047 15967 8105 16001
rect 8139 15967 8197 16001
rect 8231 15967 8289 16001
rect 8323 15967 8381 16001
rect 8415 15967 8473 16001
rect 8507 15967 8565 16001
rect 8599 15967 8657 16001
rect 8691 15967 8749 16001
rect 8783 15967 8841 16001
rect 8875 15967 8933 16001
rect 8967 15967 9025 16001
rect 9059 15967 9117 16001
rect 9151 15967 9209 16001
rect 9243 15967 9301 16001
rect 9335 15967 9393 16001
rect 9427 15967 9485 16001
rect 9519 15967 9577 16001
rect 9611 15967 9669 16001
rect 9703 15967 9761 16001
rect 9795 15967 9853 16001
rect 9887 15967 9945 16001
rect 9979 15967 10037 16001
rect 10071 15967 10129 16001
rect 10163 15967 10221 16001
rect 10255 15967 10313 16001
rect 10347 15967 10405 16001
rect 10439 15967 10497 16001
rect 7011 15958 10521 15967
rect 10573 15958 10585 16010
rect 10637 15958 10649 16010
rect 10701 16001 10713 16010
rect 10765 16001 10777 16010
rect 10829 16001 14339 16010
rect 14391 16001 14403 16010
rect 14455 16001 14467 16010
rect 10765 15967 10773 16001
rect 10829 15967 10865 16001
rect 10899 15967 10957 16001
rect 10991 15967 11049 16001
rect 11083 15967 11141 16001
rect 11175 15967 11233 16001
rect 11267 15967 11325 16001
rect 11359 15967 11417 16001
rect 11451 15967 11509 16001
rect 11543 15967 11601 16001
rect 11635 15967 11693 16001
rect 11727 15967 11785 16001
rect 11819 15967 11877 16001
rect 11911 15967 11969 16001
rect 12003 15967 12061 16001
rect 12095 15967 12153 16001
rect 12187 15967 12245 16001
rect 12279 15967 12337 16001
rect 12371 15967 12429 16001
rect 12463 15967 12521 16001
rect 12555 15967 12613 16001
rect 12647 15967 12705 16001
rect 12739 15967 12797 16001
rect 12831 15967 12889 16001
rect 12923 15967 12981 16001
rect 13015 15967 13073 16001
rect 13107 15967 13165 16001
rect 13199 15967 13257 16001
rect 13291 15967 13349 16001
rect 13383 15967 13441 16001
rect 13475 15967 13533 16001
rect 13567 15967 13625 16001
rect 13659 15967 13717 16001
rect 13751 15967 13809 16001
rect 13843 15967 13901 16001
rect 13935 15967 13993 16001
rect 14027 15967 14085 16001
rect 14119 15967 14177 16001
rect 14211 15967 14269 16001
rect 14303 15967 14339 16001
rect 14395 15967 14403 16001
rect 10701 15958 10713 15967
rect 10765 15958 10777 15967
rect 10829 15958 14339 15967
rect 14391 15958 14403 15967
rect 14455 15958 14467 15967
rect 14519 15958 14531 16010
rect 14583 15958 14595 16010
rect 14647 16001 18157 16010
rect 14671 15967 14729 16001
rect 14763 15967 14821 16001
rect 14855 15967 14913 16001
rect 14947 15967 15005 16001
rect 15039 15967 15097 16001
rect 15131 15967 15189 16001
rect 15223 15967 15281 16001
rect 15315 15967 15373 16001
rect 15407 15967 15465 16001
rect 15499 15967 15557 16001
rect 15591 15967 15649 16001
rect 15683 15967 15741 16001
rect 15775 15967 15833 16001
rect 15867 15967 15925 16001
rect 15959 15967 16017 16001
rect 16051 15967 16109 16001
rect 16143 15967 16201 16001
rect 16235 15967 16293 16001
rect 16327 15967 16385 16001
rect 16419 15967 16477 16001
rect 16511 15967 16569 16001
rect 16603 15967 16661 16001
rect 16695 15967 16753 16001
rect 16787 15967 16845 16001
rect 16879 15967 16937 16001
rect 16971 15967 17029 16001
rect 17063 15967 17121 16001
rect 17155 15967 17213 16001
rect 17247 15967 17305 16001
rect 17339 15967 17397 16001
rect 17431 15967 17489 16001
rect 17523 15967 17581 16001
rect 17615 15967 17673 16001
rect 17707 15967 17765 16001
rect 17799 15967 17857 16001
rect 17891 15967 17949 16001
rect 17983 15967 18041 16001
rect 18075 15967 18133 16001
rect 14647 15958 18157 15967
rect 18209 15958 18221 16010
rect 18273 15958 18285 16010
rect 18337 16001 18349 16010
rect 18401 16001 18413 16010
rect 18465 16001 20220 16010
rect 18401 15967 18409 16001
rect 18465 15967 18501 16001
rect 18535 15967 18593 16001
rect 18627 15967 18685 16001
rect 18719 15967 18777 16001
rect 18811 15967 18869 16001
rect 18903 15967 18961 16001
rect 18995 15967 19053 16001
rect 19087 15967 19145 16001
rect 19179 15967 19237 16001
rect 19271 15967 19329 16001
rect 19363 15967 19421 16001
rect 19455 15967 19513 16001
rect 19547 15967 19605 16001
rect 19639 15967 19697 16001
rect 19731 15967 19789 16001
rect 19823 15967 19881 16001
rect 19915 15967 19973 16001
rect 20007 15967 20065 16001
rect 20099 15967 20157 16001
rect 20191 15967 20220 16001
rect 18337 15958 18349 15967
rect 18401 15958 18413 15967
rect 18465 15958 20220 15967
rect 4948 15936 20220 15958
rect 4948 15466 20220 15488
rect 4948 15457 6043 15466
rect 6095 15457 6107 15466
rect 4948 15423 4977 15457
rect 5011 15423 5069 15457
rect 5103 15423 5161 15457
rect 5195 15423 5253 15457
rect 5287 15423 5345 15457
rect 5379 15423 5437 15457
rect 5471 15423 5529 15457
rect 5563 15423 5621 15457
rect 5655 15423 5713 15457
rect 5747 15423 5805 15457
rect 5839 15423 5897 15457
rect 5931 15423 5989 15457
rect 6023 15423 6043 15457
rect 4948 15414 6043 15423
rect 6095 15414 6107 15423
rect 6159 15414 6171 15466
rect 6223 15414 6235 15466
rect 6287 15457 6299 15466
rect 6287 15414 6299 15423
rect 6351 15457 9861 15466
rect 6351 15423 6357 15457
rect 6391 15423 6449 15457
rect 6483 15423 6541 15457
rect 6575 15423 6633 15457
rect 6667 15423 6725 15457
rect 6759 15423 6817 15457
rect 6851 15423 6909 15457
rect 6943 15423 7001 15457
rect 7035 15423 7093 15457
rect 7127 15423 7185 15457
rect 7219 15423 7277 15457
rect 7311 15423 7369 15457
rect 7403 15423 7461 15457
rect 7495 15423 7553 15457
rect 7587 15423 7645 15457
rect 7679 15423 7737 15457
rect 7771 15423 7829 15457
rect 7863 15423 7921 15457
rect 7955 15423 8013 15457
rect 8047 15423 8105 15457
rect 8139 15423 8197 15457
rect 8231 15423 8289 15457
rect 8323 15423 8381 15457
rect 8415 15423 8473 15457
rect 8507 15423 8565 15457
rect 8599 15423 8657 15457
rect 8691 15423 8749 15457
rect 8783 15423 8841 15457
rect 8875 15423 8933 15457
rect 8967 15423 9025 15457
rect 9059 15423 9117 15457
rect 9151 15423 9209 15457
rect 9243 15423 9301 15457
rect 9335 15423 9393 15457
rect 9427 15423 9485 15457
rect 9519 15423 9577 15457
rect 9611 15423 9669 15457
rect 9703 15423 9761 15457
rect 9795 15423 9853 15457
rect 6351 15414 9861 15423
rect 9913 15414 9925 15466
rect 9977 15457 9989 15466
rect 10041 15457 10053 15466
rect 9979 15423 9989 15457
rect 9977 15414 9989 15423
rect 10041 15414 10053 15423
rect 10105 15414 10117 15466
rect 10169 15457 13679 15466
rect 13731 15457 13743 15466
rect 10169 15423 10221 15457
rect 10255 15423 10313 15457
rect 10347 15423 10405 15457
rect 10439 15423 10497 15457
rect 10531 15423 10589 15457
rect 10623 15423 10681 15457
rect 10715 15423 10773 15457
rect 10807 15423 10865 15457
rect 10899 15423 10957 15457
rect 10991 15423 11049 15457
rect 11083 15423 11141 15457
rect 11175 15423 11233 15457
rect 11267 15423 11325 15457
rect 11359 15423 11417 15457
rect 11451 15423 11509 15457
rect 11543 15423 11601 15457
rect 11635 15423 11693 15457
rect 11727 15423 11785 15457
rect 11819 15423 11877 15457
rect 11911 15423 11969 15457
rect 12003 15423 12061 15457
rect 12095 15423 12153 15457
rect 12187 15423 12245 15457
rect 12279 15423 12337 15457
rect 12371 15423 12429 15457
rect 12463 15423 12521 15457
rect 12555 15423 12613 15457
rect 12647 15423 12705 15457
rect 12739 15423 12797 15457
rect 12831 15423 12889 15457
rect 12923 15423 12981 15457
rect 13015 15423 13073 15457
rect 13107 15423 13165 15457
rect 13199 15423 13257 15457
rect 13291 15423 13349 15457
rect 13383 15423 13441 15457
rect 13475 15423 13533 15457
rect 13567 15423 13625 15457
rect 13659 15423 13679 15457
rect 10169 15414 13679 15423
rect 13731 15414 13743 15423
rect 13795 15414 13807 15466
rect 13859 15414 13871 15466
rect 13923 15457 13935 15466
rect 13923 15414 13935 15423
rect 13987 15457 17497 15466
rect 13987 15423 13993 15457
rect 14027 15423 14085 15457
rect 14119 15423 14177 15457
rect 14211 15423 14269 15457
rect 14303 15423 14361 15457
rect 14395 15423 14453 15457
rect 14487 15423 14545 15457
rect 14579 15423 14637 15457
rect 14671 15423 14729 15457
rect 14763 15423 14821 15457
rect 14855 15423 14913 15457
rect 14947 15423 15005 15457
rect 15039 15423 15097 15457
rect 15131 15423 15189 15457
rect 15223 15423 15281 15457
rect 15315 15423 15373 15457
rect 15407 15423 15465 15457
rect 15499 15423 15557 15457
rect 15591 15423 15649 15457
rect 15683 15423 15741 15457
rect 15775 15423 15833 15457
rect 15867 15423 15925 15457
rect 15959 15423 16017 15457
rect 16051 15423 16109 15457
rect 16143 15423 16201 15457
rect 16235 15423 16293 15457
rect 16327 15423 16385 15457
rect 16419 15423 16477 15457
rect 16511 15423 16569 15457
rect 16603 15423 16661 15457
rect 16695 15423 16753 15457
rect 16787 15423 16845 15457
rect 16879 15423 16937 15457
rect 16971 15423 17029 15457
rect 17063 15423 17121 15457
rect 17155 15423 17213 15457
rect 17247 15423 17305 15457
rect 17339 15423 17397 15457
rect 17431 15423 17489 15457
rect 13987 15414 17497 15423
rect 17549 15414 17561 15466
rect 17613 15457 17625 15466
rect 17677 15457 17689 15466
rect 17615 15423 17625 15457
rect 17613 15414 17625 15423
rect 17677 15414 17689 15423
rect 17741 15414 17753 15466
rect 17805 15457 20220 15466
rect 17805 15423 17857 15457
rect 17891 15423 17949 15457
rect 17983 15423 18041 15457
rect 18075 15423 18133 15457
rect 18167 15423 18225 15457
rect 18259 15423 18317 15457
rect 18351 15423 18409 15457
rect 18443 15423 18501 15457
rect 18535 15423 18593 15457
rect 18627 15423 18685 15457
rect 18719 15423 18777 15457
rect 18811 15423 18869 15457
rect 18903 15423 18961 15457
rect 18995 15423 19053 15457
rect 19087 15423 19145 15457
rect 19179 15423 19237 15457
rect 19271 15423 19329 15457
rect 19363 15423 19421 15457
rect 19455 15423 19513 15457
rect 19547 15423 19605 15457
rect 19639 15423 19697 15457
rect 19731 15423 19789 15457
rect 19823 15423 19881 15457
rect 19915 15423 19973 15457
rect 20007 15423 20065 15457
rect 20099 15423 20157 15457
rect 20191 15423 20220 15457
rect 17805 15414 20220 15423
rect 4948 15392 20220 15414
rect 12874 15108 12880 15160
rect 12932 15108 12938 15160
rect 15358 15108 15364 15160
rect 15416 15108 15422 15160
rect 13426 14972 13432 15024
rect 13484 14972 13490 15024
rect 16005 15015 16063 15021
rect 16005 14981 16017 15015
rect 16051 15012 16063 15015
rect 16094 15012 16100 15024
rect 16051 14984 16100 15012
rect 16051 14981 16063 14984
rect 16005 14975 16063 14981
rect 16094 14972 16100 14984
rect 16152 14972 16158 15024
rect 4948 14922 20220 14944
rect 4948 14913 6703 14922
rect 6755 14913 6767 14922
rect 6819 14913 6831 14922
rect 4948 14879 4977 14913
rect 5011 14879 5069 14913
rect 5103 14879 5161 14913
rect 5195 14879 5253 14913
rect 5287 14879 5345 14913
rect 5379 14879 5437 14913
rect 5471 14879 5529 14913
rect 5563 14879 5621 14913
rect 5655 14879 5713 14913
rect 5747 14879 5805 14913
rect 5839 14879 5897 14913
rect 5931 14879 5989 14913
rect 6023 14879 6081 14913
rect 6115 14879 6173 14913
rect 6207 14879 6265 14913
rect 6299 14879 6357 14913
rect 6391 14879 6449 14913
rect 6483 14879 6541 14913
rect 6575 14879 6633 14913
rect 6667 14879 6703 14913
rect 6759 14879 6767 14913
rect 4948 14870 6703 14879
rect 6755 14870 6767 14879
rect 6819 14870 6831 14879
rect 6883 14870 6895 14922
rect 6947 14870 6959 14922
rect 7011 14913 10521 14922
rect 7035 14879 7093 14913
rect 7127 14879 7185 14913
rect 7219 14879 7277 14913
rect 7311 14879 7369 14913
rect 7403 14879 7461 14913
rect 7495 14879 7553 14913
rect 7587 14879 7645 14913
rect 7679 14879 7737 14913
rect 7771 14879 7829 14913
rect 7863 14879 7921 14913
rect 7955 14879 8013 14913
rect 8047 14879 8105 14913
rect 8139 14879 8197 14913
rect 8231 14879 8289 14913
rect 8323 14879 8381 14913
rect 8415 14879 8473 14913
rect 8507 14879 8565 14913
rect 8599 14879 8657 14913
rect 8691 14879 8749 14913
rect 8783 14879 8841 14913
rect 8875 14879 8933 14913
rect 8967 14879 9025 14913
rect 9059 14879 9117 14913
rect 9151 14879 9209 14913
rect 9243 14879 9301 14913
rect 9335 14879 9393 14913
rect 9427 14879 9485 14913
rect 9519 14879 9577 14913
rect 9611 14879 9669 14913
rect 9703 14879 9761 14913
rect 9795 14879 9853 14913
rect 9887 14879 9945 14913
rect 9979 14879 10037 14913
rect 10071 14879 10129 14913
rect 10163 14879 10221 14913
rect 10255 14879 10313 14913
rect 10347 14879 10405 14913
rect 10439 14879 10497 14913
rect 7011 14870 10521 14879
rect 10573 14870 10585 14922
rect 10637 14870 10649 14922
rect 10701 14913 10713 14922
rect 10765 14913 10777 14922
rect 10829 14913 14339 14922
rect 14391 14913 14403 14922
rect 14455 14913 14467 14922
rect 10765 14879 10773 14913
rect 10829 14879 10865 14913
rect 10899 14879 10957 14913
rect 10991 14879 11049 14913
rect 11083 14879 11141 14913
rect 11175 14879 11233 14913
rect 11267 14879 11325 14913
rect 11359 14879 11417 14913
rect 11451 14879 11509 14913
rect 11543 14879 11601 14913
rect 11635 14879 11693 14913
rect 11727 14879 11785 14913
rect 11819 14879 11877 14913
rect 11911 14879 11969 14913
rect 12003 14879 12061 14913
rect 12095 14879 12153 14913
rect 12187 14879 12245 14913
rect 12279 14879 12337 14913
rect 12371 14879 12429 14913
rect 12463 14879 12521 14913
rect 12555 14879 12613 14913
rect 12647 14879 12705 14913
rect 12739 14879 12797 14913
rect 12831 14879 12889 14913
rect 12923 14879 12981 14913
rect 13015 14879 13073 14913
rect 13107 14879 13165 14913
rect 13199 14879 13257 14913
rect 13291 14879 13349 14913
rect 13383 14879 13441 14913
rect 13475 14879 13533 14913
rect 13567 14879 13625 14913
rect 13659 14879 13717 14913
rect 13751 14879 13809 14913
rect 13843 14879 13901 14913
rect 13935 14879 13993 14913
rect 14027 14879 14085 14913
rect 14119 14879 14177 14913
rect 14211 14879 14269 14913
rect 14303 14879 14339 14913
rect 14395 14879 14403 14913
rect 10701 14870 10713 14879
rect 10765 14870 10777 14879
rect 10829 14870 14339 14879
rect 14391 14870 14403 14879
rect 14455 14870 14467 14879
rect 14519 14870 14531 14922
rect 14583 14870 14595 14922
rect 14647 14913 18157 14922
rect 14671 14879 14729 14913
rect 14763 14879 14821 14913
rect 14855 14879 14913 14913
rect 14947 14879 15005 14913
rect 15039 14879 15097 14913
rect 15131 14879 15189 14913
rect 15223 14879 15281 14913
rect 15315 14879 15373 14913
rect 15407 14879 15465 14913
rect 15499 14879 15557 14913
rect 15591 14879 15649 14913
rect 15683 14879 15741 14913
rect 15775 14879 15833 14913
rect 15867 14879 15925 14913
rect 15959 14879 16017 14913
rect 16051 14879 16109 14913
rect 16143 14879 16201 14913
rect 16235 14879 16293 14913
rect 16327 14879 16385 14913
rect 16419 14879 16477 14913
rect 16511 14879 16569 14913
rect 16603 14879 16661 14913
rect 16695 14879 16753 14913
rect 16787 14879 16845 14913
rect 16879 14879 16937 14913
rect 16971 14879 17029 14913
rect 17063 14879 17121 14913
rect 17155 14879 17213 14913
rect 17247 14879 17305 14913
rect 17339 14879 17397 14913
rect 17431 14879 17489 14913
rect 17523 14879 17581 14913
rect 17615 14879 17673 14913
rect 17707 14879 17765 14913
rect 17799 14879 17857 14913
rect 17891 14879 17949 14913
rect 17983 14879 18041 14913
rect 18075 14879 18133 14913
rect 14647 14870 18157 14879
rect 18209 14870 18221 14922
rect 18273 14870 18285 14922
rect 18337 14913 18349 14922
rect 18401 14913 18413 14922
rect 18465 14913 20220 14922
rect 18401 14879 18409 14913
rect 18465 14879 18501 14913
rect 18535 14879 18593 14913
rect 18627 14879 18685 14913
rect 18719 14879 18777 14913
rect 18811 14879 18869 14913
rect 18903 14879 18961 14913
rect 18995 14879 19053 14913
rect 19087 14879 19145 14913
rect 19179 14879 19237 14913
rect 19271 14879 19329 14913
rect 19363 14879 19421 14913
rect 19455 14879 19513 14913
rect 19547 14879 19605 14913
rect 19639 14879 19697 14913
rect 19731 14879 19789 14913
rect 19823 14879 19881 14913
rect 19915 14879 19973 14913
rect 20007 14879 20065 14913
rect 20099 14879 20157 14913
rect 20191 14879 20220 14913
rect 18337 14870 18349 14879
rect 18401 14870 18413 14879
rect 18465 14870 20220 14879
rect 4948 14848 20220 14870
rect 13426 14808 13432 14820
rect 13076 14780 13432 14808
rect 10853 14675 10911 14681
rect 10853 14641 10865 14675
rect 10899 14672 10911 14675
rect 11678 14672 11684 14684
rect 10899 14644 11684 14672
rect 10899 14641 10911 14644
rect 10853 14635 10911 14641
rect 11678 14632 11684 14644
rect 11736 14672 11742 14684
rect 12877 14675 12935 14681
rect 12877 14672 12889 14675
rect 11736 14644 12889 14672
rect 11736 14632 11742 14644
rect 12877 14641 12889 14644
rect 12923 14641 12935 14675
rect 12877 14635 12935 14641
rect 11034 14564 11040 14616
rect 11092 14564 11098 14616
rect 12892 14536 12920 14635
rect 13076 14613 13104 14780
rect 13426 14768 13432 14780
rect 13484 14768 13490 14820
rect 14441 14743 14499 14749
rect 14441 14709 14453 14743
rect 14487 14740 14499 14743
rect 14990 14740 14996 14752
rect 14487 14712 14996 14740
rect 14487 14709 14499 14712
rect 14441 14703 14499 14709
rect 14990 14700 14996 14712
rect 15048 14700 15054 14752
rect 15105 14743 15163 14749
rect 15105 14709 15117 14743
rect 15151 14740 15163 14743
rect 15729 14743 15787 14749
rect 15729 14740 15741 14743
rect 15151 14712 15741 14740
rect 15151 14709 15163 14712
rect 15105 14703 15163 14709
rect 15729 14709 15741 14712
rect 15775 14740 15787 14743
rect 16107 14743 16165 14749
rect 16107 14740 16119 14743
rect 15775 14712 16119 14740
rect 15775 14709 15787 14712
rect 15729 14703 15787 14709
rect 16107 14709 16119 14712
rect 16153 14709 16165 14743
rect 16107 14703 16165 14709
rect 13061 14607 13119 14613
rect 13061 14573 13073 14607
rect 13107 14573 13119 14607
rect 13061 14567 13119 14573
rect 14254 14564 14260 14616
rect 14312 14564 14318 14616
rect 14889 14602 14947 14608
rect 14889 14568 14901 14602
rect 14935 14568 14947 14602
rect 14889 14545 14947 14568
rect 15105 14607 15163 14613
rect 15105 14573 15117 14607
rect 15151 14604 15163 14607
rect 15821 14607 15879 14613
rect 15821 14604 15833 14607
rect 15151 14576 15833 14604
rect 15151 14573 15163 14576
rect 15105 14567 15163 14573
rect 15821 14573 15833 14576
rect 15867 14604 15879 14607
rect 16188 14607 16246 14613
rect 16188 14604 16200 14607
rect 15867 14576 16200 14604
rect 15867 14573 15879 14576
rect 15821 14567 15879 14573
rect 16188 14573 16200 14576
rect 16234 14573 16246 14607
rect 16188 14567 16246 14573
rect 16278 14564 16284 14616
rect 16336 14564 16342 14616
rect 15542 14545 15548 14548
rect 14829 14539 14947 14545
rect 12892 14508 14392 14536
rect 14364 14480 14392 14508
rect 14829 14505 14841 14539
rect 14875 14536 14947 14539
rect 15477 14539 15548 14545
rect 15600 14545 15606 14548
rect 15477 14536 15489 14539
rect 14875 14508 15489 14536
rect 14875 14505 14887 14508
rect 14829 14499 14887 14505
rect 15477 14505 15489 14508
rect 15523 14505 15548 14539
rect 15477 14499 15548 14505
rect 15542 14496 15548 14499
rect 15600 14499 15607 14545
rect 15600 14496 15606 14499
rect 16002 14496 16008 14548
rect 16060 14496 16066 14548
rect 10206 14428 10212 14480
rect 10264 14468 10270 14480
rect 10945 14471 11003 14477
rect 10945 14468 10957 14471
rect 10264 14440 10957 14468
rect 10264 14428 10270 14440
rect 10945 14437 10957 14440
rect 10991 14437 11003 14471
rect 10945 14431 11003 14437
rect 11402 14428 11408 14480
rect 11460 14428 11466 14480
rect 12969 14471 13027 14477
rect 12969 14437 12981 14471
rect 13015 14468 13027 14471
rect 13058 14468 13064 14480
rect 13015 14440 13064 14468
rect 13015 14437 13027 14440
rect 12969 14431 13027 14437
rect 13058 14428 13064 14440
rect 13116 14428 13122 14480
rect 13426 14428 13432 14480
rect 13484 14428 13490 14480
rect 14346 14428 14352 14480
rect 14404 14428 14410 14480
rect 14533 14471 14591 14477
rect 14533 14437 14545 14471
rect 14579 14468 14591 14471
rect 15634 14468 15640 14480
rect 14579 14440 15640 14468
rect 14579 14437 14591 14440
rect 14533 14431 14591 14437
rect 15634 14428 15640 14440
rect 15692 14428 15698 14480
rect 4948 14378 20220 14400
rect 4948 14369 6043 14378
rect 6095 14369 6107 14378
rect 4948 14335 4977 14369
rect 5011 14335 5069 14369
rect 5103 14335 5161 14369
rect 5195 14335 5253 14369
rect 5287 14335 5345 14369
rect 5379 14335 5437 14369
rect 5471 14335 5529 14369
rect 5563 14335 5621 14369
rect 5655 14335 5713 14369
rect 5747 14335 5805 14369
rect 5839 14335 5897 14369
rect 5931 14335 5989 14369
rect 6023 14335 6043 14369
rect 4948 14326 6043 14335
rect 6095 14326 6107 14335
rect 6159 14326 6171 14378
rect 6223 14326 6235 14378
rect 6287 14369 6299 14378
rect 6287 14326 6299 14335
rect 6351 14369 9861 14378
rect 6351 14335 6357 14369
rect 6391 14335 6449 14369
rect 6483 14335 6541 14369
rect 6575 14335 6633 14369
rect 6667 14335 6725 14369
rect 6759 14335 6817 14369
rect 6851 14335 6909 14369
rect 6943 14335 7001 14369
rect 7035 14335 7093 14369
rect 7127 14335 7185 14369
rect 7219 14335 7277 14369
rect 7311 14335 7369 14369
rect 7403 14335 7461 14369
rect 7495 14335 7553 14369
rect 7587 14335 7645 14369
rect 7679 14335 7737 14369
rect 7771 14335 7829 14369
rect 7863 14335 7921 14369
rect 7955 14335 8013 14369
rect 8047 14335 8105 14369
rect 8139 14335 8197 14369
rect 8231 14335 8289 14369
rect 8323 14335 8381 14369
rect 8415 14335 8473 14369
rect 8507 14335 8565 14369
rect 8599 14335 8657 14369
rect 8691 14335 8749 14369
rect 8783 14335 8841 14369
rect 8875 14335 8933 14369
rect 8967 14335 9025 14369
rect 9059 14335 9117 14369
rect 9151 14335 9209 14369
rect 9243 14335 9301 14369
rect 9335 14335 9393 14369
rect 9427 14335 9485 14369
rect 9519 14335 9577 14369
rect 9611 14335 9669 14369
rect 9703 14335 9761 14369
rect 9795 14335 9853 14369
rect 6351 14326 9861 14335
rect 9913 14326 9925 14378
rect 9977 14369 9989 14378
rect 10041 14369 10053 14378
rect 9979 14335 9989 14369
rect 9977 14326 9989 14335
rect 10041 14326 10053 14335
rect 10105 14326 10117 14378
rect 10169 14369 13679 14378
rect 13731 14369 13743 14378
rect 10169 14335 10221 14369
rect 10255 14335 10313 14369
rect 10347 14335 10405 14369
rect 10439 14335 10497 14369
rect 10531 14335 10589 14369
rect 10623 14335 10681 14369
rect 10715 14335 10773 14369
rect 10807 14335 10865 14369
rect 10899 14335 10957 14369
rect 10991 14335 11049 14369
rect 11083 14335 11141 14369
rect 11175 14335 11233 14369
rect 11267 14335 11325 14369
rect 11359 14335 11417 14369
rect 11451 14335 11509 14369
rect 11543 14335 11601 14369
rect 11635 14335 11693 14369
rect 11727 14335 11785 14369
rect 11819 14335 11877 14369
rect 11911 14335 11969 14369
rect 12003 14335 12061 14369
rect 12095 14335 12153 14369
rect 12187 14335 12245 14369
rect 12279 14335 12337 14369
rect 12371 14335 12429 14369
rect 12463 14335 12521 14369
rect 12555 14335 12613 14369
rect 12647 14335 12705 14369
rect 12739 14335 12797 14369
rect 12831 14335 12889 14369
rect 12923 14335 12981 14369
rect 13015 14335 13073 14369
rect 13107 14335 13165 14369
rect 13199 14335 13257 14369
rect 13291 14335 13349 14369
rect 13383 14335 13441 14369
rect 13475 14335 13533 14369
rect 13567 14335 13625 14369
rect 13659 14335 13679 14369
rect 10169 14326 13679 14335
rect 13731 14326 13743 14335
rect 13795 14326 13807 14378
rect 13859 14326 13871 14378
rect 13923 14369 13935 14378
rect 13923 14326 13935 14335
rect 13987 14369 17497 14378
rect 13987 14335 13993 14369
rect 14027 14335 14085 14369
rect 14119 14335 14177 14369
rect 14211 14335 14269 14369
rect 14303 14335 14361 14369
rect 14395 14335 14453 14369
rect 14487 14335 14545 14369
rect 14579 14335 14637 14369
rect 14671 14335 14729 14369
rect 14763 14335 14821 14369
rect 14855 14335 14913 14369
rect 14947 14335 15005 14369
rect 15039 14335 15097 14369
rect 15131 14335 15189 14369
rect 15223 14335 15281 14369
rect 15315 14335 15373 14369
rect 15407 14335 15465 14369
rect 15499 14335 15557 14369
rect 15591 14335 15649 14369
rect 15683 14335 15741 14369
rect 15775 14335 15833 14369
rect 15867 14335 15925 14369
rect 15959 14335 16017 14369
rect 16051 14335 16109 14369
rect 16143 14335 16201 14369
rect 16235 14335 16293 14369
rect 16327 14335 16385 14369
rect 16419 14335 16477 14369
rect 16511 14335 16569 14369
rect 16603 14335 16661 14369
rect 16695 14335 16753 14369
rect 16787 14335 16845 14369
rect 16879 14335 16937 14369
rect 16971 14335 17029 14369
rect 17063 14335 17121 14369
rect 17155 14335 17213 14369
rect 17247 14335 17305 14369
rect 17339 14335 17397 14369
rect 17431 14335 17489 14369
rect 13987 14326 17497 14335
rect 17549 14326 17561 14378
rect 17613 14369 17625 14378
rect 17677 14369 17689 14378
rect 17615 14335 17625 14369
rect 17613 14326 17625 14335
rect 17677 14326 17689 14335
rect 17741 14326 17753 14378
rect 17805 14369 20220 14378
rect 17805 14335 17857 14369
rect 17891 14335 17949 14369
rect 17983 14335 18041 14369
rect 18075 14335 18133 14369
rect 18167 14335 18225 14369
rect 18259 14335 18317 14369
rect 18351 14335 18409 14369
rect 18443 14335 18501 14369
rect 18535 14335 18593 14369
rect 18627 14335 18685 14369
rect 18719 14335 18777 14369
rect 18811 14335 18869 14369
rect 18903 14335 18961 14369
rect 18995 14335 19053 14369
rect 19087 14335 19145 14369
rect 19179 14335 19237 14369
rect 19271 14335 19329 14369
rect 19363 14335 19421 14369
rect 19455 14335 19513 14369
rect 19547 14335 19605 14369
rect 19639 14335 19697 14369
rect 19731 14335 19789 14369
rect 19823 14335 19881 14369
rect 19915 14335 19973 14369
rect 20007 14335 20065 14369
rect 20099 14335 20157 14369
rect 20191 14335 20220 14369
rect 17805 14326 20220 14335
rect 4948 14304 20220 14326
rect 11402 14224 11408 14276
rect 11460 14224 11466 14276
rect 15177 14267 15235 14273
rect 15177 14233 15189 14267
rect 15223 14264 15235 14267
rect 15358 14264 15364 14276
rect 15223 14236 15364 14264
rect 15223 14233 15235 14236
rect 15177 14227 15235 14233
rect 15358 14224 15364 14236
rect 15416 14224 15422 14276
rect 15634 14224 15640 14276
rect 15692 14224 15698 14276
rect 16002 14224 16008 14276
rect 16060 14224 16066 14276
rect 16094 14224 16100 14276
rect 16152 14224 16158 14276
rect 5790 14156 5796 14208
rect 5848 14196 5854 14208
rect 10413 14199 10471 14205
rect 10413 14196 10425 14199
rect 5848 14168 10425 14196
rect 5848 14156 5854 14168
rect 10408 14165 10425 14168
rect 10459 14196 10471 14199
rect 11061 14199 11191 14205
rect 11061 14196 11073 14199
rect 10459 14168 11073 14196
rect 10459 14165 10531 14168
rect 10408 14159 10531 14165
rect 11061 14165 11073 14168
rect 11107 14165 11145 14199
rect 11179 14165 11191 14199
rect 11420 14196 11448 14224
rect 11420 14168 11908 14196
rect 11061 14159 11191 14165
rect 10408 14060 10436 14159
rect 10473 14136 10531 14159
rect 10473 14102 10485 14136
rect 10519 14102 10531 14136
rect 10473 14096 10531 14102
rect 10689 14131 10747 14137
rect 10689 14097 10701 14131
rect 10735 14128 10747 14131
rect 11405 14131 11463 14137
rect 11405 14128 11417 14131
rect 10735 14100 11417 14128
rect 10735 14097 10747 14100
rect 10689 14091 10747 14097
rect 11405 14097 11417 14100
rect 11451 14128 11463 14131
rect 11772 14131 11830 14137
rect 11772 14128 11784 14131
rect 11451 14100 11784 14128
rect 11451 14097 11463 14100
rect 11405 14091 11463 14097
rect 11772 14097 11784 14100
rect 11818 14097 11830 14131
rect 11880 14128 11908 14168
rect 13978 14156 13984 14208
rect 14036 14156 14042 14208
rect 12141 14131 12199 14137
rect 12141 14128 12153 14131
rect 11880 14100 12153 14128
rect 11772 14091 11830 14097
rect 12141 14097 12153 14100
rect 12187 14097 12199 14131
rect 12141 14091 12199 14097
rect 14901 14131 14959 14137
rect 14901 14097 14913 14131
rect 14947 14128 14959 14131
rect 15545 14131 15603 14137
rect 15545 14128 15557 14131
rect 14947 14100 15557 14128
rect 14947 14097 14959 14100
rect 14901 14091 14959 14097
rect 15545 14097 15557 14100
rect 15591 14097 15603 14131
rect 16112 14128 16140 14224
rect 16189 14131 16247 14137
rect 16189 14128 16201 14131
rect 16112 14100 16201 14128
rect 15545 14091 15603 14097
rect 16189 14097 16201 14100
rect 16235 14097 16247 14131
rect 16189 14091 16247 14097
rect 16462 14088 16468 14140
rect 16520 14088 16526 14140
rect 10850 14060 10856 14072
rect 10408 14032 10856 14060
rect 10850 14020 10856 14032
rect 10908 14020 10914 14072
rect 11589 14063 11647 14069
rect 11589 14029 11601 14063
rect 11635 14060 11647 14063
rect 11635 14032 11816 14060
rect 11635 14029 11647 14032
rect 11589 14023 11647 14029
rect 10689 13995 10747 14001
rect 10689 13961 10701 13995
rect 10735 13992 10747 13995
rect 11313 13995 11371 14001
rect 11313 13992 11325 13995
rect 10735 13964 11325 13992
rect 10735 13961 10747 13964
rect 10689 13955 10747 13961
rect 11313 13961 11325 13964
rect 11359 13992 11371 13995
rect 11691 13995 11749 14001
rect 11691 13992 11703 13995
rect 11359 13964 11703 13992
rect 11359 13961 11371 13964
rect 11313 13955 11371 13961
rect 11691 13961 11703 13964
rect 11737 13961 11749 13995
rect 11691 13955 11749 13961
rect 10117 13927 10175 13933
rect 10117 13893 10129 13927
rect 10163 13924 10175 13927
rect 10206 13924 10212 13936
rect 10163 13896 10212 13924
rect 10163 13893 10175 13896
rect 10117 13887 10175 13893
rect 10206 13884 10212 13896
rect 10264 13884 10270 13936
rect 11788 13924 11816 14032
rect 11862 14020 11868 14072
rect 11920 14020 11926 14072
rect 14162 14020 14168 14072
rect 14220 14060 14226 14072
rect 14257 14063 14315 14069
rect 14257 14060 14269 14063
rect 14220 14032 14269 14060
rect 14220 14020 14226 14032
rect 14257 14029 14269 14032
rect 14303 14029 14315 14063
rect 14257 14023 14315 14029
rect 14346 14020 14352 14072
rect 14404 14060 14410 14072
rect 14806 14060 14812 14072
rect 14404 14032 14812 14060
rect 14404 14020 14410 14032
rect 14806 14020 14812 14032
rect 14864 14060 14870 14072
rect 15821 14063 15879 14069
rect 15821 14060 15833 14063
rect 14864 14032 15833 14060
rect 14864 14020 14870 14032
rect 15821 14029 15833 14032
rect 15867 14060 15879 14063
rect 15867 14032 17152 14060
rect 15867 14029 15879 14032
rect 15821 14023 15879 14029
rect 11957 13995 12015 14001
rect 11957 13961 11969 13995
rect 12003 13961 12015 13995
rect 11957 13955 12015 13961
rect 11972 13924 12000 13955
rect 17124 13936 17152 14032
rect 11788 13896 12000 13924
rect 12690 13884 12696 13936
rect 12748 13924 12754 13936
rect 14714 13924 14720 13936
rect 12748 13896 14720 13924
rect 12748 13884 12754 13896
rect 14714 13884 14720 13896
rect 14772 13884 14778 13936
rect 15726 13884 15732 13936
rect 15784 13924 15790 13936
rect 16281 13927 16339 13933
rect 16281 13924 16293 13927
rect 15784 13896 16293 13924
rect 15784 13884 15790 13896
rect 16281 13893 16293 13896
rect 16327 13893 16339 13927
rect 16281 13887 16339 13893
rect 17106 13884 17112 13936
rect 17164 13884 17170 13936
rect 4948 13834 20220 13856
rect 4948 13825 6703 13834
rect 6755 13825 6767 13834
rect 6819 13825 6831 13834
rect 4948 13791 4977 13825
rect 5011 13791 5069 13825
rect 5103 13791 5161 13825
rect 5195 13791 5253 13825
rect 5287 13791 5345 13825
rect 5379 13791 5437 13825
rect 5471 13791 5529 13825
rect 5563 13791 5621 13825
rect 5655 13791 5713 13825
rect 5747 13791 5805 13825
rect 5839 13791 5897 13825
rect 5931 13791 5989 13825
rect 6023 13791 6081 13825
rect 6115 13791 6173 13825
rect 6207 13791 6265 13825
rect 6299 13791 6357 13825
rect 6391 13791 6449 13825
rect 6483 13791 6541 13825
rect 6575 13791 6633 13825
rect 6667 13791 6703 13825
rect 6759 13791 6767 13825
rect 4948 13782 6703 13791
rect 6755 13782 6767 13791
rect 6819 13782 6831 13791
rect 6883 13782 6895 13834
rect 6947 13782 6959 13834
rect 7011 13825 10521 13834
rect 7035 13791 7093 13825
rect 7127 13791 7185 13825
rect 7219 13791 7277 13825
rect 7311 13791 7369 13825
rect 7403 13791 7461 13825
rect 7495 13791 7553 13825
rect 7587 13791 7645 13825
rect 7679 13791 7737 13825
rect 7771 13791 7829 13825
rect 7863 13791 7921 13825
rect 7955 13791 8013 13825
rect 8047 13791 8105 13825
rect 8139 13791 8197 13825
rect 8231 13791 8289 13825
rect 8323 13791 8381 13825
rect 8415 13791 8473 13825
rect 8507 13791 8565 13825
rect 8599 13791 8657 13825
rect 8691 13791 8749 13825
rect 8783 13791 8841 13825
rect 8875 13791 8933 13825
rect 8967 13791 9025 13825
rect 9059 13791 9117 13825
rect 9151 13791 9209 13825
rect 9243 13791 9301 13825
rect 9335 13791 9393 13825
rect 9427 13791 9485 13825
rect 9519 13791 9577 13825
rect 9611 13791 9669 13825
rect 9703 13791 9761 13825
rect 9795 13791 9853 13825
rect 9887 13791 9945 13825
rect 9979 13791 10037 13825
rect 10071 13791 10129 13825
rect 10163 13791 10221 13825
rect 10255 13791 10313 13825
rect 10347 13791 10405 13825
rect 10439 13791 10497 13825
rect 7011 13782 10521 13791
rect 10573 13782 10585 13834
rect 10637 13782 10649 13834
rect 10701 13825 10713 13834
rect 10765 13825 10777 13834
rect 10829 13825 14339 13834
rect 14391 13825 14403 13834
rect 14455 13825 14467 13834
rect 10765 13791 10773 13825
rect 10829 13791 10865 13825
rect 10899 13791 10957 13825
rect 10991 13791 11049 13825
rect 11083 13791 11141 13825
rect 11175 13791 11233 13825
rect 11267 13791 11325 13825
rect 11359 13791 11417 13825
rect 11451 13791 11509 13825
rect 11543 13791 11601 13825
rect 11635 13791 11693 13825
rect 11727 13791 11785 13825
rect 11819 13791 11877 13825
rect 11911 13791 11969 13825
rect 12003 13791 12061 13825
rect 12095 13791 12153 13825
rect 12187 13791 12245 13825
rect 12279 13791 12337 13825
rect 12371 13791 12429 13825
rect 12463 13791 12521 13825
rect 12555 13791 12613 13825
rect 12647 13791 12705 13825
rect 12739 13791 12797 13825
rect 12831 13791 12889 13825
rect 12923 13791 12981 13825
rect 13015 13791 13073 13825
rect 13107 13791 13165 13825
rect 13199 13791 13257 13825
rect 13291 13791 13349 13825
rect 13383 13791 13441 13825
rect 13475 13791 13533 13825
rect 13567 13791 13625 13825
rect 13659 13791 13717 13825
rect 13751 13791 13809 13825
rect 13843 13791 13901 13825
rect 13935 13791 13993 13825
rect 14027 13791 14085 13825
rect 14119 13791 14177 13825
rect 14211 13791 14269 13825
rect 14303 13791 14339 13825
rect 14395 13791 14403 13825
rect 10701 13782 10713 13791
rect 10765 13782 10777 13791
rect 10829 13782 14339 13791
rect 14391 13782 14403 13791
rect 14455 13782 14467 13791
rect 14519 13782 14531 13834
rect 14583 13782 14595 13834
rect 14647 13825 18157 13834
rect 14671 13791 14729 13825
rect 14763 13791 14821 13825
rect 14855 13791 14913 13825
rect 14947 13791 15005 13825
rect 15039 13791 15097 13825
rect 15131 13791 15189 13825
rect 15223 13791 15281 13825
rect 15315 13791 15373 13825
rect 15407 13791 15465 13825
rect 15499 13791 15557 13825
rect 15591 13791 15649 13825
rect 15683 13791 15741 13825
rect 15775 13791 15833 13825
rect 15867 13791 15925 13825
rect 15959 13791 16017 13825
rect 16051 13791 16109 13825
rect 16143 13791 16201 13825
rect 16235 13791 16293 13825
rect 16327 13791 16385 13825
rect 16419 13791 16477 13825
rect 16511 13791 16569 13825
rect 16603 13791 16661 13825
rect 16695 13791 16753 13825
rect 16787 13791 16845 13825
rect 16879 13791 16937 13825
rect 16971 13791 17029 13825
rect 17063 13791 17121 13825
rect 17155 13791 17213 13825
rect 17247 13791 17305 13825
rect 17339 13791 17397 13825
rect 17431 13791 17489 13825
rect 17523 13791 17581 13825
rect 17615 13791 17673 13825
rect 17707 13791 17765 13825
rect 17799 13791 17857 13825
rect 17891 13791 17949 13825
rect 17983 13791 18041 13825
rect 18075 13791 18133 13825
rect 14647 13782 18157 13791
rect 18209 13782 18221 13834
rect 18273 13782 18285 13834
rect 18337 13825 18349 13834
rect 18401 13825 18413 13834
rect 18465 13825 20220 13834
rect 18401 13791 18409 13825
rect 18465 13791 18501 13825
rect 18535 13791 18593 13825
rect 18627 13791 18685 13825
rect 18719 13791 18777 13825
rect 18811 13791 18869 13825
rect 18903 13791 18961 13825
rect 18995 13791 19053 13825
rect 19087 13791 19145 13825
rect 19179 13791 19237 13825
rect 19271 13791 19329 13825
rect 19363 13791 19421 13825
rect 19455 13791 19513 13825
rect 19547 13791 19605 13825
rect 19639 13791 19697 13825
rect 19731 13791 19789 13825
rect 19823 13791 19881 13825
rect 19915 13791 19973 13825
rect 20007 13791 20065 13825
rect 20099 13791 20157 13825
rect 20191 13791 20220 13825
rect 18337 13782 18349 13791
rect 18401 13782 18413 13791
rect 18465 13782 20220 13791
rect 4948 13760 20220 13782
rect 10393 13723 10451 13729
rect 10393 13689 10405 13723
rect 10439 13720 10451 13723
rect 11862 13720 11868 13732
rect 10439 13692 11868 13720
rect 10439 13689 10451 13692
rect 10393 13683 10451 13689
rect 11862 13680 11868 13692
rect 11920 13680 11926 13732
rect 12690 13680 12696 13732
rect 12748 13680 12754 13732
rect 12877 13723 12935 13729
rect 12877 13689 12889 13723
rect 12923 13720 12935 13723
rect 13058 13720 13064 13732
rect 12923 13692 13064 13720
rect 12923 13689 12935 13692
rect 12877 13683 12935 13689
rect 13058 13680 13064 13692
rect 13116 13680 13122 13732
rect 16189 13723 16247 13729
rect 16189 13689 16201 13723
rect 16235 13720 16247 13723
rect 16278 13720 16284 13732
rect 16235 13692 16284 13720
rect 16235 13689 16247 13692
rect 16189 13683 16247 13689
rect 12708 13584 12736 13680
rect 13449 13655 13507 13661
rect 13449 13621 13461 13655
rect 13495 13652 13507 13655
rect 14073 13655 14131 13661
rect 14073 13652 14085 13655
rect 13495 13624 14085 13652
rect 13495 13621 13507 13624
rect 13449 13615 13507 13621
rect 14073 13621 14085 13624
rect 14119 13652 14131 13655
rect 14451 13655 14509 13661
rect 14451 13652 14463 13655
rect 14119 13624 14463 13652
rect 14119 13621 14131 13624
rect 14073 13615 14131 13621
rect 14451 13621 14463 13624
rect 14497 13621 14509 13655
rect 14451 13615 14509 13621
rect 11696 13556 12736 13584
rect 14625 13587 14683 13593
rect 9654 13476 9660 13528
rect 9712 13476 9718 13528
rect 10850 13476 10856 13528
rect 10908 13476 10914 13528
rect 11696 13525 11724 13556
rect 14625 13553 14637 13587
rect 14671 13584 14683 13587
rect 15082 13584 15088 13596
rect 14671 13556 15088 13584
rect 14671 13553 14683 13556
rect 14625 13547 14683 13553
rect 15082 13544 15088 13556
rect 15140 13584 15146 13596
rect 16204 13584 16232 13683
rect 16278 13680 16284 13692
rect 16336 13680 16342 13732
rect 16462 13680 16468 13732
rect 16520 13720 16526 13732
rect 16557 13723 16615 13729
rect 16557 13720 16569 13723
rect 16520 13692 16569 13720
rect 16520 13680 16526 13692
rect 16557 13689 16569 13692
rect 16603 13689 16615 13723
rect 16557 13683 16615 13689
rect 15140 13556 16232 13584
rect 15140 13544 15146 13556
rect 17106 13544 17112 13596
rect 17164 13584 17170 13596
rect 18762 13584 18768 13596
rect 17164 13556 18768 13584
rect 17164 13544 17170 13556
rect 18762 13544 18768 13556
rect 18820 13544 18826 13596
rect 11681 13519 11739 13525
rect 11681 13485 11693 13519
rect 11727 13485 11739 13519
rect 11681 13479 11739 13485
rect 12690 13476 12696 13528
rect 12748 13476 12754 13528
rect 13233 13514 13291 13520
rect 13233 13480 13245 13514
rect 13279 13480 13291 13514
rect 10868 13448 10896 13476
rect 13233 13457 13291 13480
rect 13449 13519 13507 13525
rect 13449 13485 13461 13519
rect 13495 13516 13507 13519
rect 14165 13519 14223 13525
rect 14165 13516 14177 13519
rect 13495 13488 14177 13516
rect 13495 13485 13507 13488
rect 13449 13479 13507 13485
rect 14165 13485 14177 13488
rect 14211 13516 14223 13519
rect 14532 13519 14590 13525
rect 14532 13516 14544 13519
rect 14211 13488 14544 13516
rect 14211 13485 14223 13488
rect 14165 13479 14223 13485
rect 14532 13485 14544 13488
rect 14578 13485 14590 13519
rect 14532 13479 14590 13485
rect 14714 13476 14720 13528
rect 14772 13476 14778 13528
rect 15634 13476 15640 13528
rect 15692 13516 15698 13528
rect 16922 13516 16928 13528
rect 15692 13488 16928 13516
rect 15692 13476 15698 13488
rect 16922 13476 16928 13488
rect 16980 13476 16986 13528
rect 13173 13451 13291 13457
rect 13173 13448 13185 13451
rect 10868 13420 13185 13448
rect 9841 13383 9899 13389
rect 9841 13349 9853 13383
rect 9887 13380 9899 13383
rect 10574 13380 10580 13392
rect 9887 13352 10580 13380
rect 9887 13349 9899 13352
rect 9841 13343 9899 13349
rect 10574 13340 10580 13352
rect 10632 13340 10638 13392
rect 12506 13340 12512 13392
rect 12564 13340 12570 13392
rect 13076 13380 13104 13420
rect 13173 13417 13185 13420
rect 13219 13448 13291 13451
rect 13821 13451 13951 13457
rect 13821 13448 13833 13451
rect 13219 13420 13833 13448
rect 13219 13417 13231 13420
rect 13173 13411 13231 13417
rect 13821 13417 13833 13420
rect 13867 13417 13905 13451
rect 13939 13417 13951 13451
rect 13821 13411 13951 13417
rect 14070 13408 14076 13460
rect 14128 13448 14134 13460
rect 14349 13451 14407 13457
rect 14349 13448 14361 13451
rect 14128 13420 14361 13448
rect 14128 13408 14134 13420
rect 14349 13417 14361 13420
rect 14395 13417 14407 13451
rect 14349 13411 14407 13417
rect 14438 13380 14444 13392
rect 13076 13352 14444 13380
rect 14438 13340 14444 13352
rect 14496 13340 14502 13392
rect 17014 13340 17020 13392
rect 17072 13340 17078 13392
rect 4948 13290 20220 13312
rect 4948 13281 6043 13290
rect 6095 13281 6107 13290
rect 4948 13247 4977 13281
rect 5011 13247 5069 13281
rect 5103 13247 5161 13281
rect 5195 13247 5253 13281
rect 5287 13247 5345 13281
rect 5379 13247 5437 13281
rect 5471 13247 5529 13281
rect 5563 13247 5621 13281
rect 5655 13247 5713 13281
rect 5747 13247 5805 13281
rect 5839 13247 5897 13281
rect 5931 13247 5989 13281
rect 6023 13247 6043 13281
rect 4948 13238 6043 13247
rect 6095 13238 6107 13247
rect 6159 13238 6171 13290
rect 6223 13238 6235 13290
rect 6287 13281 6299 13290
rect 6287 13238 6299 13247
rect 6351 13281 9861 13290
rect 6351 13247 6357 13281
rect 6391 13247 6449 13281
rect 6483 13247 6541 13281
rect 6575 13247 6633 13281
rect 6667 13247 6725 13281
rect 6759 13247 6817 13281
rect 6851 13247 6909 13281
rect 6943 13247 7001 13281
rect 7035 13247 7093 13281
rect 7127 13247 7185 13281
rect 7219 13247 7277 13281
rect 7311 13247 7369 13281
rect 7403 13247 7461 13281
rect 7495 13247 7553 13281
rect 7587 13247 7645 13281
rect 7679 13247 7737 13281
rect 7771 13247 7829 13281
rect 7863 13247 7921 13281
rect 7955 13247 8013 13281
rect 8047 13247 8105 13281
rect 8139 13247 8197 13281
rect 8231 13247 8289 13281
rect 8323 13247 8381 13281
rect 8415 13247 8473 13281
rect 8507 13247 8565 13281
rect 8599 13247 8657 13281
rect 8691 13247 8749 13281
rect 8783 13247 8841 13281
rect 8875 13247 8933 13281
rect 8967 13247 9025 13281
rect 9059 13247 9117 13281
rect 9151 13247 9209 13281
rect 9243 13247 9301 13281
rect 9335 13247 9393 13281
rect 9427 13247 9485 13281
rect 9519 13247 9577 13281
rect 9611 13247 9669 13281
rect 9703 13247 9761 13281
rect 9795 13247 9853 13281
rect 6351 13238 9861 13247
rect 9913 13238 9925 13290
rect 9977 13281 9989 13290
rect 10041 13281 10053 13290
rect 9979 13247 9989 13281
rect 9977 13238 9989 13247
rect 10041 13238 10053 13247
rect 10105 13238 10117 13290
rect 10169 13281 13679 13290
rect 13731 13281 13743 13290
rect 10169 13247 10221 13281
rect 10255 13247 10313 13281
rect 10347 13247 10405 13281
rect 10439 13247 10497 13281
rect 10531 13247 10589 13281
rect 10623 13247 10681 13281
rect 10715 13247 10773 13281
rect 10807 13247 10865 13281
rect 10899 13247 10957 13281
rect 10991 13247 11049 13281
rect 11083 13247 11141 13281
rect 11175 13247 11233 13281
rect 11267 13247 11325 13281
rect 11359 13247 11417 13281
rect 11451 13247 11509 13281
rect 11543 13247 11601 13281
rect 11635 13247 11693 13281
rect 11727 13247 11785 13281
rect 11819 13247 11877 13281
rect 11911 13247 11969 13281
rect 12003 13247 12061 13281
rect 12095 13247 12153 13281
rect 12187 13247 12245 13281
rect 12279 13247 12337 13281
rect 12371 13247 12429 13281
rect 12463 13247 12521 13281
rect 12555 13247 12613 13281
rect 12647 13247 12705 13281
rect 12739 13247 12797 13281
rect 12831 13247 12889 13281
rect 12923 13247 12981 13281
rect 13015 13247 13073 13281
rect 13107 13247 13165 13281
rect 13199 13247 13257 13281
rect 13291 13247 13349 13281
rect 13383 13247 13441 13281
rect 13475 13247 13533 13281
rect 13567 13247 13625 13281
rect 13659 13247 13679 13281
rect 10169 13238 13679 13247
rect 13731 13238 13743 13247
rect 13795 13238 13807 13290
rect 13859 13238 13871 13290
rect 13923 13281 13935 13290
rect 13923 13238 13935 13247
rect 13987 13281 17497 13290
rect 13987 13247 13993 13281
rect 14027 13247 14085 13281
rect 14119 13247 14177 13281
rect 14211 13247 14269 13281
rect 14303 13247 14361 13281
rect 14395 13247 14453 13281
rect 14487 13247 14545 13281
rect 14579 13247 14637 13281
rect 14671 13247 14729 13281
rect 14763 13247 14821 13281
rect 14855 13247 14913 13281
rect 14947 13247 15005 13281
rect 15039 13247 15097 13281
rect 15131 13247 15189 13281
rect 15223 13247 15281 13281
rect 15315 13247 15373 13281
rect 15407 13247 15465 13281
rect 15499 13247 15557 13281
rect 15591 13247 15649 13281
rect 15683 13247 15741 13281
rect 15775 13247 15833 13281
rect 15867 13247 15925 13281
rect 15959 13247 16017 13281
rect 16051 13247 16109 13281
rect 16143 13247 16201 13281
rect 16235 13247 16293 13281
rect 16327 13247 16385 13281
rect 16419 13247 16477 13281
rect 16511 13247 16569 13281
rect 16603 13247 16661 13281
rect 16695 13247 16753 13281
rect 16787 13247 16845 13281
rect 16879 13247 16937 13281
rect 16971 13247 17029 13281
rect 17063 13247 17121 13281
rect 17155 13247 17213 13281
rect 17247 13247 17305 13281
rect 17339 13247 17397 13281
rect 17431 13247 17489 13281
rect 13987 13238 17497 13247
rect 17549 13238 17561 13290
rect 17613 13281 17625 13290
rect 17677 13281 17689 13290
rect 17615 13247 17625 13281
rect 17613 13238 17625 13247
rect 17677 13238 17689 13247
rect 17741 13238 17753 13290
rect 17805 13281 20220 13290
rect 17805 13247 17857 13281
rect 17891 13247 17949 13281
rect 17983 13247 18041 13281
rect 18075 13247 18133 13281
rect 18167 13247 18225 13281
rect 18259 13247 18317 13281
rect 18351 13247 18409 13281
rect 18443 13247 18501 13281
rect 18535 13247 18593 13281
rect 18627 13247 18685 13281
rect 18719 13247 18777 13281
rect 18811 13247 18869 13281
rect 18903 13247 18961 13281
rect 18995 13247 19053 13281
rect 19087 13247 19145 13281
rect 19179 13247 19237 13281
rect 19271 13247 19329 13281
rect 19363 13247 19421 13281
rect 19455 13247 19513 13281
rect 19547 13247 19605 13281
rect 19639 13247 19697 13281
rect 19731 13247 19789 13281
rect 19823 13247 19881 13281
rect 19915 13247 19973 13281
rect 20007 13247 20065 13281
rect 20099 13247 20157 13281
rect 20191 13247 20220 13281
rect 17805 13238 20220 13247
rect 4948 13216 20220 13238
rect 10574 13136 10580 13188
rect 10632 13136 10638 13188
rect 11862 13136 11868 13188
rect 11920 13136 11926 13188
rect 14438 13176 14444 13188
rect 13996 13148 14444 13176
rect 9194 12932 9200 12984
rect 9252 12972 9258 12984
rect 10393 12975 10451 12981
rect 10393 12972 10405 12975
rect 9252 12944 10405 12972
rect 9252 12932 9258 12944
rect 10393 12941 10405 12944
rect 10439 12941 10451 12975
rect 10592 12972 10620 13136
rect 10689 13111 10747 13117
rect 10689 13077 10701 13111
rect 10735 13108 10747 13111
rect 10850 13108 10856 13120
rect 10735 13080 10856 13108
rect 10735 13077 10807 13080
rect 10689 13071 10807 13077
rect 10749 13048 10807 13071
rect 10850 13068 10856 13080
rect 10908 13108 10914 13120
rect 11337 13111 11467 13117
rect 11337 13108 11349 13111
rect 10908 13080 11349 13108
rect 10908 13068 10914 13080
rect 11337 13077 11349 13080
rect 11383 13077 11421 13111
rect 11455 13077 11467 13111
rect 11880 13108 11908 13136
rect 12965 13111 13095 13117
rect 11880 13080 12184 13108
rect 11337 13071 11467 13077
rect 12156 13049 12184 13080
rect 12965 13077 12977 13111
rect 13011 13077 13049 13111
rect 13083 13108 13095 13111
rect 13685 13111 13743 13117
rect 13685 13108 13697 13111
rect 13083 13080 13697 13108
rect 13083 13077 13095 13080
rect 12965 13071 13095 13077
rect 13625 13077 13697 13080
rect 13731 13108 13743 13111
rect 13996 13108 14024 13148
rect 14438 13136 14444 13148
rect 14496 13176 14502 13188
rect 14496 13148 15496 13176
rect 14496 13136 14502 13148
rect 13731 13080 14024 13108
rect 14533 13111 14591 13117
rect 13731 13077 13743 13080
rect 13625 13071 13743 13077
rect 14533 13077 14545 13111
rect 14579 13108 14591 13111
rect 14714 13108 14720 13120
rect 14579 13080 14720 13108
rect 14579 13077 14591 13080
rect 14533 13071 14591 13077
rect 10749 13014 10761 13048
rect 10795 13014 10807 13048
rect 10749 13008 10807 13014
rect 10965 13043 11023 13049
rect 10965 13009 10977 13043
rect 11011 13040 11023 13043
rect 11681 13043 11739 13049
rect 11681 13040 11693 13043
rect 11011 13012 11693 13040
rect 11011 13009 11023 13012
rect 10965 13003 11023 13009
rect 11681 13009 11693 13012
rect 11727 13040 11739 13043
rect 12048 13043 12106 13049
rect 12048 13040 12060 13043
rect 11727 13012 12060 13040
rect 11727 13009 11739 13012
rect 11681 13003 11739 13009
rect 12048 13009 12060 13012
rect 12094 13009 12106 13043
rect 12048 13003 12106 13009
rect 12141 13043 12199 13049
rect 12141 13009 12153 13043
rect 12187 13040 12199 13043
rect 12233 13043 12291 13049
rect 12233 13040 12245 13043
rect 12187 13012 12245 13040
rect 12187 13009 12199 13012
rect 12141 13003 12199 13009
rect 12233 13009 12245 13012
rect 12279 13009 12291 13043
rect 12233 13003 12291 13009
rect 12326 13043 12384 13049
rect 12326 13009 12338 13043
rect 12372 13040 12384 13043
rect 12693 13043 12751 13049
rect 12693 13040 12705 13043
rect 12372 13012 12705 13040
rect 12372 13009 12384 13012
rect 12326 13003 12384 13009
rect 12693 13009 12705 13012
rect 12739 13040 12751 13043
rect 13409 13043 13467 13049
rect 13409 13040 13421 13043
rect 12739 13012 13421 13040
rect 12739 13009 12751 13012
rect 12693 13003 12751 13009
rect 13409 13009 13421 13012
rect 13455 13009 13467 13043
rect 13409 13003 13467 13009
rect 13625 13048 13683 13071
rect 14714 13068 14720 13080
rect 14772 13068 14778 13120
rect 14806 13068 14812 13120
rect 14864 13068 14870 13120
rect 14990 13068 14996 13120
rect 15048 13068 15054 13120
rect 15381 13111 15439 13117
rect 15381 13077 15393 13111
rect 15427 13108 15439 13111
rect 15468 13108 15496 13148
rect 16278 13136 16284 13188
rect 16336 13136 16342 13188
rect 16925 13179 16983 13185
rect 16925 13145 16937 13179
rect 16971 13176 16983 13179
rect 17014 13176 17020 13188
rect 16971 13148 17020 13176
rect 16971 13145 16983 13148
rect 16925 13139 16983 13145
rect 17014 13136 17020 13148
rect 17072 13136 17078 13188
rect 16029 13111 16159 13117
rect 16029 13108 16041 13111
rect 15427 13080 16041 13108
rect 15427 13077 15499 13080
rect 15381 13071 15499 13077
rect 16029 13077 16041 13080
rect 16075 13077 16113 13111
rect 16147 13077 16159 13111
rect 16296 13108 16324 13136
rect 16296 13080 16876 13108
rect 16029 13071 16159 13077
rect 13625 13014 13637 13048
rect 13671 13014 13683 13048
rect 13625 13008 13683 13014
rect 14441 13043 14499 13049
rect 14441 13009 14453 13043
rect 14487 13009 14499 13043
rect 14441 13003 14499 13009
rect 11865 12975 11923 12981
rect 11865 12972 11877 12975
rect 10592 12944 11877 12972
rect 10393 12935 10451 12941
rect 11865 12941 11877 12944
rect 11911 12941 11923 12975
rect 11865 12935 11923 12941
rect 12506 12932 12512 12984
rect 12564 12932 12570 12984
rect 13058 12932 13064 12984
rect 13116 12972 13122 12984
rect 14456 12972 14484 13003
rect 13116 12944 14484 12972
rect 14717 12975 14775 12981
rect 13116 12932 13122 12944
rect 14717 12941 14729 12975
rect 14763 12972 14775 12975
rect 14824 12972 14852 13068
rect 14763 12944 14852 12972
rect 15008 12972 15036 13068
rect 15441 13048 15499 13071
rect 15441 13014 15453 13048
rect 15487 13040 15499 13048
rect 15542 13040 15548 13052
rect 15487 13014 15548 13040
rect 15441 13012 15548 13014
rect 15441 13008 15499 13012
rect 15542 13000 15548 13012
rect 15600 13000 15606 13052
rect 16848 13049 16876 13080
rect 15657 13043 15715 13049
rect 15657 13009 15669 13043
rect 15703 13040 15715 13043
rect 16373 13043 16431 13049
rect 16373 13040 16385 13043
rect 15703 13012 16385 13040
rect 15703 13009 15715 13012
rect 15657 13003 15715 13009
rect 16373 13009 16385 13012
rect 16419 13040 16431 13043
rect 16740 13043 16798 13049
rect 16740 13040 16752 13043
rect 16419 13012 16752 13040
rect 16419 13009 16431 13012
rect 16373 13003 16431 13009
rect 16740 13009 16752 13012
rect 16786 13009 16798 13043
rect 16740 13003 16798 13009
rect 16833 13043 16891 13049
rect 16833 13009 16845 13043
rect 16879 13009 16891 13043
rect 16833 13003 16891 13009
rect 16557 12975 16615 12981
rect 16557 12972 16569 12975
rect 15008 12944 16569 12972
rect 14763 12941 14775 12944
rect 14717 12935 14775 12941
rect 16557 12941 16569 12944
rect 16603 12941 16615 12975
rect 16557 12935 16615 12941
rect 17566 12932 17572 12984
rect 17624 12932 17630 12984
rect 10965 12907 11023 12913
rect 10965 12873 10977 12907
rect 11011 12904 11023 12907
rect 11589 12907 11647 12913
rect 11589 12904 11601 12907
rect 11011 12876 11601 12904
rect 11011 12873 11023 12876
rect 10965 12867 11023 12873
rect 11589 12873 11601 12876
rect 11635 12904 11647 12907
rect 11967 12907 12025 12913
rect 11967 12904 11979 12907
rect 11635 12876 11979 12904
rect 11635 12873 11647 12876
rect 11589 12867 11647 12873
rect 11967 12873 11979 12876
rect 12013 12873 12025 12907
rect 11967 12867 12025 12873
rect 12407 12907 12465 12913
rect 12407 12873 12419 12907
rect 12453 12904 12465 12907
rect 12785 12907 12843 12913
rect 12785 12904 12797 12907
rect 12453 12876 12797 12904
rect 12453 12873 12465 12876
rect 12407 12867 12465 12873
rect 12785 12873 12797 12876
rect 12831 12904 12843 12907
rect 13409 12907 13467 12913
rect 13409 12904 13421 12907
rect 12831 12876 13421 12904
rect 12831 12873 12843 12876
rect 12785 12867 12843 12873
rect 13409 12873 13421 12876
rect 13455 12873 13467 12907
rect 13409 12867 13467 12873
rect 14073 12907 14131 12913
rect 14073 12873 14085 12907
rect 14119 12904 14131 12907
rect 14254 12904 14260 12916
rect 14119 12876 14260 12904
rect 14119 12873 14131 12876
rect 14073 12867 14131 12873
rect 14254 12864 14260 12876
rect 14312 12864 14318 12916
rect 15657 12907 15715 12913
rect 15657 12873 15669 12907
rect 15703 12904 15715 12907
rect 16281 12907 16339 12913
rect 16281 12904 16293 12907
rect 15703 12876 16293 12904
rect 15703 12873 15715 12876
rect 15657 12867 15715 12873
rect 16281 12873 16293 12876
rect 16327 12904 16339 12907
rect 16659 12907 16717 12913
rect 16659 12904 16671 12907
rect 16327 12876 16671 12904
rect 16327 12873 16339 12876
rect 16281 12867 16339 12873
rect 16659 12873 16671 12876
rect 16705 12873 16717 12907
rect 16659 12867 16717 12873
rect 9746 12796 9752 12848
rect 9804 12796 9810 12848
rect 10206 12796 10212 12848
rect 10264 12836 10270 12848
rect 11494 12836 11500 12848
rect 10264 12808 11500 12836
rect 10264 12796 10270 12808
rect 11494 12796 11500 12808
rect 11552 12796 11558 12848
rect 12874 12796 12880 12848
rect 12932 12836 12938 12848
rect 13981 12839 14039 12845
rect 13981 12836 13993 12839
rect 12932 12808 13993 12836
rect 12932 12796 12938 12808
rect 13981 12805 13993 12808
rect 14027 12805 14039 12839
rect 13981 12799 14039 12805
rect 14162 12796 14168 12848
rect 14220 12836 14226 12848
rect 15085 12839 15143 12845
rect 15085 12836 15097 12839
rect 14220 12808 15097 12836
rect 14220 12796 14226 12808
rect 15085 12805 15097 12808
rect 15131 12805 15143 12839
rect 15085 12799 15143 12805
rect 4948 12746 20220 12768
rect 4948 12737 6703 12746
rect 6755 12737 6767 12746
rect 6819 12737 6831 12746
rect 4948 12703 4977 12737
rect 5011 12703 5069 12737
rect 5103 12703 5161 12737
rect 5195 12703 5253 12737
rect 5287 12703 5345 12737
rect 5379 12703 5437 12737
rect 5471 12703 5529 12737
rect 5563 12703 5621 12737
rect 5655 12703 5713 12737
rect 5747 12703 5805 12737
rect 5839 12703 5897 12737
rect 5931 12703 5989 12737
rect 6023 12703 6081 12737
rect 6115 12703 6173 12737
rect 6207 12703 6265 12737
rect 6299 12703 6357 12737
rect 6391 12703 6449 12737
rect 6483 12703 6541 12737
rect 6575 12703 6633 12737
rect 6667 12703 6703 12737
rect 6759 12703 6767 12737
rect 4948 12694 6703 12703
rect 6755 12694 6767 12703
rect 6819 12694 6831 12703
rect 6883 12694 6895 12746
rect 6947 12694 6959 12746
rect 7011 12737 10521 12746
rect 7035 12703 7093 12737
rect 7127 12703 7185 12737
rect 7219 12703 7277 12737
rect 7311 12703 7369 12737
rect 7403 12703 7461 12737
rect 7495 12703 7553 12737
rect 7587 12703 7645 12737
rect 7679 12703 7737 12737
rect 7771 12703 7829 12737
rect 7863 12703 7921 12737
rect 7955 12703 8013 12737
rect 8047 12703 8105 12737
rect 8139 12703 8197 12737
rect 8231 12703 8289 12737
rect 8323 12703 8381 12737
rect 8415 12703 8473 12737
rect 8507 12703 8565 12737
rect 8599 12703 8657 12737
rect 8691 12703 8749 12737
rect 8783 12703 8841 12737
rect 8875 12703 8933 12737
rect 8967 12703 9025 12737
rect 9059 12703 9117 12737
rect 9151 12703 9209 12737
rect 9243 12703 9301 12737
rect 9335 12703 9393 12737
rect 9427 12703 9485 12737
rect 9519 12703 9577 12737
rect 9611 12703 9669 12737
rect 9703 12703 9761 12737
rect 9795 12703 9853 12737
rect 9887 12703 9945 12737
rect 9979 12703 10037 12737
rect 10071 12703 10129 12737
rect 10163 12703 10221 12737
rect 10255 12703 10313 12737
rect 10347 12703 10405 12737
rect 10439 12703 10497 12737
rect 7011 12694 10521 12703
rect 10573 12694 10585 12746
rect 10637 12694 10649 12746
rect 10701 12737 10713 12746
rect 10765 12737 10777 12746
rect 10829 12737 14339 12746
rect 14391 12737 14403 12746
rect 14455 12737 14467 12746
rect 10765 12703 10773 12737
rect 10829 12703 10865 12737
rect 10899 12703 10957 12737
rect 10991 12703 11049 12737
rect 11083 12703 11141 12737
rect 11175 12703 11233 12737
rect 11267 12703 11325 12737
rect 11359 12703 11417 12737
rect 11451 12703 11509 12737
rect 11543 12703 11601 12737
rect 11635 12703 11693 12737
rect 11727 12703 11785 12737
rect 11819 12703 11877 12737
rect 11911 12703 11969 12737
rect 12003 12703 12061 12737
rect 12095 12703 12153 12737
rect 12187 12703 12245 12737
rect 12279 12703 12337 12737
rect 12371 12703 12429 12737
rect 12463 12703 12521 12737
rect 12555 12703 12613 12737
rect 12647 12703 12705 12737
rect 12739 12703 12797 12737
rect 12831 12703 12889 12737
rect 12923 12703 12981 12737
rect 13015 12703 13073 12737
rect 13107 12703 13165 12737
rect 13199 12703 13257 12737
rect 13291 12703 13349 12737
rect 13383 12703 13441 12737
rect 13475 12703 13533 12737
rect 13567 12703 13625 12737
rect 13659 12703 13717 12737
rect 13751 12703 13809 12737
rect 13843 12703 13901 12737
rect 13935 12703 13993 12737
rect 14027 12703 14085 12737
rect 14119 12703 14177 12737
rect 14211 12703 14269 12737
rect 14303 12703 14339 12737
rect 14395 12703 14403 12737
rect 10701 12694 10713 12703
rect 10765 12694 10777 12703
rect 10829 12694 14339 12703
rect 14391 12694 14403 12703
rect 14455 12694 14467 12703
rect 14519 12694 14531 12746
rect 14583 12694 14595 12746
rect 14647 12737 18157 12746
rect 14671 12703 14729 12737
rect 14763 12703 14821 12737
rect 14855 12703 14913 12737
rect 14947 12703 15005 12737
rect 15039 12703 15097 12737
rect 15131 12703 15189 12737
rect 15223 12703 15281 12737
rect 15315 12703 15373 12737
rect 15407 12703 15465 12737
rect 15499 12703 15557 12737
rect 15591 12703 15649 12737
rect 15683 12703 15741 12737
rect 15775 12703 15833 12737
rect 15867 12703 15925 12737
rect 15959 12703 16017 12737
rect 16051 12703 16109 12737
rect 16143 12703 16201 12737
rect 16235 12703 16293 12737
rect 16327 12703 16385 12737
rect 16419 12703 16477 12737
rect 16511 12703 16569 12737
rect 16603 12703 16661 12737
rect 16695 12703 16753 12737
rect 16787 12703 16845 12737
rect 16879 12703 16937 12737
rect 16971 12703 17029 12737
rect 17063 12703 17121 12737
rect 17155 12703 17213 12737
rect 17247 12703 17305 12737
rect 17339 12703 17397 12737
rect 17431 12703 17489 12737
rect 17523 12703 17581 12737
rect 17615 12703 17673 12737
rect 17707 12703 17765 12737
rect 17799 12703 17857 12737
rect 17891 12703 17949 12737
rect 17983 12703 18041 12737
rect 18075 12703 18133 12737
rect 14647 12694 18157 12703
rect 18209 12694 18221 12746
rect 18273 12694 18285 12746
rect 18337 12737 18349 12746
rect 18401 12737 18413 12746
rect 18465 12737 20220 12746
rect 18401 12703 18409 12737
rect 18465 12703 18501 12737
rect 18535 12703 18593 12737
rect 18627 12703 18685 12737
rect 18719 12703 18777 12737
rect 18811 12703 18869 12737
rect 18903 12703 18961 12737
rect 18995 12703 19053 12737
rect 19087 12703 19145 12737
rect 19179 12703 19237 12737
rect 19271 12703 19329 12737
rect 19363 12703 19421 12737
rect 19455 12703 19513 12737
rect 19547 12703 19605 12737
rect 19639 12703 19697 12737
rect 19731 12703 19789 12737
rect 19823 12703 19881 12737
rect 19915 12703 19973 12737
rect 20007 12703 20065 12737
rect 20099 12703 20157 12737
rect 20191 12703 20220 12737
rect 18337 12694 18349 12703
rect 18401 12694 18413 12703
rect 18465 12694 20220 12703
rect 4948 12672 20220 12694
rect 9654 12592 9660 12644
rect 9712 12592 9718 12644
rect 10206 12592 10212 12644
rect 10264 12592 10270 12644
rect 12141 12635 12199 12641
rect 12141 12601 12153 12635
rect 12187 12632 12199 12635
rect 12690 12632 12696 12644
rect 12187 12604 12696 12632
rect 12187 12601 12199 12604
rect 12141 12595 12199 12601
rect 12690 12592 12696 12604
rect 12748 12592 12754 12644
rect 13981 12635 14039 12641
rect 13981 12601 13993 12635
rect 14027 12632 14039 12635
rect 14070 12632 14076 12644
rect 14027 12604 14076 12632
rect 14027 12601 14039 12604
rect 13981 12595 14039 12601
rect 14070 12592 14076 12604
rect 14128 12592 14134 12644
rect 14714 12592 14720 12644
rect 14772 12592 14778 12644
rect 9672 12564 9700 12592
rect 10485 12567 10543 12573
rect 10485 12564 10497 12567
rect 9672 12536 10497 12564
rect 10485 12533 10497 12536
rect 10531 12533 10543 12567
rect 10485 12527 10543 12533
rect 15259 12567 15317 12573
rect 15259 12533 15271 12567
rect 15305 12564 15317 12567
rect 15637 12567 15695 12573
rect 15637 12564 15649 12567
rect 15305 12536 15649 12564
rect 15305 12533 15317 12536
rect 15259 12527 15317 12533
rect 15637 12533 15649 12536
rect 15683 12564 15695 12567
rect 16261 12567 16319 12573
rect 16261 12564 16273 12567
rect 15683 12536 16273 12564
rect 15683 12533 15695 12536
rect 15637 12527 15695 12533
rect 16261 12533 16273 12536
rect 16307 12533 16319 12567
rect 16261 12527 16319 12533
rect 9746 12456 9752 12508
rect 9804 12496 9810 12508
rect 10945 12499 11003 12505
rect 10945 12496 10957 12499
rect 9804 12468 10957 12496
rect 9804 12456 9810 12468
rect 10945 12465 10957 12468
rect 10991 12465 11003 12499
rect 10945 12459 11003 12465
rect 11129 12499 11187 12505
rect 11129 12465 11141 12499
rect 11175 12496 11187 12499
rect 11589 12499 11647 12505
rect 11589 12496 11601 12499
rect 11175 12468 11601 12496
rect 11175 12465 11187 12468
rect 11129 12459 11187 12465
rect 11589 12465 11601 12468
rect 11635 12496 11647 12499
rect 11678 12496 11684 12508
rect 11635 12468 11684 12496
rect 11635 12465 11647 12468
rect 11589 12459 11647 12465
rect 5238 12388 5244 12440
rect 5296 12388 5302 12440
rect 9194 12388 9200 12440
rect 9252 12388 9258 12440
rect 10114 12428 10120 12440
rect 9764 12400 10120 12428
rect 7081 12363 7139 12369
rect 7081 12329 7093 12363
rect 7127 12360 7139 12363
rect 9764 12360 9792 12400
rect 10114 12388 10120 12400
rect 10172 12428 10178 12440
rect 10853 12431 10911 12437
rect 10853 12428 10865 12431
rect 10172 12400 10865 12428
rect 10172 12388 10178 12400
rect 10853 12397 10865 12400
rect 10899 12397 10911 12431
rect 10960 12428 10988 12459
rect 11678 12456 11684 12468
rect 11736 12456 11742 12508
rect 14162 12496 14168 12508
rect 13076 12468 14168 12496
rect 13076 12437 13104 12468
rect 14162 12456 14168 12468
rect 14220 12456 14226 12508
rect 15082 12456 15088 12508
rect 15140 12456 15146 12508
rect 15361 12499 15419 12505
rect 15361 12465 15373 12499
rect 15407 12496 15419 12499
rect 15726 12496 15732 12508
rect 15407 12468 15732 12496
rect 15407 12465 15419 12468
rect 15361 12459 15419 12465
rect 15726 12456 15732 12468
rect 15784 12456 15790 12508
rect 16833 12499 16891 12505
rect 16833 12465 16845 12499
rect 16879 12496 16891 12499
rect 16879 12468 17612 12496
rect 16879 12465 16891 12468
rect 16833 12459 16891 12465
rect 17584 12440 17612 12468
rect 11773 12431 11831 12437
rect 11773 12428 11785 12431
rect 10960 12400 11785 12428
rect 10853 12391 10911 12397
rect 11773 12397 11785 12400
rect 11819 12397 11831 12431
rect 11773 12391 11831 12397
rect 13061 12431 13119 12437
rect 13061 12397 13073 12431
rect 13107 12397 13119 12431
rect 13061 12391 13119 12397
rect 13150 12388 13156 12440
rect 13208 12428 13214 12440
rect 13337 12431 13395 12437
rect 13337 12428 13349 12431
rect 13208 12400 13349 12428
rect 13208 12388 13214 12400
rect 13337 12397 13349 12400
rect 13383 12397 13395 12431
rect 13337 12391 13395 12397
rect 13426 12388 13432 12440
rect 13484 12428 13490 12440
rect 13797 12431 13855 12437
rect 13797 12428 13809 12431
rect 13484 12400 13809 12428
rect 13484 12388 13490 12400
rect 13797 12397 13809 12400
rect 13843 12397 13855 12431
rect 13797 12391 13855 12397
rect 15178 12431 15236 12437
rect 15178 12397 15190 12431
rect 15224 12428 15236 12431
rect 15545 12431 15603 12437
rect 15545 12428 15557 12431
rect 15224 12400 15557 12428
rect 15224 12397 15236 12400
rect 15178 12391 15236 12397
rect 15545 12397 15557 12400
rect 15591 12428 15603 12431
rect 16261 12431 16319 12437
rect 16261 12428 16273 12431
rect 15591 12400 16273 12428
rect 15591 12397 15603 12400
rect 15545 12391 15603 12397
rect 16261 12397 16273 12400
rect 16307 12397 16319 12431
rect 16261 12391 16319 12397
rect 16477 12426 16535 12432
rect 16477 12392 16489 12426
rect 16523 12392 16535 12426
rect 7127 12332 9792 12360
rect 10301 12363 10359 12369
rect 7127 12329 7139 12332
rect 7081 12323 7139 12329
rect 10301 12329 10313 12363
rect 10347 12360 10359 12363
rect 15634 12360 15640 12372
rect 10347 12332 11724 12360
rect 10347 12329 10359 12332
rect 10301 12323 10359 12329
rect 6989 12295 7047 12301
rect 6989 12261 7001 12295
rect 7035 12292 7047 12295
rect 7262 12292 7268 12304
rect 7035 12264 7268 12292
rect 7035 12261 7047 12264
rect 6989 12255 7047 12261
rect 7262 12252 7268 12264
rect 7320 12252 7326 12304
rect 9105 12295 9163 12301
rect 9105 12261 9117 12295
rect 9151 12292 9163 12295
rect 9378 12292 9384 12304
rect 9151 12264 9384 12292
rect 9151 12261 9163 12264
rect 9105 12255 9163 12261
rect 9378 12252 9384 12264
rect 9436 12252 9442 12304
rect 11696 12301 11724 12332
rect 13536 12332 15640 12360
rect 11681 12295 11739 12301
rect 11681 12261 11693 12295
rect 11727 12292 11739 12295
rect 12874 12292 12880 12304
rect 11727 12264 12880 12292
rect 11727 12261 11739 12264
rect 11681 12255 11739 12261
rect 12874 12252 12880 12264
rect 12932 12252 12938 12304
rect 12969 12295 13027 12301
rect 12969 12261 12981 12295
rect 13015 12292 13027 12295
rect 13536 12292 13564 12332
rect 15634 12320 15640 12332
rect 15692 12320 15698 12372
rect 16477 12369 16535 12392
rect 16922 12388 16928 12440
rect 16980 12428 16986 12440
rect 17109 12431 17167 12437
rect 17109 12428 17121 12431
rect 16980 12400 17121 12428
rect 16980 12388 16986 12400
rect 17109 12397 17121 12400
rect 17155 12397 17167 12431
rect 17109 12391 17167 12397
rect 17566 12388 17572 12440
rect 17624 12428 17630 12440
rect 19501 12431 19559 12437
rect 19501 12428 19513 12431
rect 17624 12400 19513 12428
rect 17624 12388 17630 12400
rect 19501 12397 19513 12400
rect 19547 12397 19559 12431
rect 19501 12391 19559 12397
rect 15817 12363 15947 12369
rect 15817 12360 15829 12363
rect 15744 12332 15829 12360
rect 13015 12264 13564 12292
rect 13015 12261 13027 12264
rect 12969 12255 13027 12261
rect 13610 12252 13616 12304
rect 13668 12252 13674 12304
rect 15542 12252 15548 12304
rect 15600 12292 15606 12304
rect 15744 12292 15772 12332
rect 15817 12329 15829 12332
rect 15863 12329 15901 12363
rect 15935 12360 15947 12363
rect 16477 12363 16595 12369
rect 16477 12360 16549 12363
rect 15935 12332 16549 12360
rect 15935 12329 15947 12332
rect 15817 12323 15947 12329
rect 16537 12329 16549 12332
rect 16583 12329 16595 12363
rect 16537 12323 16595 12329
rect 17477 12363 17535 12369
rect 17477 12329 17489 12363
rect 17523 12360 17535 12363
rect 17842 12360 17848 12372
rect 17523 12332 17848 12360
rect 17523 12329 17535 12332
rect 17477 12323 17535 12329
rect 17842 12320 17848 12332
rect 17900 12320 17906 12372
rect 19869 12363 19927 12369
rect 19869 12329 19881 12363
rect 19915 12360 19927 12363
rect 19958 12360 19964 12372
rect 19915 12332 19964 12360
rect 19915 12329 19927 12332
rect 19869 12323 19927 12329
rect 19958 12320 19964 12332
rect 20016 12320 20022 12372
rect 15600 12264 15772 12292
rect 15600 12252 15606 12264
rect 4948 12202 20220 12224
rect 4948 12193 6043 12202
rect 6095 12193 6107 12202
rect 4948 12159 4977 12193
rect 5011 12159 5069 12193
rect 5103 12159 5161 12193
rect 5195 12159 5253 12193
rect 5287 12159 5345 12193
rect 5379 12159 5437 12193
rect 5471 12159 5529 12193
rect 5563 12159 5621 12193
rect 5655 12159 5713 12193
rect 5747 12159 5805 12193
rect 5839 12159 5897 12193
rect 5931 12159 5989 12193
rect 6023 12159 6043 12193
rect 4948 12150 6043 12159
rect 6095 12150 6107 12159
rect 6159 12150 6171 12202
rect 6223 12150 6235 12202
rect 6287 12193 6299 12202
rect 6287 12150 6299 12159
rect 6351 12193 9861 12202
rect 6351 12159 6357 12193
rect 6391 12159 6449 12193
rect 6483 12159 6541 12193
rect 6575 12159 6633 12193
rect 6667 12159 6725 12193
rect 6759 12159 6817 12193
rect 6851 12159 6909 12193
rect 6943 12159 7001 12193
rect 7035 12159 7093 12193
rect 7127 12159 7185 12193
rect 7219 12159 7277 12193
rect 7311 12159 7369 12193
rect 7403 12159 7461 12193
rect 7495 12159 7553 12193
rect 7587 12159 7645 12193
rect 7679 12159 7737 12193
rect 7771 12159 7829 12193
rect 7863 12159 7921 12193
rect 7955 12159 8013 12193
rect 8047 12159 8105 12193
rect 8139 12159 8197 12193
rect 8231 12159 8289 12193
rect 8323 12159 8381 12193
rect 8415 12159 8473 12193
rect 8507 12159 8565 12193
rect 8599 12159 8657 12193
rect 8691 12159 8749 12193
rect 8783 12159 8841 12193
rect 8875 12159 8933 12193
rect 8967 12159 9025 12193
rect 9059 12159 9117 12193
rect 9151 12159 9209 12193
rect 9243 12159 9301 12193
rect 9335 12159 9393 12193
rect 9427 12159 9485 12193
rect 9519 12159 9577 12193
rect 9611 12159 9669 12193
rect 9703 12159 9761 12193
rect 9795 12159 9853 12193
rect 6351 12150 9861 12159
rect 9913 12150 9925 12202
rect 9977 12193 9989 12202
rect 10041 12193 10053 12202
rect 9979 12159 9989 12193
rect 9977 12150 9989 12159
rect 10041 12150 10053 12159
rect 10105 12150 10117 12202
rect 10169 12193 13679 12202
rect 13731 12193 13743 12202
rect 10169 12159 10221 12193
rect 10255 12159 10313 12193
rect 10347 12159 10405 12193
rect 10439 12159 10497 12193
rect 10531 12159 10589 12193
rect 10623 12159 10681 12193
rect 10715 12159 10773 12193
rect 10807 12159 10865 12193
rect 10899 12159 10957 12193
rect 10991 12159 11049 12193
rect 11083 12159 11141 12193
rect 11175 12159 11233 12193
rect 11267 12159 11325 12193
rect 11359 12159 11417 12193
rect 11451 12159 11509 12193
rect 11543 12159 11601 12193
rect 11635 12159 11693 12193
rect 11727 12159 11785 12193
rect 11819 12159 11877 12193
rect 11911 12159 11969 12193
rect 12003 12159 12061 12193
rect 12095 12159 12153 12193
rect 12187 12159 12245 12193
rect 12279 12159 12337 12193
rect 12371 12159 12429 12193
rect 12463 12159 12521 12193
rect 12555 12159 12613 12193
rect 12647 12159 12705 12193
rect 12739 12159 12797 12193
rect 12831 12159 12889 12193
rect 12923 12159 12981 12193
rect 13015 12159 13073 12193
rect 13107 12159 13165 12193
rect 13199 12159 13257 12193
rect 13291 12159 13349 12193
rect 13383 12159 13441 12193
rect 13475 12159 13533 12193
rect 13567 12159 13625 12193
rect 13659 12159 13679 12193
rect 10169 12150 13679 12159
rect 13731 12150 13743 12159
rect 13795 12150 13807 12202
rect 13859 12150 13871 12202
rect 13923 12193 13935 12202
rect 13923 12150 13935 12159
rect 13987 12193 17497 12202
rect 13987 12159 13993 12193
rect 14027 12159 14085 12193
rect 14119 12159 14177 12193
rect 14211 12159 14269 12193
rect 14303 12159 14361 12193
rect 14395 12159 14453 12193
rect 14487 12159 14545 12193
rect 14579 12159 14637 12193
rect 14671 12159 14729 12193
rect 14763 12159 14821 12193
rect 14855 12159 14913 12193
rect 14947 12159 15005 12193
rect 15039 12159 15097 12193
rect 15131 12159 15189 12193
rect 15223 12159 15281 12193
rect 15315 12159 15373 12193
rect 15407 12159 15465 12193
rect 15499 12159 15557 12193
rect 15591 12159 15649 12193
rect 15683 12159 15741 12193
rect 15775 12159 15833 12193
rect 15867 12159 15925 12193
rect 15959 12159 16017 12193
rect 16051 12159 16109 12193
rect 16143 12159 16201 12193
rect 16235 12159 16293 12193
rect 16327 12159 16385 12193
rect 16419 12159 16477 12193
rect 16511 12159 16569 12193
rect 16603 12159 16661 12193
rect 16695 12159 16753 12193
rect 16787 12159 16845 12193
rect 16879 12159 16937 12193
rect 16971 12159 17029 12193
rect 17063 12159 17121 12193
rect 17155 12159 17213 12193
rect 17247 12159 17305 12193
rect 17339 12159 17397 12193
rect 17431 12159 17489 12193
rect 13987 12150 17497 12159
rect 17549 12150 17561 12202
rect 17613 12193 17625 12202
rect 17677 12193 17689 12202
rect 17615 12159 17625 12193
rect 17613 12150 17625 12159
rect 17677 12150 17689 12159
rect 17741 12150 17753 12202
rect 17805 12193 20220 12202
rect 17805 12159 17857 12193
rect 17891 12159 17949 12193
rect 17983 12159 18041 12193
rect 18075 12159 18133 12193
rect 18167 12159 18225 12193
rect 18259 12159 18317 12193
rect 18351 12159 18409 12193
rect 18443 12159 18501 12193
rect 18535 12159 18593 12193
rect 18627 12159 18685 12193
rect 18719 12159 18777 12193
rect 18811 12159 18869 12193
rect 18903 12159 18961 12193
rect 18995 12159 19053 12193
rect 19087 12159 19145 12193
rect 19179 12159 19237 12193
rect 19271 12159 19329 12193
rect 19363 12159 19421 12193
rect 19455 12159 19513 12193
rect 19547 12159 19605 12193
rect 19639 12159 19697 12193
rect 19731 12159 19789 12193
rect 19823 12159 19881 12193
rect 19915 12159 19973 12193
rect 20007 12159 20065 12193
rect 20099 12159 20157 12193
rect 20191 12159 20220 12193
rect 17805 12150 20220 12159
rect 4948 12128 20220 12150
rect 750 10160 5300 10200
rect 750 10020 5160 10160
rect 5260 10020 5300 10160
rect 750 10000 5300 10020
rect 7200 10150 7400 10200
rect -200 3630 620 3640
rect -200 3450 430 3630
rect 610 3450 620 3630
rect -200 3440 620 3450
rect -200 2690 0 2700
rect 200 2690 680 2700
rect -200 2510 440 2690
rect 620 2510 680 2690
rect -200 2500 680 2510
rect 750 2060 950 10000
rect 7200 9980 7240 10150
rect 7370 9980 7400 10150
rect 7200 9700 7400 9980
rect 4030 9500 7400 9700
rect 9300 10190 9500 10300
rect 9300 10020 9340 10190
rect 9470 10020 9500 10190
rect 3400 6720 3700 6750
rect 3400 6480 3430 6720
rect 3650 6480 3700 6720
rect 3400 5852 3700 6480
rect 3400 5650 3532 5852
rect 3526 5455 3532 5650
rect 3570 5650 3700 5852
rect 3570 5455 3576 5650
rect 3526 5443 3576 5455
rect 3526 5221 3576 5233
rect 3526 4940 3532 5221
rect 3450 4824 3532 4940
rect 3570 4940 3576 5221
rect 3570 4824 3650 4940
rect 1470 4311 1530 4330
rect 1470 4310 1482 4311
rect 1450 4277 1482 4310
rect 1516 4310 1530 4311
rect 1516 4277 1570 4310
rect 1450 4213 1570 4277
rect 1432 4201 1570 4213
rect 1432 3713 1438 4201
rect 1472 4180 1526 4201
rect 1472 3713 1478 4180
rect 1432 3701 1478 3713
rect 1520 3713 1526 4180
rect 1560 4180 1570 4201
rect 1760 4304 3010 4330
rect 1760 4270 1995 4304
rect 2029 4270 2187 4304
rect 2221 4270 2379 4304
rect 2413 4270 2571 4304
rect 2605 4270 2763 4304
rect 2797 4270 2955 4304
rect 2989 4270 3010 4304
rect 3170 4311 3230 4330
rect 3170 4277 3182 4311
rect 3216 4277 3230 4311
rect 3170 4270 3230 4277
rect 1560 3820 1566 4180
rect 1670 3911 1730 3930
rect 1670 3877 1682 3911
rect 1716 3877 1730 3911
rect 1670 3870 1730 3877
rect 1760 3830 1800 4270
rect 1983 4264 2041 4270
rect 2175 4264 2233 4270
rect 2367 4264 2425 4270
rect 2559 4264 2617 4270
rect 2751 4264 2809 4270
rect 2943 4264 3001 4270
rect 3132 4218 3178 4230
rect 1632 3820 1678 3830
rect 1560 3818 1678 3820
rect 1560 3713 1638 3818
rect 1040 3620 1260 3640
rect 1040 3440 1050 3620
rect 1230 3590 1260 3620
rect 1520 3590 1638 3713
rect 1230 3580 1638 3590
rect 1230 3490 1310 3580
rect 1360 3490 1638 3580
rect 1230 3480 1638 3490
rect 1230 3440 1260 3480
rect 1040 3430 1240 3440
rect 1520 3250 1638 3480
rect 1632 3242 1638 3250
rect 1672 3242 1678 3818
rect 1632 3230 1678 3242
rect 1720 3818 1800 3830
rect 1720 3242 1726 3818
rect 1760 3720 1800 3818
rect 1845 4200 1891 4206
rect 2037 4200 2083 4206
rect 2229 4200 2275 4206
rect 2421 4200 2467 4206
rect 2613 4200 2659 4206
rect 2805 4200 2851 4206
rect 2997 4200 3043 4206
rect 1845 4194 3043 4200
rect 1760 3380 1766 3720
rect 1845 3706 1851 4194
rect 1885 4050 2043 4194
rect 1885 3950 1890 4050
rect 2030 3950 2043 4050
rect 1885 3820 2043 3950
rect 1885 3706 1891 3820
rect 1845 3694 1891 3706
rect 1941 3740 1987 3752
rect 1941 3550 1947 3740
rect 1760 3242 1790 3380
rect 1930 3270 1947 3550
rect 1720 3230 1790 3242
rect 1941 3252 1947 3270
rect 1981 3550 1987 3740
rect 2037 3706 2043 3820
rect 2077 3820 2235 4194
rect 2077 3706 2083 3820
rect 2037 3694 2083 3706
rect 2133 3740 2179 3752
rect 2133 3550 2139 3740
rect 1981 3270 2139 3550
rect 1981 3252 1987 3270
rect 1941 3240 1987 3252
rect 2133 3252 2139 3270
rect 2173 3550 2179 3740
rect 2229 3706 2235 3820
rect 2269 3820 2427 4194
rect 2269 3706 2275 3820
rect 2229 3694 2275 3706
rect 2325 3740 2371 3752
rect 2325 3550 2331 3740
rect 2173 3270 2331 3550
rect 2173 3252 2179 3270
rect 2133 3240 2179 3252
rect 2325 3252 2331 3270
rect 2365 3550 2371 3740
rect 2421 3706 2427 3820
rect 2461 3820 2619 4194
rect 2461 3706 2467 3820
rect 2421 3694 2467 3706
rect 2517 3740 2563 3752
rect 2517 3550 2523 3740
rect 2365 3270 2523 3550
rect 2365 3252 2371 3270
rect 2325 3240 2371 3252
rect 2517 3252 2523 3270
rect 2557 3550 2563 3740
rect 2613 3706 2619 3820
rect 2653 3820 2811 4194
rect 2653 3706 2659 3820
rect 2613 3694 2659 3706
rect 2709 3740 2755 3752
rect 2709 3550 2715 3740
rect 2557 3270 2715 3550
rect 2557 3252 2563 3270
rect 2517 3240 2563 3252
rect 2709 3252 2715 3270
rect 2749 3550 2755 3740
rect 2805 3706 2811 3820
rect 2845 3820 3003 4194
rect 2845 3706 2851 3820
rect 2805 3694 2851 3706
rect 2901 3740 2947 3752
rect 2901 3550 2907 3740
rect 2749 3270 2907 3550
rect 2749 3252 2755 3270
rect 2709 3240 2755 3252
rect 2901 3252 2907 3270
rect 2941 3550 2947 3740
rect 2997 3706 3003 3820
rect 3037 3706 3043 4194
rect 2997 3694 3043 3706
rect 2941 3340 3080 3550
rect 3132 3340 3138 4218
rect 2941 3270 3138 3340
rect 2941 3252 2947 3270
rect 2980 3260 3138 3270
rect 2901 3240 2947 3252
rect 3050 3242 3138 3260
rect 3172 3340 3178 4218
rect 3220 4218 3266 4230
rect 3220 3340 3226 4218
rect 3172 3242 3226 3340
rect 3260 3340 3266 4218
rect 3260 3242 3290 3340
rect 1450 3183 1530 3190
rect 1450 3149 1482 3183
rect 1516 3149 1530 3183
rect 1450 3130 1530 3149
rect 1670 3183 1730 3190
rect 1670 3149 1682 3183
rect 1716 3149 1730 3183
rect 1440 2780 1560 2800
rect 1440 2746 1486 2780
rect 1520 2746 1560 2780
rect 1040 2690 1260 2700
rect 1440 2691 1560 2746
rect 1670 2786 1730 3149
rect 1670 2780 1732 2786
rect 1670 2746 1686 2780
rect 1720 2746 1732 2780
rect 1670 2740 1732 2746
rect 1760 2708 1790 3230
rect 1900 3182 2910 3190
rect 1887 3176 2910 3182
rect 1887 3142 1899 3176
rect 1933 3142 2091 3176
rect 2125 3142 2283 3176
rect 2317 3142 2475 3176
rect 2509 3142 2667 3176
rect 2701 3142 2859 3176
rect 2893 3142 2910 3176
rect 1887 3136 2910 3142
rect 1900 3130 2910 3136
rect 3050 3183 3290 3242
rect 3050 3149 3182 3183
rect 3216 3149 3290 3183
rect 3050 3100 3290 3149
rect 3450 3100 3650 4824
rect 3050 3000 3650 3100
rect 1990 2779 3010 2800
rect 1987 2773 3010 2779
rect 1987 2739 1999 2773
rect 2033 2740 2191 2773
rect 2033 2739 2045 2740
rect 1987 2733 2045 2739
rect 2179 2739 2191 2740
rect 2225 2740 2383 2773
rect 2225 2739 2237 2740
rect 2179 2733 2237 2739
rect 2371 2739 2383 2740
rect 2417 2740 2575 2773
rect 2417 2739 2429 2740
rect 2371 2733 2429 2739
rect 2563 2739 2575 2740
rect 2609 2740 2767 2773
rect 2609 2739 2621 2740
rect 2563 2733 2621 2739
rect 2755 2739 2767 2740
rect 2801 2740 2959 2773
rect 2801 2739 2813 2740
rect 2755 2733 2813 2739
rect 2947 2739 2959 2740
rect 2993 2740 3010 2773
rect 2993 2739 3005 2740
rect 2947 2733 3005 2739
rect 1636 2696 1682 2708
rect 1040 2510 1060 2690
rect 1240 2680 1260 2690
rect 1436 2680 1570 2691
rect 1636 2680 1642 2696
rect 1240 2679 1642 2680
rect 1240 2670 1442 2679
rect 1240 2540 1300 2670
rect 1360 2540 1442 2670
rect 1240 2530 1442 2540
rect 1240 2510 1260 2530
rect 1420 2520 1442 2530
rect 1040 2500 1260 2510
rect 1436 2191 1442 2520
rect 1476 2520 1530 2679
rect 1476 2191 1482 2520
rect 1436 2179 1482 2191
rect 1524 2191 1530 2520
rect 1564 2530 1642 2679
rect 1564 2191 1570 2530
rect 1636 2520 1642 2530
rect 1676 2520 1682 2696
rect 1636 2508 1682 2520
rect 1724 2696 1790 2708
rect 1724 2520 1730 2696
rect 1764 2600 1790 2696
rect 3050 2690 3080 3000
rect 3150 2780 3220 2800
rect 3150 2746 3166 2780
rect 3200 2746 3220 2780
rect 3150 2730 3220 2746
rect 3010 2684 3080 2690
rect 1849 2680 1895 2684
rect 2041 2680 2087 2684
rect 2233 2680 2279 2684
rect 2425 2680 2471 2684
rect 2617 2680 2663 2684
rect 2809 2680 2855 2684
rect 3001 2680 3080 2684
rect 1849 2672 3080 2680
rect 1764 2520 1770 2600
rect 1724 2508 1770 2520
rect 1670 2476 1730 2480
rect 1670 2470 1732 2476
rect 1670 2436 1686 2470
rect 1720 2436 1732 2470
rect 1670 2430 1732 2436
rect 1670 2420 1730 2430
rect 1524 2179 1570 2191
rect 750 1975 1250 2060
rect 1680 1975 1730 2420
rect 1849 2184 1855 2672
rect 1889 2470 2047 2672
rect 1889 2184 1895 2470
rect 1849 2172 1895 2184
rect 1945 2218 1991 2230
rect 1945 2120 1951 2218
rect 750 1925 1730 1975
rect 1920 2100 1951 2120
rect 1985 2120 1991 2218
rect 2041 2184 2047 2470
rect 2081 2470 2239 2672
rect 2081 2184 2087 2470
rect 2041 2172 2087 2184
rect 2137 2218 2183 2230
rect 2137 2120 2143 2218
rect 1985 2100 2143 2120
rect 1920 2000 1930 2100
rect 2040 2000 2143 2100
rect 1920 1980 1951 2000
rect 1985 1980 2143 2000
rect 750 1860 1250 1925
rect 1470 1676 1530 1690
rect 1470 1670 1532 1676
rect 1470 1636 1486 1670
rect 1520 1636 1532 1670
rect 1470 1630 1532 1636
rect 1675 1675 1725 1925
rect 1920 1880 1930 1980
rect 2040 1880 2143 1980
rect 1920 1860 1951 1880
rect 1985 1860 2143 1880
rect 1920 1760 1930 1860
rect 2040 1760 2143 1860
rect 1920 1730 1951 1760
rect 1985 1730 2143 1760
rect 2177 2120 2183 2218
rect 2233 2184 2239 2470
rect 2273 2470 2431 2672
rect 2273 2184 2279 2470
rect 2233 2172 2279 2184
rect 2329 2218 2375 2230
rect 2329 2120 2335 2218
rect 2177 1730 2335 2120
rect 2369 2120 2375 2218
rect 2425 2184 2431 2470
rect 2465 2470 2623 2672
rect 2465 2184 2471 2470
rect 2425 2172 2471 2184
rect 2521 2218 2567 2230
rect 2521 2120 2527 2218
rect 2369 1730 2527 2120
rect 2561 2120 2567 2218
rect 2617 2184 2623 2470
rect 2657 2470 2815 2672
rect 2657 2184 2663 2470
rect 2617 2172 2663 2184
rect 2713 2218 2759 2230
rect 2713 2120 2719 2218
rect 2561 1730 2719 2120
rect 2753 2120 2759 2218
rect 2809 2184 2815 2470
rect 2849 2470 3007 2672
rect 2849 2184 2855 2470
rect 2809 2172 2855 2184
rect 2905 2218 2951 2230
rect 2905 2120 2911 2218
rect 2753 1730 2911 2120
rect 2945 1870 2951 2218
rect 3001 2184 3007 2470
rect 3041 2470 3080 2672
rect 3041 2184 3047 2470
rect 3001 2172 3047 2184
rect 3116 2225 3162 2237
rect 3116 1870 3122 2225
rect 2945 1790 3122 1870
rect 2945 1730 2951 1790
rect 1945 1718 1991 1730
rect 2137 1718 2183 1730
rect 2329 1718 2375 1730
rect 2521 1718 2567 1730
rect 2713 1718 2759 1730
rect 2905 1718 2951 1730
rect 3110 1737 3122 1790
rect 3156 1870 3162 2225
rect 3204 2225 3250 2237
rect 3204 1870 3210 2225
rect 3156 1737 3210 1870
rect 3244 1870 3250 2225
rect 4030 2060 4230 9500
rect 7260 9400 7460 9450
rect 9300 9400 9500 10020
rect 11400 10190 11600 10300
rect 11400 10020 11430 10190
rect 11560 10020 11600 10190
rect 11400 9450 11600 10020
rect 13500 10190 14210 10200
rect 13500 10020 13600 10190
rect 13730 10020 14210 10190
rect 13500 10000 14210 10020
rect 7260 9200 9500 9400
rect 10500 9250 11600 9450
rect 6700 6610 7000 6650
rect 6700 6490 6730 6610
rect 6940 6490 7000 6610
rect 6700 5756 7000 6490
rect 6700 5550 6832 5756
rect 6826 5359 6832 5550
rect 6870 5550 7000 5756
rect 6870 5359 6876 5550
rect 6826 5347 6876 5359
rect 6826 5221 6876 5233
rect 6826 4940 6832 5221
rect 6750 4824 6832 4940
rect 6870 4940 6876 5221
rect 6870 4824 6950 4940
rect 4770 4311 4830 4330
rect 4770 4310 4782 4311
rect 4750 4277 4782 4310
rect 4816 4310 4830 4311
rect 4816 4277 4870 4310
rect 4750 4213 4870 4277
rect 4732 4201 4870 4213
rect 4732 3713 4738 4201
rect 4772 4180 4826 4201
rect 4772 3713 4778 4180
rect 4732 3701 4778 3713
rect 4820 3713 4826 4180
rect 4860 4180 4870 4201
rect 5060 4304 6310 4330
rect 5060 4270 5295 4304
rect 5329 4270 5487 4304
rect 5521 4270 5679 4304
rect 5713 4270 5871 4304
rect 5905 4270 6063 4304
rect 6097 4270 6255 4304
rect 6289 4270 6310 4304
rect 6470 4311 6530 4330
rect 6470 4277 6482 4311
rect 6516 4277 6530 4311
rect 6470 4270 6530 4277
rect 4860 3820 4866 4180
rect 4970 3911 5030 3930
rect 4970 3877 4982 3911
rect 5016 3877 5030 3911
rect 4970 3870 5030 3877
rect 5060 3830 5100 4270
rect 5283 4264 5341 4270
rect 5475 4264 5533 4270
rect 5667 4264 5725 4270
rect 5859 4264 5917 4270
rect 6051 4264 6109 4270
rect 6243 4264 6301 4270
rect 6432 4218 6478 4230
rect 4932 3820 4978 3830
rect 4860 3818 4978 3820
rect 4860 3713 4938 3818
rect 4340 3630 4560 3640
rect 4340 3450 4360 3630
rect 4540 3590 4560 3630
rect 4820 3590 4938 3713
rect 4540 3580 4938 3590
rect 4540 3490 4610 3580
rect 4660 3490 4938 3580
rect 4540 3480 4938 3490
rect 4540 3450 4560 3480
rect 4340 3440 4560 3450
rect 4820 3250 4938 3480
rect 4932 3242 4938 3250
rect 4972 3242 4978 3818
rect 4932 3230 4978 3242
rect 5020 3818 5100 3830
rect 5020 3242 5026 3818
rect 5060 3720 5100 3818
rect 5145 4200 5191 4206
rect 5337 4200 5383 4206
rect 5529 4200 5575 4206
rect 5721 4200 5767 4206
rect 5913 4200 5959 4206
rect 6105 4200 6151 4206
rect 6297 4200 6343 4206
rect 5145 4194 6343 4200
rect 5060 3380 5066 3720
rect 5145 3706 5151 4194
rect 5185 4050 5343 4194
rect 5185 3950 5190 4050
rect 5330 3950 5343 4050
rect 5185 3820 5343 3950
rect 5185 3706 5191 3820
rect 5145 3694 5191 3706
rect 5241 3740 5287 3752
rect 5241 3550 5247 3740
rect 5060 3242 5090 3380
rect 5230 3270 5247 3550
rect 5020 3230 5090 3242
rect 5241 3252 5247 3270
rect 5281 3550 5287 3740
rect 5337 3706 5343 3820
rect 5377 3820 5535 4194
rect 5377 3706 5383 3820
rect 5337 3694 5383 3706
rect 5433 3740 5479 3752
rect 5433 3550 5439 3740
rect 5281 3270 5439 3550
rect 5281 3252 5287 3270
rect 5241 3240 5287 3252
rect 5433 3252 5439 3270
rect 5473 3550 5479 3740
rect 5529 3706 5535 3820
rect 5569 3820 5727 4194
rect 5569 3706 5575 3820
rect 5529 3694 5575 3706
rect 5625 3740 5671 3752
rect 5625 3550 5631 3740
rect 5473 3270 5631 3550
rect 5473 3252 5479 3270
rect 5433 3240 5479 3252
rect 5625 3252 5631 3270
rect 5665 3550 5671 3740
rect 5721 3706 5727 3820
rect 5761 3820 5919 4194
rect 5761 3706 5767 3820
rect 5721 3694 5767 3706
rect 5817 3740 5863 3752
rect 5817 3550 5823 3740
rect 5665 3270 5823 3550
rect 5665 3252 5671 3270
rect 5625 3240 5671 3252
rect 5817 3252 5823 3270
rect 5857 3550 5863 3740
rect 5913 3706 5919 3820
rect 5953 3820 6111 4194
rect 5953 3706 5959 3820
rect 5913 3694 5959 3706
rect 6009 3740 6055 3752
rect 6009 3550 6015 3740
rect 5857 3270 6015 3550
rect 5857 3252 5863 3270
rect 5817 3240 5863 3252
rect 6009 3252 6015 3270
rect 6049 3550 6055 3740
rect 6105 3706 6111 3820
rect 6145 3820 6303 4194
rect 6145 3706 6151 3820
rect 6105 3694 6151 3706
rect 6201 3740 6247 3752
rect 6201 3550 6207 3740
rect 6049 3270 6207 3550
rect 6049 3252 6055 3270
rect 6009 3240 6055 3252
rect 6201 3252 6207 3270
rect 6241 3550 6247 3740
rect 6297 3706 6303 3820
rect 6337 3706 6343 4194
rect 6297 3694 6343 3706
rect 6241 3340 6380 3550
rect 6432 3340 6438 4218
rect 6241 3270 6438 3340
rect 6241 3252 6247 3270
rect 6280 3260 6438 3270
rect 6201 3240 6247 3252
rect 6350 3242 6438 3260
rect 6472 3340 6478 4218
rect 6520 4218 6566 4230
rect 6520 3340 6526 4218
rect 6472 3242 6526 3340
rect 6560 3340 6566 4218
rect 6560 3242 6590 3340
rect 4750 3183 4830 3190
rect 4750 3149 4782 3183
rect 4816 3149 4830 3183
rect 4750 3130 4830 3149
rect 4970 3183 5030 3190
rect 4970 3149 4982 3183
rect 5016 3149 5030 3183
rect 4740 2780 4860 2800
rect 4740 2746 4786 2780
rect 4820 2746 4860 2780
rect 4340 2690 4560 2700
rect 4740 2691 4860 2746
rect 4970 2786 5030 3149
rect 4970 2780 5032 2786
rect 4970 2746 4986 2780
rect 5020 2746 5032 2780
rect 4970 2740 5032 2746
rect 5060 2708 5090 3230
rect 5200 3182 6210 3190
rect 5187 3176 6210 3182
rect 5187 3142 5199 3176
rect 5233 3142 5391 3176
rect 5425 3142 5583 3176
rect 5617 3142 5775 3176
rect 5809 3142 5967 3176
rect 6001 3142 6159 3176
rect 6193 3142 6210 3176
rect 5187 3136 6210 3142
rect 5200 3130 6210 3136
rect 6350 3183 6590 3242
rect 6350 3149 6482 3183
rect 6516 3149 6590 3183
rect 6350 3100 6590 3149
rect 6750 3100 6950 4824
rect 6350 3000 6950 3100
rect 5290 2779 6310 2800
rect 5287 2773 6310 2779
rect 5287 2739 5299 2773
rect 5333 2740 5491 2773
rect 5333 2739 5345 2740
rect 5287 2733 5345 2739
rect 5479 2739 5491 2740
rect 5525 2740 5683 2773
rect 5525 2739 5537 2740
rect 5479 2733 5537 2739
rect 5671 2739 5683 2740
rect 5717 2740 5875 2773
rect 5717 2739 5729 2740
rect 5671 2733 5729 2739
rect 5863 2739 5875 2740
rect 5909 2740 6067 2773
rect 5909 2739 5921 2740
rect 5863 2733 5921 2739
rect 6055 2739 6067 2740
rect 6101 2740 6259 2773
rect 6101 2739 6113 2740
rect 6055 2733 6113 2739
rect 6247 2739 6259 2740
rect 6293 2740 6310 2773
rect 6293 2739 6305 2740
rect 6247 2733 6305 2739
rect 4936 2696 4982 2708
rect 4340 2510 4350 2690
rect 4530 2680 4560 2690
rect 4736 2680 4870 2691
rect 4936 2680 4942 2696
rect 4530 2679 4942 2680
rect 4530 2670 4742 2679
rect 4530 2540 4600 2670
rect 4660 2540 4742 2670
rect 4530 2530 4742 2540
rect 4530 2510 4560 2530
rect 4720 2520 4742 2530
rect 4340 2500 4560 2510
rect 4736 2191 4742 2520
rect 4776 2520 4830 2679
rect 4776 2191 4782 2520
rect 4736 2179 4782 2191
rect 4824 2191 4830 2520
rect 4864 2530 4942 2679
rect 4864 2191 4870 2530
rect 4936 2520 4942 2530
rect 4976 2520 4982 2696
rect 4936 2508 4982 2520
rect 5024 2696 5090 2708
rect 5024 2520 5030 2696
rect 5064 2600 5090 2696
rect 6350 2690 6380 3000
rect 6450 2780 6520 2800
rect 6450 2746 6466 2780
rect 6500 2746 6520 2780
rect 6450 2730 6520 2746
rect 6310 2684 6380 2690
rect 5149 2680 5195 2684
rect 5341 2680 5387 2684
rect 5533 2680 5579 2684
rect 5725 2680 5771 2684
rect 5917 2680 5963 2684
rect 6109 2680 6155 2684
rect 6301 2680 6380 2684
rect 5149 2672 6380 2680
rect 5064 2520 5070 2600
rect 5024 2508 5070 2520
rect 4970 2476 5030 2480
rect 4970 2470 5032 2476
rect 4970 2436 4986 2470
rect 5020 2436 5032 2470
rect 4970 2430 5032 2436
rect 4970 2420 5030 2430
rect 4824 2179 4870 2191
rect 4030 1975 4550 2060
rect 4980 1975 5030 2420
rect 5149 2184 5155 2672
rect 5189 2470 5347 2672
rect 5189 2184 5195 2470
rect 5149 2172 5195 2184
rect 5245 2218 5291 2230
rect 5245 2120 5251 2218
rect 4030 1925 5030 1975
rect 5220 2100 5251 2120
rect 5285 2120 5291 2218
rect 5341 2184 5347 2470
rect 5381 2470 5539 2672
rect 5381 2184 5387 2470
rect 5341 2172 5387 2184
rect 5437 2218 5483 2230
rect 5437 2120 5443 2218
rect 5285 2100 5443 2120
rect 5220 2000 5230 2100
rect 5340 2000 5443 2100
rect 5220 1980 5251 2000
rect 5285 1980 5443 2000
rect 3450 1870 3650 1920
rect 3244 1790 3650 1870
rect 4030 1860 4550 1925
rect 3244 1737 3250 1790
rect 1675 1669 1905 1675
rect 3110 1670 3250 1737
rect 1675 1663 1949 1669
rect 1675 1629 1903 1663
rect 1937 1660 1949 1663
rect 2083 1663 2141 1669
rect 2083 1660 2095 1663
rect 1937 1629 2095 1660
rect 2129 1660 2141 1663
rect 2275 1663 2333 1669
rect 2275 1660 2287 1663
rect 2129 1629 2287 1660
rect 2321 1660 2333 1663
rect 2467 1663 2525 1669
rect 2467 1660 2479 1663
rect 2321 1629 2479 1660
rect 2513 1660 2525 1663
rect 2659 1663 2717 1669
rect 2659 1660 2671 1663
rect 2513 1629 2671 1660
rect 2705 1660 2717 1663
rect 2851 1663 2909 1669
rect 2851 1660 2863 1663
rect 2705 1629 2863 1660
rect 2897 1660 2909 1663
rect 2897 1629 2910 1660
rect 3110 1636 3166 1670
rect 3200 1636 3250 1670
rect 3110 1630 3250 1636
rect 1675 1625 2910 1629
rect 1890 1600 2910 1625
rect 3150 1620 3210 1630
rect 3450 1250 3650 1790
rect 4770 1676 4830 1690
rect 4770 1670 4832 1676
rect 4770 1636 4786 1670
rect 4820 1636 4832 1670
rect 4770 1630 4832 1636
rect 4975 1675 5025 1925
rect 5220 1880 5230 1980
rect 5340 1880 5443 1980
rect 5220 1860 5251 1880
rect 5285 1860 5443 1880
rect 5220 1760 5230 1860
rect 5340 1760 5443 1860
rect 5220 1730 5251 1760
rect 5285 1730 5443 1760
rect 5477 2120 5483 2218
rect 5533 2184 5539 2470
rect 5573 2470 5731 2672
rect 5573 2184 5579 2470
rect 5533 2172 5579 2184
rect 5629 2218 5675 2230
rect 5629 2120 5635 2218
rect 5477 1730 5635 2120
rect 5669 2120 5675 2218
rect 5725 2184 5731 2470
rect 5765 2470 5923 2672
rect 5765 2184 5771 2470
rect 5725 2172 5771 2184
rect 5821 2218 5867 2230
rect 5821 2120 5827 2218
rect 5669 1730 5827 2120
rect 5861 2120 5867 2218
rect 5917 2184 5923 2470
rect 5957 2470 6115 2672
rect 5957 2184 5963 2470
rect 5917 2172 5963 2184
rect 6013 2218 6059 2230
rect 6013 2120 6019 2218
rect 5861 1730 6019 2120
rect 6053 2120 6059 2218
rect 6109 2184 6115 2470
rect 6149 2470 6307 2672
rect 6149 2184 6155 2470
rect 6109 2172 6155 2184
rect 6205 2218 6251 2230
rect 6205 2120 6211 2218
rect 6053 1730 6211 2120
rect 6245 1870 6251 2218
rect 6301 2184 6307 2470
rect 6341 2470 6380 2672
rect 6341 2184 6347 2470
rect 6301 2172 6347 2184
rect 6416 2225 6462 2237
rect 6416 1870 6422 2225
rect 6245 1790 6422 1870
rect 6245 1730 6251 1790
rect 5245 1718 5291 1730
rect 5437 1718 5483 1730
rect 5629 1718 5675 1730
rect 5821 1718 5867 1730
rect 6013 1718 6059 1730
rect 6205 1718 6251 1730
rect 6410 1737 6422 1790
rect 6456 1870 6462 2225
rect 6504 2225 6550 2237
rect 6504 1870 6510 2225
rect 6456 1737 6510 1870
rect 6544 1870 6550 2225
rect 7260 2060 7460 9200
rect 10000 6730 10300 6770
rect 10000 6470 10040 6730
rect 10240 6470 10300 6730
rect 10000 5896 10300 6470
rect 10000 5670 10132 5896
rect 10126 5499 10132 5670
rect 10170 5670 10300 5896
rect 10170 5499 10176 5670
rect 10126 5487 10176 5499
rect 10126 5221 10176 5233
rect 10126 4940 10132 5221
rect 10050 4824 10132 4940
rect 10170 4940 10176 5221
rect 10170 4824 10250 4940
rect 8070 4311 8130 4330
rect 8070 4310 8082 4311
rect 8050 4277 8082 4310
rect 8116 4310 8130 4311
rect 8116 4277 8170 4310
rect 8050 4213 8170 4277
rect 8032 4201 8170 4213
rect 8032 3713 8038 4201
rect 8072 4180 8126 4201
rect 8072 3713 8078 4180
rect 8032 3701 8078 3713
rect 8120 3713 8126 4180
rect 8160 4180 8170 4201
rect 8360 4304 9610 4330
rect 8360 4270 8595 4304
rect 8629 4270 8787 4304
rect 8821 4270 8979 4304
rect 9013 4270 9171 4304
rect 9205 4270 9363 4304
rect 9397 4270 9555 4304
rect 9589 4270 9610 4304
rect 9770 4311 9830 4330
rect 9770 4277 9782 4311
rect 9816 4277 9830 4311
rect 9770 4270 9830 4277
rect 8160 3820 8166 4180
rect 8270 3911 8330 3930
rect 8270 3877 8282 3911
rect 8316 3877 8330 3911
rect 8270 3870 8330 3877
rect 8360 3830 8400 4270
rect 8583 4264 8641 4270
rect 8775 4264 8833 4270
rect 8967 4264 9025 4270
rect 9159 4264 9217 4270
rect 9351 4264 9409 4270
rect 9543 4264 9601 4270
rect 9732 4218 9778 4230
rect 8232 3820 8278 3830
rect 8160 3818 8278 3820
rect 8160 3713 8238 3818
rect 7640 3630 7860 3640
rect 7640 3450 7660 3630
rect 7840 3590 7860 3630
rect 8120 3590 8238 3713
rect 7840 3580 8238 3590
rect 7840 3490 7910 3580
rect 7960 3490 8238 3580
rect 7840 3480 8238 3490
rect 7840 3450 7860 3480
rect 7640 3440 7860 3450
rect 8120 3250 8238 3480
rect 8232 3242 8238 3250
rect 8272 3242 8278 3818
rect 8232 3230 8278 3242
rect 8320 3818 8400 3830
rect 8320 3242 8326 3818
rect 8360 3720 8400 3818
rect 8445 4200 8491 4206
rect 8637 4200 8683 4206
rect 8829 4200 8875 4206
rect 9021 4200 9067 4206
rect 9213 4200 9259 4206
rect 9405 4200 9451 4206
rect 9597 4200 9643 4206
rect 8445 4194 9643 4200
rect 8360 3380 8366 3720
rect 8445 3706 8451 4194
rect 8485 4050 8643 4194
rect 8485 3950 8490 4050
rect 8630 3950 8643 4050
rect 8485 3820 8643 3950
rect 8485 3706 8491 3820
rect 8445 3694 8491 3706
rect 8541 3740 8587 3752
rect 8541 3550 8547 3740
rect 8360 3242 8390 3380
rect 8530 3270 8547 3550
rect 8320 3230 8390 3242
rect 8541 3252 8547 3270
rect 8581 3550 8587 3740
rect 8637 3706 8643 3820
rect 8677 3820 8835 4194
rect 8677 3706 8683 3820
rect 8637 3694 8683 3706
rect 8733 3740 8779 3752
rect 8733 3550 8739 3740
rect 8581 3270 8739 3550
rect 8581 3252 8587 3270
rect 8541 3240 8587 3252
rect 8733 3252 8739 3270
rect 8773 3550 8779 3740
rect 8829 3706 8835 3820
rect 8869 3820 9027 4194
rect 8869 3706 8875 3820
rect 8829 3694 8875 3706
rect 8925 3740 8971 3752
rect 8925 3550 8931 3740
rect 8773 3270 8931 3550
rect 8773 3252 8779 3270
rect 8733 3240 8779 3252
rect 8925 3252 8931 3270
rect 8965 3550 8971 3740
rect 9021 3706 9027 3820
rect 9061 3820 9219 4194
rect 9061 3706 9067 3820
rect 9021 3694 9067 3706
rect 9117 3740 9163 3752
rect 9117 3550 9123 3740
rect 8965 3270 9123 3550
rect 8965 3252 8971 3270
rect 8925 3240 8971 3252
rect 9117 3252 9123 3270
rect 9157 3550 9163 3740
rect 9213 3706 9219 3820
rect 9253 3820 9411 4194
rect 9253 3706 9259 3820
rect 9213 3694 9259 3706
rect 9309 3740 9355 3752
rect 9309 3550 9315 3740
rect 9157 3270 9315 3550
rect 9157 3252 9163 3270
rect 9117 3240 9163 3252
rect 9309 3252 9315 3270
rect 9349 3550 9355 3740
rect 9405 3706 9411 3820
rect 9445 3820 9603 4194
rect 9445 3706 9451 3820
rect 9405 3694 9451 3706
rect 9501 3740 9547 3752
rect 9501 3550 9507 3740
rect 9349 3270 9507 3550
rect 9349 3252 9355 3270
rect 9309 3240 9355 3252
rect 9501 3252 9507 3270
rect 9541 3550 9547 3740
rect 9597 3706 9603 3820
rect 9637 3706 9643 4194
rect 9597 3694 9643 3706
rect 9541 3340 9680 3550
rect 9732 3340 9738 4218
rect 9541 3270 9738 3340
rect 9541 3252 9547 3270
rect 9580 3260 9738 3270
rect 9501 3240 9547 3252
rect 9650 3242 9738 3260
rect 9772 3340 9778 4218
rect 9820 4218 9866 4230
rect 9820 3340 9826 4218
rect 9772 3242 9826 3340
rect 9860 3340 9866 4218
rect 9860 3242 9890 3340
rect 8050 3183 8130 3190
rect 8050 3149 8082 3183
rect 8116 3149 8130 3183
rect 8050 3130 8130 3149
rect 8270 3183 8330 3190
rect 8270 3149 8282 3183
rect 8316 3149 8330 3183
rect 8040 2780 8160 2800
rect 8040 2746 8086 2780
rect 8120 2746 8160 2780
rect 7640 2690 7860 2700
rect 8040 2691 8160 2746
rect 8270 2786 8330 3149
rect 8270 2780 8332 2786
rect 8270 2746 8286 2780
rect 8320 2746 8332 2780
rect 8270 2740 8332 2746
rect 8360 2708 8390 3230
rect 8500 3182 9510 3190
rect 8487 3176 9510 3182
rect 8487 3142 8499 3176
rect 8533 3142 8691 3176
rect 8725 3142 8883 3176
rect 8917 3142 9075 3176
rect 9109 3142 9267 3176
rect 9301 3142 9459 3176
rect 9493 3142 9510 3176
rect 8487 3136 9510 3142
rect 8500 3130 9510 3136
rect 9650 3183 9890 3242
rect 9650 3149 9782 3183
rect 9816 3149 9890 3183
rect 9650 3100 9890 3149
rect 10050 3100 10250 4824
rect 9650 3000 10250 3100
rect 8590 2779 9610 2800
rect 8587 2773 9610 2779
rect 8587 2739 8599 2773
rect 8633 2740 8791 2773
rect 8633 2739 8645 2740
rect 8587 2733 8645 2739
rect 8779 2739 8791 2740
rect 8825 2740 8983 2773
rect 8825 2739 8837 2740
rect 8779 2733 8837 2739
rect 8971 2739 8983 2740
rect 9017 2740 9175 2773
rect 9017 2739 9029 2740
rect 8971 2733 9029 2739
rect 9163 2739 9175 2740
rect 9209 2740 9367 2773
rect 9209 2739 9221 2740
rect 9163 2733 9221 2739
rect 9355 2739 9367 2740
rect 9401 2740 9559 2773
rect 9401 2739 9413 2740
rect 9355 2733 9413 2739
rect 9547 2739 9559 2740
rect 9593 2740 9610 2773
rect 9593 2739 9605 2740
rect 9547 2733 9605 2739
rect 8236 2696 8282 2708
rect 7640 2510 7660 2690
rect 7840 2680 7860 2690
rect 8036 2680 8170 2691
rect 8236 2680 8242 2696
rect 7840 2679 8242 2680
rect 7840 2670 8042 2679
rect 7840 2540 7900 2670
rect 7960 2540 8042 2670
rect 7840 2530 8042 2540
rect 7840 2510 7860 2530
rect 8020 2520 8042 2530
rect 7640 2500 7860 2510
rect 8036 2191 8042 2520
rect 8076 2520 8130 2679
rect 8076 2191 8082 2520
rect 8036 2179 8082 2191
rect 8124 2191 8130 2520
rect 8164 2530 8242 2679
rect 8164 2191 8170 2530
rect 8236 2520 8242 2530
rect 8276 2520 8282 2696
rect 8236 2508 8282 2520
rect 8324 2696 8390 2708
rect 8324 2520 8330 2696
rect 8364 2600 8390 2696
rect 9650 2690 9680 3000
rect 9750 2780 9820 2800
rect 9750 2746 9766 2780
rect 9800 2746 9820 2780
rect 9750 2730 9820 2746
rect 9610 2684 9680 2690
rect 8449 2680 8495 2684
rect 8641 2680 8687 2684
rect 8833 2680 8879 2684
rect 9025 2680 9071 2684
rect 9217 2680 9263 2684
rect 9409 2680 9455 2684
rect 9601 2680 9680 2684
rect 8449 2672 9680 2680
rect 8364 2520 8370 2600
rect 8324 2508 8370 2520
rect 8270 2476 8330 2480
rect 8270 2470 8332 2476
rect 8270 2436 8286 2470
rect 8320 2436 8332 2470
rect 8270 2430 8332 2436
rect 8270 2420 8330 2430
rect 8124 2179 8170 2191
rect 7260 1975 7850 2060
rect 8280 1975 8330 2420
rect 8449 2184 8455 2672
rect 8489 2470 8647 2672
rect 8489 2184 8495 2470
rect 8449 2172 8495 2184
rect 8545 2218 8591 2230
rect 8545 2120 8551 2218
rect 7260 1925 8330 1975
rect 8520 2100 8551 2120
rect 8585 2120 8591 2218
rect 8641 2184 8647 2470
rect 8681 2470 8839 2672
rect 8681 2184 8687 2470
rect 8641 2172 8687 2184
rect 8737 2218 8783 2230
rect 8737 2120 8743 2218
rect 8585 2100 8743 2120
rect 8520 2000 8530 2100
rect 8640 2000 8743 2100
rect 8520 1980 8551 2000
rect 8585 1980 8743 2000
rect 6750 1870 6950 1920
rect 6544 1790 6950 1870
rect 7260 1860 7850 1925
rect 6544 1737 6550 1790
rect 4975 1669 5205 1675
rect 6410 1670 6550 1737
rect 4975 1663 5249 1669
rect 4975 1629 5203 1663
rect 5237 1660 5249 1663
rect 5383 1663 5441 1669
rect 5383 1660 5395 1663
rect 5237 1629 5395 1660
rect 5429 1660 5441 1663
rect 5575 1663 5633 1669
rect 5575 1660 5587 1663
rect 5429 1629 5587 1660
rect 5621 1660 5633 1663
rect 5767 1663 5825 1669
rect 5767 1660 5779 1663
rect 5621 1629 5779 1660
rect 5813 1660 5825 1663
rect 5959 1663 6017 1669
rect 5959 1660 5971 1663
rect 5813 1629 5971 1660
rect 6005 1660 6017 1663
rect 6151 1663 6209 1669
rect 6151 1660 6163 1663
rect 6005 1629 6163 1660
rect 6197 1660 6209 1663
rect 6197 1629 6210 1660
rect 6410 1636 6466 1670
rect 6500 1636 6550 1670
rect 6410 1630 6550 1636
rect 4975 1625 6210 1629
rect 5190 1600 6210 1625
rect 6450 1620 6510 1630
rect 6750 1250 6950 1790
rect 8070 1676 8130 1690
rect 8070 1670 8132 1676
rect 8070 1636 8086 1670
rect 8120 1636 8132 1670
rect 8070 1630 8132 1636
rect 8275 1675 8325 1925
rect 8520 1880 8530 1980
rect 8640 1880 8743 1980
rect 8520 1860 8551 1880
rect 8585 1860 8743 1880
rect 8520 1760 8530 1860
rect 8640 1760 8743 1860
rect 8520 1730 8551 1760
rect 8585 1730 8743 1760
rect 8777 2120 8783 2218
rect 8833 2184 8839 2470
rect 8873 2470 9031 2672
rect 8873 2184 8879 2470
rect 8833 2172 8879 2184
rect 8929 2218 8975 2230
rect 8929 2120 8935 2218
rect 8777 1730 8935 2120
rect 8969 2120 8975 2218
rect 9025 2184 9031 2470
rect 9065 2470 9223 2672
rect 9065 2184 9071 2470
rect 9025 2172 9071 2184
rect 9121 2218 9167 2230
rect 9121 2120 9127 2218
rect 8969 1730 9127 2120
rect 9161 2120 9167 2218
rect 9217 2184 9223 2470
rect 9257 2470 9415 2672
rect 9257 2184 9263 2470
rect 9217 2172 9263 2184
rect 9313 2218 9359 2230
rect 9313 2120 9319 2218
rect 9161 1730 9319 2120
rect 9353 2120 9359 2218
rect 9409 2184 9415 2470
rect 9449 2470 9607 2672
rect 9449 2184 9455 2470
rect 9409 2172 9455 2184
rect 9505 2218 9551 2230
rect 9505 2120 9511 2218
rect 9353 1730 9511 2120
rect 9545 1870 9551 2218
rect 9601 2184 9607 2470
rect 9641 2470 9680 2672
rect 9641 2184 9647 2470
rect 9601 2172 9647 2184
rect 9716 2225 9762 2237
rect 9716 1870 9722 2225
rect 9545 1790 9722 1870
rect 9545 1730 9551 1790
rect 8545 1718 8591 1730
rect 8737 1718 8783 1730
rect 8929 1718 8975 1730
rect 9121 1718 9167 1730
rect 9313 1718 9359 1730
rect 9505 1718 9551 1730
rect 9710 1737 9722 1790
rect 9756 1870 9762 2225
rect 9804 2225 9850 2237
rect 9804 1870 9810 2225
rect 9756 1737 9810 1870
rect 9844 1870 9850 2225
rect 10500 2060 10700 9250
rect 13310 6790 13610 6890
rect 13310 6480 13360 6790
rect 13560 6480 13610 6790
rect 13310 6176 13610 6480
rect 13310 5790 13432 6176
rect 13426 5779 13432 5790
rect 13470 5790 13610 6176
rect 13470 5779 13476 5790
rect 13426 5767 13476 5779
rect 13426 5221 13476 5233
rect 13426 4940 13432 5221
rect 13350 4824 13432 4940
rect 13470 4940 13476 5221
rect 13470 4824 13550 4940
rect 11370 4311 11430 4330
rect 11370 4310 11382 4311
rect 11350 4277 11382 4310
rect 11416 4310 11430 4311
rect 11416 4277 11470 4310
rect 11350 4213 11470 4277
rect 11332 4201 11470 4213
rect 11332 3713 11338 4201
rect 11372 4180 11426 4201
rect 11372 3713 11378 4180
rect 11332 3701 11378 3713
rect 11420 3713 11426 4180
rect 11460 4180 11470 4201
rect 11660 4304 12910 4330
rect 11660 4270 11895 4304
rect 11929 4270 12087 4304
rect 12121 4270 12279 4304
rect 12313 4270 12471 4304
rect 12505 4270 12663 4304
rect 12697 4270 12855 4304
rect 12889 4270 12910 4304
rect 13070 4311 13130 4330
rect 13070 4277 13082 4311
rect 13116 4277 13130 4311
rect 13070 4270 13130 4277
rect 11460 3820 11466 4180
rect 11570 3911 11630 3930
rect 11570 3877 11582 3911
rect 11616 3877 11630 3911
rect 11570 3870 11630 3877
rect 11660 3830 11700 4270
rect 11883 4264 11941 4270
rect 12075 4264 12133 4270
rect 12267 4264 12325 4270
rect 12459 4264 12517 4270
rect 12651 4264 12709 4270
rect 12843 4264 12901 4270
rect 13032 4218 13078 4230
rect 11532 3820 11578 3830
rect 11460 3818 11578 3820
rect 11460 3713 11538 3818
rect 10940 3630 11160 3640
rect 10940 3450 10960 3630
rect 11140 3590 11160 3630
rect 11420 3590 11538 3713
rect 11140 3580 11538 3590
rect 11140 3490 11210 3580
rect 11260 3490 11538 3580
rect 11140 3480 11538 3490
rect 11140 3450 11160 3480
rect 10940 3440 11160 3450
rect 11420 3250 11538 3480
rect 11532 3242 11538 3250
rect 11572 3242 11578 3818
rect 11532 3230 11578 3242
rect 11620 3818 11700 3830
rect 11620 3242 11626 3818
rect 11660 3720 11700 3818
rect 11745 4200 11791 4206
rect 11937 4200 11983 4206
rect 12129 4200 12175 4206
rect 12321 4200 12367 4206
rect 12513 4200 12559 4206
rect 12705 4200 12751 4206
rect 12897 4200 12943 4206
rect 11745 4194 12943 4200
rect 11660 3380 11666 3720
rect 11745 3706 11751 4194
rect 11785 4050 11943 4194
rect 11785 3950 11790 4050
rect 11930 3950 11943 4050
rect 11785 3820 11943 3950
rect 11785 3706 11791 3820
rect 11745 3694 11791 3706
rect 11841 3740 11887 3752
rect 11841 3550 11847 3740
rect 11660 3242 11690 3380
rect 11830 3270 11847 3550
rect 11620 3230 11690 3242
rect 11841 3252 11847 3270
rect 11881 3550 11887 3740
rect 11937 3706 11943 3820
rect 11977 3820 12135 4194
rect 11977 3706 11983 3820
rect 11937 3694 11983 3706
rect 12033 3740 12079 3752
rect 12033 3550 12039 3740
rect 11881 3270 12039 3550
rect 11881 3252 11887 3270
rect 11841 3240 11887 3252
rect 12033 3252 12039 3270
rect 12073 3550 12079 3740
rect 12129 3706 12135 3820
rect 12169 3820 12327 4194
rect 12169 3706 12175 3820
rect 12129 3694 12175 3706
rect 12225 3740 12271 3752
rect 12225 3550 12231 3740
rect 12073 3270 12231 3550
rect 12073 3252 12079 3270
rect 12033 3240 12079 3252
rect 12225 3252 12231 3270
rect 12265 3550 12271 3740
rect 12321 3706 12327 3820
rect 12361 3820 12519 4194
rect 12361 3706 12367 3820
rect 12321 3694 12367 3706
rect 12417 3740 12463 3752
rect 12417 3550 12423 3740
rect 12265 3270 12423 3550
rect 12265 3252 12271 3270
rect 12225 3240 12271 3252
rect 12417 3252 12423 3270
rect 12457 3550 12463 3740
rect 12513 3706 12519 3820
rect 12553 3820 12711 4194
rect 12553 3706 12559 3820
rect 12513 3694 12559 3706
rect 12609 3740 12655 3752
rect 12609 3550 12615 3740
rect 12457 3270 12615 3550
rect 12457 3252 12463 3270
rect 12417 3240 12463 3252
rect 12609 3252 12615 3270
rect 12649 3550 12655 3740
rect 12705 3706 12711 3820
rect 12745 3820 12903 4194
rect 12745 3706 12751 3820
rect 12705 3694 12751 3706
rect 12801 3740 12847 3752
rect 12801 3550 12807 3740
rect 12649 3270 12807 3550
rect 12649 3252 12655 3270
rect 12609 3240 12655 3252
rect 12801 3252 12807 3270
rect 12841 3550 12847 3740
rect 12897 3706 12903 3820
rect 12937 3706 12943 4194
rect 12897 3694 12943 3706
rect 12841 3340 12980 3550
rect 13032 3340 13038 4218
rect 12841 3270 13038 3340
rect 12841 3252 12847 3270
rect 12880 3260 13038 3270
rect 12801 3240 12847 3252
rect 12950 3242 13038 3260
rect 13072 3340 13078 4218
rect 13120 4218 13166 4230
rect 13120 3340 13126 4218
rect 13072 3242 13126 3340
rect 13160 3340 13166 4218
rect 13160 3242 13190 3340
rect 11350 3183 11430 3190
rect 11350 3149 11382 3183
rect 11416 3149 11430 3183
rect 11350 3130 11430 3149
rect 11570 3183 11630 3190
rect 11570 3149 11582 3183
rect 11616 3149 11630 3183
rect 11340 2780 11460 2800
rect 11340 2746 11386 2780
rect 11420 2746 11460 2780
rect 10940 2690 11160 2700
rect 11340 2691 11460 2746
rect 11570 2786 11630 3149
rect 11570 2780 11632 2786
rect 11570 2746 11586 2780
rect 11620 2746 11632 2780
rect 11570 2740 11632 2746
rect 11660 2708 11690 3230
rect 11800 3182 12810 3190
rect 11787 3176 12810 3182
rect 11787 3142 11799 3176
rect 11833 3142 11991 3176
rect 12025 3142 12183 3176
rect 12217 3142 12375 3176
rect 12409 3142 12567 3176
rect 12601 3142 12759 3176
rect 12793 3142 12810 3176
rect 11787 3136 12810 3142
rect 11800 3130 12810 3136
rect 12950 3183 13190 3242
rect 12950 3149 13082 3183
rect 13116 3149 13190 3183
rect 12950 3100 13190 3149
rect 13350 3100 13550 4824
rect 12950 3000 13550 3100
rect 11890 2779 12910 2800
rect 11887 2773 12910 2779
rect 11887 2739 11899 2773
rect 11933 2740 12091 2773
rect 11933 2739 11945 2740
rect 11887 2733 11945 2739
rect 12079 2739 12091 2740
rect 12125 2740 12283 2773
rect 12125 2739 12137 2740
rect 12079 2733 12137 2739
rect 12271 2739 12283 2740
rect 12317 2740 12475 2773
rect 12317 2739 12329 2740
rect 12271 2733 12329 2739
rect 12463 2739 12475 2740
rect 12509 2740 12667 2773
rect 12509 2739 12521 2740
rect 12463 2733 12521 2739
rect 12655 2739 12667 2740
rect 12701 2740 12859 2773
rect 12701 2739 12713 2740
rect 12655 2733 12713 2739
rect 12847 2739 12859 2740
rect 12893 2740 12910 2773
rect 12893 2739 12905 2740
rect 12847 2733 12905 2739
rect 11536 2696 11582 2708
rect 10940 2510 10960 2690
rect 11140 2680 11160 2690
rect 11336 2680 11470 2691
rect 11536 2680 11542 2696
rect 11140 2679 11542 2680
rect 11140 2670 11342 2679
rect 11140 2540 11200 2670
rect 11260 2540 11342 2670
rect 11140 2530 11342 2540
rect 11140 2510 11160 2530
rect 11320 2520 11342 2530
rect 10940 2500 11160 2510
rect 11336 2191 11342 2520
rect 11376 2520 11430 2679
rect 11376 2191 11382 2520
rect 11336 2179 11382 2191
rect 11424 2191 11430 2520
rect 11464 2530 11542 2679
rect 11464 2191 11470 2530
rect 11536 2520 11542 2530
rect 11576 2520 11582 2696
rect 11536 2508 11582 2520
rect 11624 2696 11690 2708
rect 11624 2520 11630 2696
rect 11664 2600 11690 2696
rect 12950 2690 12980 3000
rect 13050 2780 13120 2800
rect 13050 2746 13066 2780
rect 13100 2746 13120 2780
rect 13050 2730 13120 2746
rect 12910 2684 12980 2690
rect 11749 2680 11795 2684
rect 11941 2680 11987 2684
rect 12133 2680 12179 2684
rect 12325 2680 12371 2684
rect 12517 2680 12563 2684
rect 12709 2680 12755 2684
rect 12901 2680 12980 2684
rect 11749 2672 12980 2680
rect 11664 2520 11670 2600
rect 11624 2508 11670 2520
rect 11570 2476 11630 2480
rect 11570 2470 11632 2476
rect 11570 2436 11586 2470
rect 11620 2436 11632 2470
rect 11570 2430 11632 2436
rect 11570 2420 11630 2430
rect 11424 2179 11470 2191
rect 10500 1975 11150 2060
rect 11580 1975 11630 2420
rect 11749 2184 11755 2672
rect 11789 2470 11947 2672
rect 11789 2184 11795 2470
rect 11749 2172 11795 2184
rect 11845 2218 11891 2230
rect 11845 2120 11851 2218
rect 10500 1925 11630 1975
rect 11820 2100 11851 2120
rect 11885 2120 11891 2218
rect 11941 2184 11947 2470
rect 11981 2470 12139 2672
rect 11981 2184 11987 2470
rect 11941 2172 11987 2184
rect 12037 2218 12083 2230
rect 12037 2120 12043 2218
rect 11885 2100 12043 2120
rect 11820 2000 11830 2100
rect 11940 2000 12043 2100
rect 11820 1980 11851 2000
rect 11885 1980 12043 2000
rect 10050 1870 10250 1920
rect 9844 1790 10250 1870
rect 10500 1860 11150 1925
rect 9844 1737 9850 1790
rect 8275 1669 8505 1675
rect 9710 1670 9850 1737
rect 8275 1663 8549 1669
rect 8275 1629 8503 1663
rect 8537 1660 8549 1663
rect 8683 1663 8741 1669
rect 8683 1660 8695 1663
rect 8537 1629 8695 1660
rect 8729 1660 8741 1663
rect 8875 1663 8933 1669
rect 8875 1660 8887 1663
rect 8729 1629 8887 1660
rect 8921 1660 8933 1663
rect 9067 1663 9125 1669
rect 9067 1660 9079 1663
rect 8921 1629 9079 1660
rect 9113 1660 9125 1663
rect 9259 1663 9317 1669
rect 9259 1660 9271 1663
rect 9113 1629 9271 1660
rect 9305 1660 9317 1663
rect 9451 1663 9509 1669
rect 9451 1660 9463 1663
rect 9305 1629 9463 1660
rect 9497 1660 9509 1663
rect 9497 1629 9510 1660
rect 9710 1636 9766 1670
rect 9800 1636 9850 1670
rect 9710 1630 9850 1636
rect 8275 1625 9510 1629
rect 8490 1600 9510 1625
rect 9750 1620 9810 1630
rect 10050 1250 10250 1790
rect 11370 1676 11430 1690
rect 11370 1670 11432 1676
rect 11370 1636 11386 1670
rect 11420 1636 11432 1670
rect 11370 1630 11432 1636
rect 11575 1675 11625 1925
rect 11820 1880 11830 1980
rect 11940 1880 12043 1980
rect 11820 1860 11851 1880
rect 11885 1860 12043 1880
rect 11820 1760 11830 1860
rect 11940 1760 12043 1860
rect 11820 1730 11851 1760
rect 11885 1730 12043 1760
rect 12077 2120 12083 2218
rect 12133 2184 12139 2470
rect 12173 2470 12331 2672
rect 12173 2184 12179 2470
rect 12133 2172 12179 2184
rect 12229 2218 12275 2230
rect 12229 2120 12235 2218
rect 12077 1730 12235 2120
rect 12269 2120 12275 2218
rect 12325 2184 12331 2470
rect 12365 2470 12523 2672
rect 12365 2184 12371 2470
rect 12325 2172 12371 2184
rect 12421 2218 12467 2230
rect 12421 2120 12427 2218
rect 12269 1730 12427 2120
rect 12461 2120 12467 2218
rect 12517 2184 12523 2470
rect 12557 2470 12715 2672
rect 12557 2184 12563 2470
rect 12517 2172 12563 2184
rect 12613 2218 12659 2230
rect 12613 2120 12619 2218
rect 12461 1730 12619 2120
rect 12653 2120 12659 2218
rect 12709 2184 12715 2470
rect 12749 2470 12907 2672
rect 12749 2184 12755 2470
rect 12709 2172 12755 2184
rect 12805 2218 12851 2230
rect 12805 2120 12811 2218
rect 12653 1730 12811 2120
rect 12845 1870 12851 2218
rect 12901 2184 12907 2470
rect 12941 2470 12980 2672
rect 12941 2184 12947 2470
rect 12901 2172 12947 2184
rect 13016 2225 13062 2237
rect 13016 1870 13022 2225
rect 12845 1790 13022 1870
rect 12845 1730 12851 1790
rect 11845 1718 11891 1730
rect 12037 1718 12083 1730
rect 12229 1718 12275 1730
rect 12421 1718 12467 1730
rect 12613 1718 12659 1730
rect 12805 1718 12851 1730
rect 13010 1737 13022 1790
rect 13056 1870 13062 2225
rect 13104 2225 13150 2237
rect 13104 1870 13110 2225
rect 13056 1737 13110 1870
rect 13144 1870 13150 2225
rect 14010 2060 14210 10000
rect 15700 10190 15900 10300
rect 15700 10020 15720 10190
rect 15850 10020 15900 10190
rect 15700 9450 15900 10020
rect 17700 10180 18700 10200
rect 17700 10010 17810 10180
rect 17940 10010 18700 10180
rect 17700 10000 18700 10010
rect 19900 10190 24910 10200
rect 19900 10020 19940 10190
rect 20070 10020 24910 10190
rect 19900 10000 24910 10020
rect 18500 9450 18700 10000
rect 15700 9250 17750 9450
rect 18500 9250 21380 9450
rect 16850 6810 17200 6860
rect 16850 6500 16930 6810
rect 17150 6500 17200 6810
rect 16850 6460 17032 6500
rect 17026 6339 17032 6460
rect 17070 6460 17200 6500
rect 17070 6339 17076 6460
rect 17026 6327 17076 6339
rect 17026 5221 17076 5233
rect 17026 4940 17032 5221
rect 16950 4824 17032 4940
rect 17070 4940 17076 5221
rect 17070 4824 17150 4940
rect 14970 4311 15030 4330
rect 14970 4310 14982 4311
rect 14950 4277 14982 4310
rect 15016 4310 15030 4311
rect 15016 4277 15070 4310
rect 14950 4213 15070 4277
rect 14932 4201 15070 4213
rect 14932 3713 14938 4201
rect 14972 4180 15026 4201
rect 14972 3713 14978 4180
rect 14932 3701 14978 3713
rect 15020 3713 15026 4180
rect 15060 4180 15070 4201
rect 15260 4304 16510 4330
rect 15260 4270 15495 4304
rect 15529 4270 15687 4304
rect 15721 4270 15879 4304
rect 15913 4270 16071 4304
rect 16105 4270 16263 4304
rect 16297 4270 16455 4304
rect 16489 4270 16510 4304
rect 16670 4311 16730 4330
rect 16670 4277 16682 4311
rect 16716 4277 16730 4311
rect 16670 4270 16730 4277
rect 15060 3820 15066 4180
rect 15170 3911 15230 3930
rect 15170 3877 15182 3911
rect 15216 3877 15230 3911
rect 15170 3870 15230 3877
rect 15260 3830 15300 4270
rect 15483 4264 15541 4270
rect 15675 4264 15733 4270
rect 15867 4264 15925 4270
rect 16059 4264 16117 4270
rect 16251 4264 16309 4270
rect 16443 4264 16501 4270
rect 16632 4218 16678 4230
rect 15132 3820 15178 3830
rect 15060 3818 15178 3820
rect 15060 3713 15138 3818
rect 14540 3630 14760 3640
rect 14540 3450 14560 3630
rect 14740 3590 14760 3630
rect 15020 3590 15138 3713
rect 14740 3580 15138 3590
rect 14740 3490 14810 3580
rect 14860 3490 15138 3580
rect 14740 3480 15138 3490
rect 14740 3450 14760 3480
rect 14540 3440 14760 3450
rect 15020 3250 15138 3480
rect 15132 3242 15138 3250
rect 15172 3242 15178 3818
rect 15132 3230 15178 3242
rect 15220 3818 15300 3830
rect 15220 3242 15226 3818
rect 15260 3720 15300 3818
rect 15345 4200 15391 4206
rect 15537 4200 15583 4206
rect 15729 4200 15775 4206
rect 15921 4200 15967 4206
rect 16113 4200 16159 4206
rect 16305 4200 16351 4206
rect 16497 4200 16543 4206
rect 15345 4194 16543 4200
rect 15260 3380 15266 3720
rect 15345 3706 15351 4194
rect 15385 4050 15543 4194
rect 15385 3950 15390 4050
rect 15530 3950 15543 4050
rect 15385 3820 15543 3950
rect 15385 3706 15391 3820
rect 15345 3694 15391 3706
rect 15441 3740 15487 3752
rect 15441 3550 15447 3740
rect 15260 3242 15290 3380
rect 15430 3270 15447 3550
rect 15220 3230 15290 3242
rect 15441 3252 15447 3270
rect 15481 3550 15487 3740
rect 15537 3706 15543 3820
rect 15577 3820 15735 4194
rect 15577 3706 15583 3820
rect 15537 3694 15583 3706
rect 15633 3740 15679 3752
rect 15633 3550 15639 3740
rect 15481 3270 15639 3550
rect 15481 3252 15487 3270
rect 15441 3240 15487 3252
rect 15633 3252 15639 3270
rect 15673 3550 15679 3740
rect 15729 3706 15735 3820
rect 15769 3820 15927 4194
rect 15769 3706 15775 3820
rect 15729 3694 15775 3706
rect 15825 3740 15871 3752
rect 15825 3550 15831 3740
rect 15673 3270 15831 3550
rect 15673 3252 15679 3270
rect 15633 3240 15679 3252
rect 15825 3252 15831 3270
rect 15865 3550 15871 3740
rect 15921 3706 15927 3820
rect 15961 3820 16119 4194
rect 15961 3706 15967 3820
rect 15921 3694 15967 3706
rect 16017 3740 16063 3752
rect 16017 3550 16023 3740
rect 15865 3270 16023 3550
rect 15865 3252 15871 3270
rect 15825 3240 15871 3252
rect 16017 3252 16023 3270
rect 16057 3550 16063 3740
rect 16113 3706 16119 3820
rect 16153 3820 16311 4194
rect 16153 3706 16159 3820
rect 16113 3694 16159 3706
rect 16209 3740 16255 3752
rect 16209 3550 16215 3740
rect 16057 3270 16215 3550
rect 16057 3252 16063 3270
rect 16017 3240 16063 3252
rect 16209 3252 16215 3270
rect 16249 3550 16255 3740
rect 16305 3706 16311 3820
rect 16345 3820 16503 4194
rect 16345 3706 16351 3820
rect 16305 3694 16351 3706
rect 16401 3740 16447 3752
rect 16401 3550 16407 3740
rect 16249 3270 16407 3550
rect 16249 3252 16255 3270
rect 16209 3240 16255 3252
rect 16401 3252 16407 3270
rect 16441 3550 16447 3740
rect 16497 3706 16503 3820
rect 16537 3706 16543 4194
rect 16497 3694 16543 3706
rect 16441 3340 16580 3550
rect 16632 3340 16638 4218
rect 16441 3270 16638 3340
rect 16441 3252 16447 3270
rect 16480 3260 16638 3270
rect 16401 3240 16447 3252
rect 16550 3242 16638 3260
rect 16672 3340 16678 4218
rect 16720 4218 16766 4230
rect 16720 3340 16726 4218
rect 16672 3242 16726 3340
rect 16760 3340 16766 4218
rect 16760 3242 16790 3340
rect 14950 3183 15030 3190
rect 14950 3149 14982 3183
rect 15016 3149 15030 3183
rect 14950 3130 15030 3149
rect 15170 3183 15230 3190
rect 15170 3149 15182 3183
rect 15216 3149 15230 3183
rect 14940 2780 15060 2800
rect 14940 2746 14986 2780
rect 15020 2746 15060 2780
rect 14540 2690 14760 2700
rect 14940 2691 15060 2746
rect 15170 2786 15230 3149
rect 15170 2780 15232 2786
rect 15170 2746 15186 2780
rect 15220 2746 15232 2780
rect 15170 2740 15232 2746
rect 15260 2708 15290 3230
rect 15400 3182 16410 3190
rect 15387 3176 16410 3182
rect 15387 3142 15399 3176
rect 15433 3142 15591 3176
rect 15625 3142 15783 3176
rect 15817 3142 15975 3176
rect 16009 3142 16167 3176
rect 16201 3142 16359 3176
rect 16393 3142 16410 3176
rect 15387 3136 16410 3142
rect 15400 3130 16410 3136
rect 16550 3183 16790 3242
rect 16550 3149 16682 3183
rect 16716 3149 16790 3183
rect 16550 3100 16790 3149
rect 16950 3100 17150 4824
rect 16550 3000 17150 3100
rect 15490 2779 16510 2800
rect 15487 2773 16510 2779
rect 15487 2739 15499 2773
rect 15533 2740 15691 2773
rect 15533 2739 15545 2740
rect 15487 2733 15545 2739
rect 15679 2739 15691 2740
rect 15725 2740 15883 2773
rect 15725 2739 15737 2740
rect 15679 2733 15737 2739
rect 15871 2739 15883 2740
rect 15917 2740 16075 2773
rect 15917 2739 15929 2740
rect 15871 2733 15929 2739
rect 16063 2739 16075 2740
rect 16109 2740 16267 2773
rect 16109 2739 16121 2740
rect 16063 2733 16121 2739
rect 16255 2739 16267 2740
rect 16301 2740 16459 2773
rect 16301 2739 16313 2740
rect 16255 2733 16313 2739
rect 16447 2739 16459 2740
rect 16493 2740 16510 2773
rect 16493 2739 16505 2740
rect 16447 2733 16505 2739
rect 15136 2696 15182 2708
rect 14540 2510 14550 2690
rect 14730 2680 14760 2690
rect 14936 2680 15070 2691
rect 15136 2680 15142 2696
rect 14730 2679 15142 2680
rect 14730 2670 14942 2679
rect 14730 2540 14800 2670
rect 14860 2540 14942 2670
rect 14730 2530 14942 2540
rect 14730 2510 14760 2530
rect 14920 2520 14942 2530
rect 14540 2500 14760 2510
rect 14936 2191 14942 2520
rect 14976 2520 15030 2679
rect 14976 2191 14982 2520
rect 14936 2179 14982 2191
rect 15024 2191 15030 2520
rect 15064 2530 15142 2679
rect 15064 2191 15070 2530
rect 15136 2520 15142 2530
rect 15176 2520 15182 2696
rect 15136 2508 15182 2520
rect 15224 2696 15290 2708
rect 15224 2520 15230 2696
rect 15264 2600 15290 2696
rect 16550 2690 16580 3000
rect 16650 2780 16720 2800
rect 16650 2746 16666 2780
rect 16700 2746 16720 2780
rect 16650 2730 16720 2746
rect 16510 2684 16580 2690
rect 15349 2680 15395 2684
rect 15541 2680 15587 2684
rect 15733 2680 15779 2684
rect 15925 2680 15971 2684
rect 16117 2680 16163 2684
rect 16309 2680 16355 2684
rect 16501 2680 16580 2684
rect 15349 2672 16580 2680
rect 15264 2520 15270 2600
rect 15224 2508 15270 2520
rect 15170 2476 15230 2480
rect 15170 2470 15232 2476
rect 15170 2436 15186 2470
rect 15220 2436 15232 2470
rect 15170 2430 15232 2436
rect 15170 2420 15230 2430
rect 15024 2179 15070 2191
rect 14010 1975 14750 2060
rect 15180 1975 15230 2420
rect 15349 2184 15355 2672
rect 15389 2470 15547 2672
rect 15389 2184 15395 2470
rect 15349 2172 15395 2184
rect 15445 2218 15491 2230
rect 15445 2120 15451 2218
rect 14010 1925 15230 1975
rect 15420 2100 15451 2120
rect 15485 2120 15491 2218
rect 15541 2184 15547 2470
rect 15581 2470 15739 2672
rect 15581 2184 15587 2470
rect 15541 2172 15587 2184
rect 15637 2218 15683 2230
rect 15637 2120 15643 2218
rect 15485 2100 15643 2120
rect 15420 2000 15430 2100
rect 15540 2000 15643 2100
rect 15420 1980 15451 2000
rect 15485 1980 15643 2000
rect 13350 1870 13550 1920
rect 13144 1790 13550 1870
rect 14010 1860 14750 1925
rect 13144 1737 13150 1790
rect 11575 1669 11805 1675
rect 13010 1670 13150 1737
rect 11575 1663 11849 1669
rect 11575 1629 11803 1663
rect 11837 1660 11849 1663
rect 11983 1663 12041 1669
rect 11983 1660 11995 1663
rect 11837 1629 11995 1660
rect 12029 1660 12041 1663
rect 12175 1663 12233 1669
rect 12175 1660 12187 1663
rect 12029 1629 12187 1660
rect 12221 1660 12233 1663
rect 12367 1663 12425 1669
rect 12367 1660 12379 1663
rect 12221 1629 12379 1660
rect 12413 1660 12425 1663
rect 12559 1663 12617 1669
rect 12559 1660 12571 1663
rect 12413 1629 12571 1660
rect 12605 1660 12617 1663
rect 12751 1663 12809 1669
rect 12751 1660 12763 1663
rect 12605 1629 12763 1660
rect 12797 1660 12809 1663
rect 12797 1629 12810 1660
rect 13010 1636 13066 1670
rect 13100 1636 13150 1670
rect 13010 1630 13150 1636
rect 11575 1625 12810 1629
rect 11790 1600 12810 1625
rect 13050 1620 13110 1630
rect 13350 1250 13550 1790
rect 14970 1676 15030 1690
rect 14970 1670 15032 1676
rect 14970 1636 14986 1670
rect 15020 1636 15032 1670
rect 14970 1630 15032 1636
rect 15175 1675 15225 1925
rect 15420 1880 15430 1980
rect 15540 1880 15643 1980
rect 15420 1860 15451 1880
rect 15485 1860 15643 1880
rect 15420 1760 15430 1860
rect 15540 1760 15643 1860
rect 15420 1730 15451 1760
rect 15485 1730 15643 1760
rect 15677 2120 15683 2218
rect 15733 2184 15739 2470
rect 15773 2470 15931 2672
rect 15773 2184 15779 2470
rect 15733 2172 15779 2184
rect 15829 2218 15875 2230
rect 15829 2120 15835 2218
rect 15677 1730 15835 2120
rect 15869 2120 15875 2218
rect 15925 2184 15931 2470
rect 15965 2470 16123 2672
rect 15965 2184 15971 2470
rect 15925 2172 15971 2184
rect 16021 2218 16067 2230
rect 16021 2120 16027 2218
rect 15869 1730 16027 2120
rect 16061 2120 16067 2218
rect 16117 2184 16123 2470
rect 16157 2470 16315 2672
rect 16157 2184 16163 2470
rect 16117 2172 16163 2184
rect 16213 2218 16259 2230
rect 16213 2120 16219 2218
rect 16061 1730 16219 2120
rect 16253 2120 16259 2218
rect 16309 2184 16315 2470
rect 16349 2470 16507 2672
rect 16349 2184 16355 2470
rect 16309 2172 16355 2184
rect 16405 2218 16451 2230
rect 16405 2120 16411 2218
rect 16253 1730 16411 2120
rect 16445 1870 16451 2218
rect 16501 2184 16507 2470
rect 16541 2470 16580 2672
rect 16541 2184 16547 2470
rect 16501 2172 16547 2184
rect 16616 2225 16662 2237
rect 16616 1870 16622 2225
rect 16445 1790 16622 1870
rect 16445 1730 16451 1790
rect 15445 1718 15491 1730
rect 15637 1718 15683 1730
rect 15829 1718 15875 1730
rect 16021 1718 16067 1730
rect 16213 1718 16259 1730
rect 16405 1718 16451 1730
rect 16610 1737 16622 1790
rect 16656 1870 16662 2225
rect 16704 2225 16750 2237
rect 16704 1870 16710 2225
rect 16656 1737 16710 1870
rect 16744 1870 16750 2225
rect 17550 2060 17750 9250
rect 19450 6780 19870 6840
rect 19450 6490 19490 6780
rect 19820 6490 19870 6780
rect 19450 5240 19870 6490
rect 20226 6736 20276 6748
rect 20226 6339 20232 6736
rect 20270 6710 20276 6736
rect 20544 6736 20594 6748
rect 20544 6710 20550 6736
rect 20270 6350 20550 6710
rect 20270 6339 20276 6350
rect 20226 6327 20276 6339
rect 20544 6339 20550 6350
rect 20588 6339 20594 6736
rect 20544 6327 20594 6339
rect 19450 5233 20260 5240
rect 19450 5221 20276 5233
rect 19450 4824 20232 5221
rect 20270 4824 20276 5221
rect 20544 5221 20594 5233
rect 20544 4940 20550 5221
rect 19450 4820 20276 4824
rect 20226 4812 20276 4820
rect 20450 4824 20550 4940
rect 20588 4940 20594 5221
rect 20588 4824 20650 4940
rect 18470 4311 18530 4330
rect 18470 4310 18482 4311
rect 18450 4277 18482 4310
rect 18516 4310 18530 4311
rect 18516 4277 18570 4310
rect 18450 4213 18570 4277
rect 18432 4201 18570 4213
rect 18432 3713 18438 4201
rect 18472 4180 18526 4201
rect 18472 3713 18478 4180
rect 18432 3701 18478 3713
rect 18520 3713 18526 4180
rect 18560 4180 18570 4201
rect 18760 4304 20010 4330
rect 18760 4270 18995 4304
rect 19029 4270 19187 4304
rect 19221 4270 19379 4304
rect 19413 4270 19571 4304
rect 19605 4270 19763 4304
rect 19797 4270 19955 4304
rect 19989 4270 20010 4304
rect 20170 4311 20230 4330
rect 20170 4277 20182 4311
rect 20216 4277 20230 4311
rect 20170 4270 20230 4277
rect 18560 3820 18566 4180
rect 18670 3911 18730 3930
rect 18670 3877 18682 3911
rect 18716 3877 18730 3911
rect 18670 3870 18730 3877
rect 18760 3830 18800 4270
rect 18983 4264 19041 4270
rect 19175 4264 19233 4270
rect 19367 4264 19425 4270
rect 19559 4264 19617 4270
rect 19751 4264 19809 4270
rect 19943 4264 20001 4270
rect 20132 4218 20178 4230
rect 18632 3820 18678 3830
rect 18560 3818 18678 3820
rect 18560 3713 18638 3818
rect 18040 3630 18260 3640
rect 18040 3450 18060 3630
rect 18240 3590 18260 3630
rect 18520 3590 18638 3713
rect 18240 3580 18638 3590
rect 18240 3490 18310 3580
rect 18360 3490 18638 3580
rect 18240 3480 18638 3490
rect 18240 3450 18260 3480
rect 18040 3440 18260 3450
rect 18520 3250 18638 3480
rect 18632 3242 18638 3250
rect 18672 3242 18678 3818
rect 18632 3230 18678 3242
rect 18720 3818 18800 3830
rect 18720 3242 18726 3818
rect 18760 3720 18800 3818
rect 18845 4200 18891 4206
rect 19037 4200 19083 4206
rect 19229 4200 19275 4206
rect 19421 4200 19467 4206
rect 19613 4200 19659 4206
rect 19805 4200 19851 4206
rect 19997 4200 20043 4206
rect 18845 4194 20043 4200
rect 18760 3380 18766 3720
rect 18845 3706 18851 4194
rect 18885 4050 19043 4194
rect 18885 3950 18890 4050
rect 19030 3950 19043 4050
rect 18885 3820 19043 3950
rect 18885 3706 18891 3820
rect 18845 3694 18891 3706
rect 18941 3740 18987 3752
rect 18941 3550 18947 3740
rect 18760 3242 18790 3380
rect 18930 3270 18947 3550
rect 18720 3230 18790 3242
rect 18941 3252 18947 3270
rect 18981 3550 18987 3740
rect 19037 3706 19043 3820
rect 19077 3820 19235 4194
rect 19077 3706 19083 3820
rect 19037 3694 19083 3706
rect 19133 3740 19179 3752
rect 19133 3550 19139 3740
rect 18981 3270 19139 3550
rect 18981 3252 18987 3270
rect 18941 3240 18987 3252
rect 19133 3252 19139 3270
rect 19173 3550 19179 3740
rect 19229 3706 19235 3820
rect 19269 3820 19427 4194
rect 19269 3706 19275 3820
rect 19229 3694 19275 3706
rect 19325 3740 19371 3752
rect 19325 3550 19331 3740
rect 19173 3270 19331 3550
rect 19173 3252 19179 3270
rect 19133 3240 19179 3252
rect 19325 3252 19331 3270
rect 19365 3550 19371 3740
rect 19421 3706 19427 3820
rect 19461 3820 19619 4194
rect 19461 3706 19467 3820
rect 19421 3694 19467 3706
rect 19517 3740 19563 3752
rect 19517 3550 19523 3740
rect 19365 3270 19523 3550
rect 19365 3252 19371 3270
rect 19325 3240 19371 3252
rect 19517 3252 19523 3270
rect 19557 3550 19563 3740
rect 19613 3706 19619 3820
rect 19653 3820 19811 4194
rect 19653 3706 19659 3820
rect 19613 3694 19659 3706
rect 19709 3740 19755 3752
rect 19709 3550 19715 3740
rect 19557 3270 19715 3550
rect 19557 3252 19563 3270
rect 19517 3240 19563 3252
rect 19709 3252 19715 3270
rect 19749 3550 19755 3740
rect 19805 3706 19811 3820
rect 19845 3820 20003 4194
rect 19845 3706 19851 3820
rect 19805 3694 19851 3706
rect 19901 3740 19947 3752
rect 19901 3550 19907 3740
rect 19749 3270 19907 3550
rect 19749 3252 19755 3270
rect 19709 3240 19755 3252
rect 19901 3252 19907 3270
rect 19941 3550 19947 3740
rect 19997 3706 20003 3820
rect 20037 3706 20043 4194
rect 19997 3694 20043 3706
rect 19941 3340 20080 3550
rect 20132 3340 20138 4218
rect 19941 3270 20138 3340
rect 19941 3252 19947 3270
rect 19980 3260 20138 3270
rect 19901 3240 19947 3252
rect 20050 3242 20138 3260
rect 20172 3340 20178 4218
rect 20220 4218 20266 4230
rect 20220 3340 20226 4218
rect 20172 3242 20226 3340
rect 20260 3340 20266 4218
rect 20260 3242 20290 3340
rect 18450 3183 18530 3190
rect 18450 3149 18482 3183
rect 18516 3149 18530 3183
rect 18450 3130 18530 3149
rect 18670 3183 18730 3190
rect 18670 3149 18682 3183
rect 18716 3149 18730 3183
rect 18440 2780 18560 2800
rect 18440 2746 18486 2780
rect 18520 2746 18560 2780
rect 18040 2680 18260 2700
rect 18440 2691 18560 2746
rect 18670 2786 18730 3149
rect 18670 2780 18732 2786
rect 18670 2746 18686 2780
rect 18720 2746 18732 2780
rect 18670 2740 18732 2746
rect 18760 2708 18790 3230
rect 18900 3182 19910 3190
rect 18887 3176 19910 3182
rect 18887 3142 18899 3176
rect 18933 3142 19091 3176
rect 19125 3142 19283 3176
rect 19317 3142 19475 3176
rect 19509 3142 19667 3176
rect 19701 3142 19859 3176
rect 19893 3142 19910 3176
rect 18887 3136 19910 3142
rect 18900 3130 19910 3136
rect 20050 3183 20290 3242
rect 20050 3149 20182 3183
rect 20216 3149 20290 3183
rect 20050 3100 20290 3149
rect 20450 3100 20650 4824
rect 20050 3000 20650 3100
rect 18990 2779 20010 2800
rect 18987 2773 20010 2779
rect 18987 2739 18999 2773
rect 19033 2740 19191 2773
rect 19033 2739 19045 2740
rect 18987 2733 19045 2739
rect 19179 2739 19191 2740
rect 19225 2740 19383 2773
rect 19225 2739 19237 2740
rect 19179 2733 19237 2739
rect 19371 2739 19383 2740
rect 19417 2740 19575 2773
rect 19417 2739 19429 2740
rect 19371 2733 19429 2739
rect 19563 2739 19575 2740
rect 19609 2740 19767 2773
rect 19609 2739 19621 2740
rect 19563 2733 19621 2739
rect 19755 2739 19767 2740
rect 19801 2740 19959 2773
rect 19801 2739 19813 2740
rect 19755 2733 19813 2739
rect 19947 2739 19959 2740
rect 19993 2740 20010 2773
rect 19993 2739 20005 2740
rect 19947 2733 20005 2739
rect 18636 2696 18682 2708
rect 18436 2680 18570 2691
rect 18636 2680 18642 2696
rect 18040 2500 18060 2680
rect 18240 2679 18642 2680
rect 18240 2670 18442 2679
rect 18240 2540 18300 2670
rect 18360 2540 18442 2670
rect 18240 2530 18442 2540
rect 18240 2500 18260 2530
rect 18420 2520 18442 2530
rect 18050 2490 18250 2500
rect 18436 2191 18442 2520
rect 18476 2520 18530 2679
rect 18476 2191 18482 2520
rect 18436 2179 18482 2191
rect 18524 2191 18530 2520
rect 18564 2530 18642 2679
rect 18564 2191 18570 2530
rect 18636 2520 18642 2530
rect 18676 2520 18682 2696
rect 18636 2508 18682 2520
rect 18724 2696 18790 2708
rect 18724 2520 18730 2696
rect 18764 2600 18790 2696
rect 20050 2690 20080 3000
rect 20150 2780 20220 2800
rect 20150 2746 20166 2780
rect 20200 2746 20220 2780
rect 20150 2730 20220 2746
rect 20010 2684 20080 2690
rect 18849 2680 18895 2684
rect 19041 2680 19087 2684
rect 19233 2680 19279 2684
rect 19425 2680 19471 2684
rect 19617 2680 19663 2684
rect 19809 2680 19855 2684
rect 20001 2680 20080 2684
rect 18849 2672 20080 2680
rect 18764 2520 18770 2600
rect 18724 2508 18770 2520
rect 18670 2476 18730 2480
rect 18670 2470 18732 2476
rect 18670 2436 18686 2470
rect 18720 2436 18732 2470
rect 18670 2430 18732 2436
rect 18670 2420 18730 2430
rect 18524 2179 18570 2191
rect 17550 1975 18250 2060
rect 18680 1975 18730 2420
rect 18849 2184 18855 2672
rect 18889 2470 19047 2672
rect 18889 2184 18895 2470
rect 18849 2172 18895 2184
rect 18945 2218 18991 2230
rect 18945 2120 18951 2218
rect 17550 1925 18730 1975
rect 18920 2100 18951 2120
rect 18985 2120 18991 2218
rect 19041 2184 19047 2470
rect 19081 2470 19239 2672
rect 19081 2184 19087 2470
rect 19041 2172 19087 2184
rect 19137 2218 19183 2230
rect 19137 2120 19143 2218
rect 18985 2100 19143 2120
rect 18920 2000 18930 2100
rect 19040 2000 19143 2100
rect 18920 1980 18951 2000
rect 18985 1980 19143 2000
rect 16950 1870 17150 1920
rect 16744 1790 17150 1870
rect 17550 1860 18250 1925
rect 16744 1737 16750 1790
rect 15175 1669 15405 1675
rect 16610 1670 16750 1737
rect 15175 1663 15449 1669
rect 15175 1629 15403 1663
rect 15437 1660 15449 1663
rect 15583 1663 15641 1669
rect 15583 1660 15595 1663
rect 15437 1629 15595 1660
rect 15629 1660 15641 1663
rect 15775 1663 15833 1669
rect 15775 1660 15787 1663
rect 15629 1629 15787 1660
rect 15821 1660 15833 1663
rect 15967 1663 16025 1669
rect 15967 1660 15979 1663
rect 15821 1629 15979 1660
rect 16013 1660 16025 1663
rect 16159 1663 16217 1669
rect 16159 1660 16171 1663
rect 16013 1629 16171 1660
rect 16205 1660 16217 1663
rect 16351 1663 16409 1669
rect 16351 1660 16363 1663
rect 16205 1629 16363 1660
rect 16397 1660 16409 1663
rect 16397 1629 16410 1660
rect 16610 1636 16666 1670
rect 16700 1636 16750 1670
rect 16610 1630 16750 1636
rect 15175 1625 16410 1629
rect 15390 1600 16410 1625
rect 16650 1620 16710 1630
rect 16950 1250 17150 1790
rect 18470 1676 18530 1690
rect 18470 1670 18532 1676
rect 18470 1636 18486 1670
rect 18520 1636 18532 1670
rect 18470 1630 18532 1636
rect 18675 1675 18725 1925
rect 18920 1880 18930 1980
rect 19040 1880 19143 1980
rect 18920 1860 18951 1880
rect 18985 1860 19143 1880
rect 18920 1760 18930 1860
rect 19040 1760 19143 1860
rect 18920 1730 18951 1760
rect 18985 1730 19143 1760
rect 19177 2120 19183 2218
rect 19233 2184 19239 2470
rect 19273 2470 19431 2672
rect 19273 2184 19279 2470
rect 19233 2172 19279 2184
rect 19329 2218 19375 2230
rect 19329 2120 19335 2218
rect 19177 1730 19335 2120
rect 19369 2120 19375 2218
rect 19425 2184 19431 2470
rect 19465 2470 19623 2672
rect 19465 2184 19471 2470
rect 19425 2172 19471 2184
rect 19521 2218 19567 2230
rect 19521 2120 19527 2218
rect 19369 1730 19527 2120
rect 19561 2120 19567 2218
rect 19617 2184 19623 2470
rect 19657 2470 19815 2672
rect 19657 2184 19663 2470
rect 19617 2172 19663 2184
rect 19713 2218 19759 2230
rect 19713 2120 19719 2218
rect 19561 1730 19719 2120
rect 19753 2120 19759 2218
rect 19809 2184 19815 2470
rect 19849 2470 20007 2672
rect 19849 2184 19855 2470
rect 19809 2172 19855 2184
rect 19905 2218 19951 2230
rect 19905 2120 19911 2218
rect 19753 1730 19911 2120
rect 19945 1870 19951 2218
rect 20001 2184 20007 2470
rect 20041 2470 20080 2672
rect 20041 2184 20047 2470
rect 20001 2172 20047 2184
rect 20116 2225 20162 2237
rect 20116 1870 20122 2225
rect 19945 1790 20122 1870
rect 19945 1730 19951 1790
rect 18945 1718 18991 1730
rect 19137 1718 19183 1730
rect 19329 1718 19375 1730
rect 19521 1718 19567 1730
rect 19713 1718 19759 1730
rect 19905 1718 19951 1730
rect 20110 1737 20122 1790
rect 20156 1870 20162 2225
rect 20204 2225 20250 2237
rect 20204 1870 20210 2225
rect 20156 1737 20210 1870
rect 20244 1870 20250 2225
rect 21180 2060 21380 9250
rect 22515 6780 22925 6845
rect 22515 6500 22560 6780
rect 22860 6500 22925 6780
rect 22515 5220 22925 6500
rect 23326 6736 23376 6748
rect 23326 6339 23332 6736
rect 23370 6690 23376 6736
rect 23644 6736 23694 6748
rect 23644 6690 23650 6736
rect 23370 6339 23650 6690
rect 23688 6339 23694 6736
rect 23326 6330 23694 6339
rect 23326 6327 23376 6330
rect 23644 6327 23694 6330
rect 23962 6736 24012 6748
rect 23962 6339 23968 6736
rect 24006 6710 24012 6736
rect 24280 6736 24330 6748
rect 24280 6710 24286 6736
rect 24006 6350 24286 6710
rect 24006 6339 24012 6350
rect 23962 6327 24012 6339
rect 24280 6339 24286 6350
rect 24324 6339 24330 6736
rect 24280 6327 24330 6339
rect 23326 5221 23376 5233
rect 23326 5220 23332 5221
rect 22515 4824 23332 5220
rect 23370 4824 23376 5221
rect 22515 4812 23376 4824
rect 23644 5221 23694 5233
rect 23644 4824 23650 5221
rect 23688 5170 23694 5221
rect 23962 5221 24012 5233
rect 23962 5170 23968 5221
rect 23688 4824 23968 5170
rect 24006 4824 24012 5221
rect 24280 5221 24330 5233
rect 24280 4940 24286 5221
rect 23644 4812 24012 4824
rect 24150 4824 24286 4940
rect 24324 4940 24330 5221
rect 24324 4824 24350 4940
rect 22515 4810 23360 4812
rect 23660 4810 23990 4812
rect 22170 4311 22230 4330
rect 22170 4310 22182 4311
rect 22150 4277 22182 4310
rect 22216 4310 22230 4311
rect 22216 4277 22270 4310
rect 22150 4213 22270 4277
rect 22132 4201 22270 4213
rect 22132 3713 22138 4201
rect 22172 4180 22226 4201
rect 22172 3713 22178 4180
rect 22132 3701 22178 3713
rect 22220 3713 22226 4180
rect 22260 4180 22270 4201
rect 22460 4304 23710 4330
rect 22460 4270 22695 4304
rect 22729 4270 22887 4304
rect 22921 4270 23079 4304
rect 23113 4270 23271 4304
rect 23305 4270 23463 4304
rect 23497 4270 23655 4304
rect 23689 4270 23710 4304
rect 23870 4311 23930 4330
rect 23870 4277 23882 4311
rect 23916 4277 23930 4311
rect 23870 4270 23930 4277
rect 22260 3820 22266 4180
rect 22370 3911 22430 3930
rect 22370 3877 22382 3911
rect 22416 3877 22430 3911
rect 22370 3870 22430 3877
rect 22460 3830 22500 4270
rect 22683 4264 22741 4270
rect 22875 4264 22933 4270
rect 23067 4264 23125 4270
rect 23259 4264 23317 4270
rect 23451 4264 23509 4270
rect 23643 4264 23701 4270
rect 23832 4218 23878 4230
rect 22332 3820 22378 3830
rect 22260 3818 22378 3820
rect 22260 3713 22338 3818
rect 21740 3630 21960 3640
rect 21740 3450 21760 3630
rect 21940 3590 21960 3630
rect 22220 3590 22338 3713
rect 21940 3580 22338 3590
rect 21940 3490 22010 3580
rect 22060 3490 22338 3580
rect 21940 3480 22338 3490
rect 21940 3450 21960 3480
rect 21740 3440 21960 3450
rect 22220 3250 22338 3480
rect 22332 3242 22338 3250
rect 22372 3242 22378 3818
rect 22332 3230 22378 3242
rect 22420 3818 22500 3830
rect 22420 3242 22426 3818
rect 22460 3720 22500 3818
rect 22545 4200 22591 4206
rect 22737 4200 22783 4206
rect 22929 4200 22975 4206
rect 23121 4200 23167 4206
rect 23313 4200 23359 4206
rect 23505 4200 23551 4206
rect 23697 4200 23743 4206
rect 22545 4194 23743 4200
rect 22460 3380 22466 3720
rect 22545 3706 22551 4194
rect 22585 4050 22743 4194
rect 22585 3950 22590 4050
rect 22730 3950 22743 4050
rect 22585 3820 22743 3950
rect 22585 3706 22591 3820
rect 22545 3694 22591 3706
rect 22641 3740 22687 3752
rect 22641 3550 22647 3740
rect 22460 3242 22490 3380
rect 22630 3270 22647 3550
rect 22420 3230 22490 3242
rect 22641 3252 22647 3270
rect 22681 3550 22687 3740
rect 22737 3706 22743 3820
rect 22777 3820 22935 4194
rect 22777 3706 22783 3820
rect 22737 3694 22783 3706
rect 22833 3740 22879 3752
rect 22833 3550 22839 3740
rect 22681 3270 22839 3550
rect 22681 3252 22687 3270
rect 22641 3240 22687 3252
rect 22833 3252 22839 3270
rect 22873 3550 22879 3740
rect 22929 3706 22935 3820
rect 22969 3820 23127 4194
rect 22969 3706 22975 3820
rect 22929 3694 22975 3706
rect 23025 3740 23071 3752
rect 23025 3550 23031 3740
rect 22873 3270 23031 3550
rect 22873 3252 22879 3270
rect 22833 3240 22879 3252
rect 23025 3252 23031 3270
rect 23065 3550 23071 3740
rect 23121 3706 23127 3820
rect 23161 3820 23319 4194
rect 23161 3706 23167 3820
rect 23121 3694 23167 3706
rect 23217 3740 23263 3752
rect 23217 3550 23223 3740
rect 23065 3270 23223 3550
rect 23065 3252 23071 3270
rect 23025 3240 23071 3252
rect 23217 3252 23223 3270
rect 23257 3550 23263 3740
rect 23313 3706 23319 3820
rect 23353 3820 23511 4194
rect 23353 3706 23359 3820
rect 23313 3694 23359 3706
rect 23409 3740 23455 3752
rect 23409 3550 23415 3740
rect 23257 3270 23415 3550
rect 23257 3252 23263 3270
rect 23217 3240 23263 3252
rect 23409 3252 23415 3270
rect 23449 3550 23455 3740
rect 23505 3706 23511 3820
rect 23545 3820 23703 4194
rect 23545 3706 23551 3820
rect 23505 3694 23551 3706
rect 23601 3740 23647 3752
rect 23601 3550 23607 3740
rect 23449 3270 23607 3550
rect 23449 3252 23455 3270
rect 23409 3240 23455 3252
rect 23601 3252 23607 3270
rect 23641 3550 23647 3740
rect 23697 3706 23703 3820
rect 23737 3706 23743 4194
rect 23697 3694 23743 3706
rect 23641 3340 23780 3550
rect 23832 3340 23838 4218
rect 23641 3270 23838 3340
rect 23641 3252 23647 3270
rect 23680 3260 23838 3270
rect 23601 3240 23647 3252
rect 23750 3242 23838 3260
rect 23872 3340 23878 4218
rect 23920 4218 23966 4230
rect 23920 3340 23926 4218
rect 23872 3242 23926 3340
rect 23960 3340 23966 4218
rect 23960 3242 23990 3340
rect 22150 3183 22230 3190
rect 22150 3149 22182 3183
rect 22216 3149 22230 3183
rect 22150 3130 22230 3149
rect 22370 3183 22430 3190
rect 22370 3149 22382 3183
rect 22416 3149 22430 3183
rect 22140 2780 22260 2800
rect 22140 2746 22186 2780
rect 22220 2746 22260 2780
rect 21740 2690 21960 2700
rect 22140 2691 22260 2746
rect 22370 2786 22430 3149
rect 22370 2780 22432 2786
rect 22370 2746 22386 2780
rect 22420 2746 22432 2780
rect 22370 2740 22432 2746
rect 22460 2708 22490 3230
rect 22600 3182 23610 3190
rect 22587 3176 23610 3182
rect 22587 3142 22599 3176
rect 22633 3142 22791 3176
rect 22825 3142 22983 3176
rect 23017 3142 23175 3176
rect 23209 3142 23367 3176
rect 23401 3142 23559 3176
rect 23593 3142 23610 3176
rect 22587 3136 23610 3142
rect 22600 3130 23610 3136
rect 23750 3183 23990 3242
rect 23750 3149 23882 3183
rect 23916 3149 23990 3183
rect 23750 3100 23990 3149
rect 24150 3100 24350 4824
rect 23750 3000 24350 3100
rect 22690 2779 23710 2800
rect 22687 2773 23710 2779
rect 22687 2739 22699 2773
rect 22733 2740 22891 2773
rect 22733 2739 22745 2740
rect 22687 2733 22745 2739
rect 22879 2739 22891 2740
rect 22925 2740 23083 2773
rect 22925 2739 22937 2740
rect 22879 2733 22937 2739
rect 23071 2739 23083 2740
rect 23117 2740 23275 2773
rect 23117 2739 23129 2740
rect 23071 2733 23129 2739
rect 23263 2739 23275 2740
rect 23309 2740 23467 2773
rect 23309 2739 23321 2740
rect 23263 2733 23321 2739
rect 23455 2739 23467 2740
rect 23501 2740 23659 2773
rect 23501 2739 23513 2740
rect 23455 2733 23513 2739
rect 23647 2739 23659 2740
rect 23693 2740 23710 2773
rect 23693 2739 23705 2740
rect 23647 2733 23705 2739
rect 22336 2696 22382 2708
rect 21740 2510 21760 2690
rect 21940 2680 21960 2690
rect 22136 2680 22270 2691
rect 22336 2680 22342 2696
rect 21940 2679 22342 2680
rect 21940 2670 22142 2679
rect 21940 2540 22000 2670
rect 22060 2540 22142 2670
rect 21940 2530 22142 2540
rect 21940 2510 21960 2530
rect 22120 2520 22142 2530
rect 21740 2500 21960 2510
rect 22136 2191 22142 2520
rect 22176 2520 22230 2679
rect 22176 2191 22182 2520
rect 22136 2179 22182 2191
rect 22224 2191 22230 2520
rect 22264 2530 22342 2679
rect 22264 2191 22270 2530
rect 22336 2520 22342 2530
rect 22376 2520 22382 2696
rect 22336 2508 22382 2520
rect 22424 2696 22490 2708
rect 22424 2520 22430 2696
rect 22464 2600 22490 2696
rect 23750 2690 23780 3000
rect 23850 2780 23920 2800
rect 23850 2746 23866 2780
rect 23900 2746 23920 2780
rect 23850 2730 23920 2746
rect 23710 2684 23780 2690
rect 22549 2680 22595 2684
rect 22741 2680 22787 2684
rect 22933 2680 22979 2684
rect 23125 2680 23171 2684
rect 23317 2680 23363 2684
rect 23509 2680 23555 2684
rect 23701 2680 23780 2684
rect 22549 2672 23780 2680
rect 22464 2520 22470 2600
rect 22424 2508 22470 2520
rect 22370 2476 22430 2480
rect 22370 2470 22432 2476
rect 22370 2436 22386 2470
rect 22420 2436 22432 2470
rect 22370 2430 22432 2436
rect 22370 2420 22430 2430
rect 22224 2179 22270 2191
rect 21180 1975 21950 2060
rect 22380 1975 22430 2420
rect 22549 2184 22555 2672
rect 22589 2470 22747 2672
rect 22589 2184 22595 2470
rect 22549 2172 22595 2184
rect 22645 2218 22691 2230
rect 22645 2120 22651 2218
rect 21180 1925 22430 1975
rect 22620 2100 22651 2120
rect 22685 2120 22691 2218
rect 22741 2184 22747 2470
rect 22781 2470 22939 2672
rect 22781 2184 22787 2470
rect 22741 2172 22787 2184
rect 22837 2218 22883 2230
rect 22837 2120 22843 2218
rect 22685 2100 22843 2120
rect 22620 2000 22630 2100
rect 22740 2000 22843 2100
rect 22620 1980 22651 2000
rect 22685 1980 22843 2000
rect 20450 1870 20650 1920
rect 20244 1790 20650 1870
rect 21180 1860 21950 1925
rect 20244 1737 20250 1790
rect 18675 1669 18905 1675
rect 20110 1670 20250 1737
rect 18675 1663 18949 1669
rect 18675 1629 18903 1663
rect 18937 1660 18949 1663
rect 19083 1663 19141 1669
rect 19083 1660 19095 1663
rect 18937 1629 19095 1660
rect 19129 1660 19141 1663
rect 19275 1663 19333 1669
rect 19275 1660 19287 1663
rect 19129 1629 19287 1660
rect 19321 1660 19333 1663
rect 19467 1663 19525 1669
rect 19467 1660 19479 1663
rect 19321 1629 19479 1660
rect 19513 1660 19525 1663
rect 19659 1663 19717 1669
rect 19659 1660 19671 1663
rect 19513 1629 19671 1660
rect 19705 1660 19717 1663
rect 19851 1663 19909 1669
rect 19851 1660 19863 1663
rect 19705 1629 19863 1660
rect 19897 1660 19909 1663
rect 19897 1629 19910 1660
rect 20110 1636 20166 1670
rect 20200 1636 20250 1670
rect 20110 1630 20250 1636
rect 18675 1625 19910 1629
rect 18890 1600 19910 1625
rect 20150 1620 20210 1630
rect 20450 1250 20650 1790
rect 22170 1676 22230 1690
rect 22170 1670 22232 1676
rect 22170 1636 22186 1670
rect 22220 1636 22232 1670
rect 22170 1630 22232 1636
rect 22375 1675 22425 1925
rect 22620 1880 22630 1980
rect 22740 1880 22843 1980
rect 22620 1860 22651 1880
rect 22685 1860 22843 1880
rect 22620 1760 22630 1860
rect 22740 1760 22843 1860
rect 22620 1730 22651 1760
rect 22685 1730 22843 1760
rect 22877 2120 22883 2218
rect 22933 2184 22939 2470
rect 22973 2470 23131 2672
rect 22973 2184 22979 2470
rect 22933 2172 22979 2184
rect 23029 2218 23075 2230
rect 23029 2120 23035 2218
rect 22877 1730 23035 2120
rect 23069 2120 23075 2218
rect 23125 2184 23131 2470
rect 23165 2470 23323 2672
rect 23165 2184 23171 2470
rect 23125 2172 23171 2184
rect 23221 2218 23267 2230
rect 23221 2120 23227 2218
rect 23069 1730 23227 2120
rect 23261 2120 23267 2218
rect 23317 2184 23323 2470
rect 23357 2470 23515 2672
rect 23357 2184 23363 2470
rect 23317 2172 23363 2184
rect 23413 2218 23459 2230
rect 23413 2120 23419 2218
rect 23261 1730 23419 2120
rect 23453 2120 23459 2218
rect 23509 2184 23515 2470
rect 23549 2470 23707 2672
rect 23549 2184 23555 2470
rect 23509 2172 23555 2184
rect 23605 2218 23651 2230
rect 23605 2120 23611 2218
rect 23453 1730 23611 2120
rect 23645 1870 23651 2218
rect 23701 2184 23707 2470
rect 23741 2470 23780 2672
rect 23741 2184 23747 2470
rect 23701 2172 23747 2184
rect 23816 2225 23862 2237
rect 23816 1870 23822 2225
rect 23645 1790 23822 1870
rect 23645 1730 23651 1790
rect 22645 1718 22691 1730
rect 22837 1718 22883 1730
rect 23029 1718 23075 1730
rect 23221 1718 23267 1730
rect 23413 1718 23459 1730
rect 23605 1718 23651 1730
rect 23810 1737 23822 1790
rect 23856 1870 23862 2225
rect 23904 2225 23950 2237
rect 23904 1870 23910 2225
rect 23856 1737 23910 1870
rect 23944 1870 23950 2225
rect 24710 2060 24910 10000
rect 25856 9076 25906 9088
rect 25856 8679 25862 9076
rect 25900 9070 25906 9076
rect 26174 9076 26224 9088
rect 26174 9070 26180 9076
rect 25900 8700 26180 9070
rect 25900 8679 25906 8700
rect 25856 8667 25906 8679
rect 26174 8679 26180 8700
rect 26218 8679 26224 9076
rect 26174 8667 26224 8679
rect 26492 9076 26542 9088
rect 26492 8679 26498 9076
rect 26536 9060 26542 9076
rect 26810 9076 26860 9088
rect 26810 9060 26816 9076
rect 26536 8690 26816 9060
rect 26536 8679 26542 8690
rect 26492 8667 26542 8679
rect 26810 8679 26816 8690
rect 26854 8679 26860 9076
rect 26810 8667 26860 8679
rect 27128 9076 27178 9088
rect 27128 8679 27134 9076
rect 27172 9060 27178 9076
rect 27446 9076 27496 9088
rect 27446 9060 27452 9076
rect 27172 8690 27452 9060
rect 27172 8679 27178 8690
rect 27128 8667 27178 8679
rect 27446 8679 27452 8690
rect 27490 8679 27496 9076
rect 27764 9076 27814 9088
rect 27764 9060 27770 9076
rect 27760 8690 27770 9060
rect 27446 8667 27496 8679
rect 27764 8679 27770 8690
rect 27808 9060 27814 9076
rect 28082 9076 28132 9088
rect 28082 9060 28088 9076
rect 27808 8690 28088 9060
rect 27808 8679 27814 8690
rect 27764 8667 27814 8679
rect 28082 8679 28088 8690
rect 28126 8679 28132 9076
rect 28082 8667 28132 8679
rect 25856 7561 25906 7573
rect 25856 7550 25862 7561
rect 25165 7540 25862 7550
rect 25165 7410 25210 7540
rect 25340 7530 25862 7540
rect 25340 7410 25410 7530
rect 25165 7400 25410 7410
rect 25540 7520 25862 7530
rect 25540 7400 25600 7520
rect 25165 7390 25600 7400
rect 25730 7390 25862 7520
rect 25165 7360 25862 7390
rect 25165 7230 25220 7360
rect 25350 7340 25862 7360
rect 25350 7230 25400 7340
rect 25165 7210 25400 7230
rect 25530 7330 25862 7340
rect 25530 7210 25580 7330
rect 25165 7200 25580 7210
rect 25710 7200 25862 7330
rect 25165 7164 25862 7200
rect 25900 7550 25906 7561
rect 26174 7561 26224 7573
rect 25900 7164 25930 7550
rect 25165 7140 25930 7164
rect 26174 7164 26180 7561
rect 26218 7550 26224 7561
rect 26492 7561 26542 7573
rect 26492 7550 26498 7561
rect 26218 7180 26498 7550
rect 26218 7164 26224 7180
rect 26174 7152 26224 7164
rect 26492 7164 26498 7180
rect 26536 7164 26542 7561
rect 26492 7152 26542 7164
rect 26810 7561 26860 7573
rect 26810 7164 26816 7561
rect 26854 7530 26860 7561
rect 27128 7561 27178 7573
rect 27128 7530 27134 7561
rect 26854 7164 27134 7530
rect 27172 7164 27178 7561
rect 26810 7160 27178 7164
rect 26810 7152 26860 7160
rect 27128 7152 27178 7160
rect 27446 7561 27496 7573
rect 27446 7164 27452 7561
rect 27490 7530 27496 7561
rect 27764 7561 27814 7573
rect 27764 7530 27770 7561
rect 27490 7164 27770 7530
rect 27808 7164 27814 7561
rect 28082 7561 28132 7573
rect 28082 7520 28088 7561
rect 27446 7160 27814 7164
rect 27446 7152 27496 7160
rect 27764 7152 27814 7160
rect 28050 7164 28088 7520
rect 28126 7520 28132 7561
rect 28630 7520 28900 7530
rect 28126 7164 28900 7520
rect 28050 7120 28900 7164
rect 28630 6870 28900 7120
rect 28330 6850 28900 6870
rect 25125 6710 25555 6775
rect 25125 6490 25170 6710
rect 25500 6490 25555 6710
rect 25125 5240 25555 6490
rect 25826 6736 25876 6748
rect 25826 6339 25832 6736
rect 25870 6720 25876 6736
rect 26144 6736 26194 6748
rect 26144 6720 26150 6736
rect 25870 6360 26150 6720
rect 25870 6339 25876 6360
rect 25826 6327 25876 6339
rect 26144 6339 26150 6360
rect 26188 6339 26194 6736
rect 26144 6327 26194 6339
rect 26462 6736 26512 6748
rect 26462 6339 26468 6736
rect 26506 6700 26512 6736
rect 26780 6736 26830 6748
rect 26780 6700 26786 6736
rect 26506 6340 26786 6700
rect 26506 6339 26512 6340
rect 26462 6327 26512 6339
rect 26780 6339 26786 6340
rect 26824 6339 26830 6736
rect 26780 6327 26830 6339
rect 27098 6740 27148 6748
rect 27416 6740 27466 6748
rect 27098 6736 27466 6740
rect 27098 6339 27104 6736
rect 27142 6340 27422 6736
rect 27142 6339 27148 6340
rect 27098 6327 27148 6339
rect 27416 6339 27422 6340
rect 27460 6339 27466 6736
rect 27416 6327 27466 6339
rect 27734 6740 27784 6748
rect 28052 6740 28102 6748
rect 27734 6736 28102 6740
rect 27734 6339 27740 6736
rect 27778 6340 28058 6736
rect 27778 6339 27784 6340
rect 27734 6327 27784 6339
rect 28052 6339 28058 6340
rect 28096 6339 28102 6736
rect 28330 6520 28380 6850
rect 28590 6520 28900 6850
rect 28330 6480 28900 6520
rect 28052 6327 28102 6339
rect 28700 5760 28900 6480
rect 29200 6110 29400 9640
rect 32050 7320 32250 7540
rect 32050 7180 32080 7320
rect 32230 7180 32250 7320
rect 32050 7170 32250 7180
rect 32100 7070 32220 7170
rect 29720 7050 34680 7070
rect 29720 7010 29780 7050
rect 30380 7010 34680 7050
rect 29720 6990 34680 7010
rect 29720 6950 34690 6990
rect 29760 6831 30050 6950
rect 29760 6797 29830 6831
rect 29998 6797 30050 6831
rect 29760 6750 30050 6797
rect 29760 6738 30066 6750
rect 29760 6670 29768 6738
rect 29762 6162 29768 6670
rect 29802 6670 30026 6738
rect 29802 6162 29808 6670
rect 29762 6150 29808 6162
rect 30020 6162 30026 6670
rect 30060 6162 30066 6738
rect 30120 6733 30160 6950
rect 30198 6831 30390 6837
rect 30198 6797 30210 6831
rect 30378 6797 30390 6831
rect 30198 6791 30390 6797
rect 30456 6831 30648 6837
rect 30456 6797 30468 6831
rect 30636 6797 30648 6831
rect 30456 6791 30648 6797
rect 30760 6733 30800 6950
rect 30838 6831 31030 6837
rect 30838 6797 30850 6831
rect 31018 6797 31030 6831
rect 30838 6791 31030 6797
rect 31096 6831 31288 6837
rect 31096 6797 31108 6831
rect 31276 6797 31288 6831
rect 31096 6791 31288 6797
rect 31354 6831 31546 6837
rect 31354 6797 31366 6831
rect 31534 6797 31546 6831
rect 31354 6791 31546 6797
rect 31660 6733 31700 6950
rect 31738 6831 31930 6837
rect 31738 6797 31750 6831
rect 31918 6797 31930 6831
rect 31738 6791 31930 6797
rect 31996 6831 32188 6837
rect 31996 6797 32008 6831
rect 32176 6797 32188 6831
rect 31996 6791 32188 6797
rect 32254 6831 32446 6837
rect 32254 6797 32266 6831
rect 32434 6797 32446 6831
rect 32254 6791 32446 6797
rect 32512 6831 32704 6837
rect 32512 6797 32524 6831
rect 32692 6797 32704 6831
rect 32512 6791 32704 6797
rect 32770 6831 32962 6837
rect 32770 6797 32782 6831
rect 32950 6797 32962 6831
rect 32770 6791 32962 6797
rect 33028 6831 33220 6837
rect 33028 6797 33040 6831
rect 33208 6797 33220 6831
rect 33028 6791 33220 6797
rect 33286 6831 33478 6837
rect 33286 6797 33298 6831
rect 33466 6797 33478 6831
rect 33286 6791 33478 6797
rect 33544 6831 33736 6837
rect 33544 6797 33556 6831
rect 33724 6797 33736 6831
rect 33544 6791 33736 6797
rect 33802 6831 33994 6837
rect 33802 6797 33814 6831
rect 33982 6797 33994 6831
rect 33802 6791 33994 6797
rect 34060 6831 34252 6837
rect 34060 6797 34072 6831
rect 34240 6797 34252 6831
rect 34060 6791 34252 6797
rect 34380 6831 34690 6950
rect 34380 6797 34450 6831
rect 34618 6797 34690 6831
rect 34380 6738 34690 6797
rect 30120 6721 30188 6733
rect 30120 6570 30148 6721
rect 30142 6433 30148 6570
rect 30182 6690 30188 6721
rect 30658 6721 30704 6733
rect 30658 6690 30664 6721
rect 30182 6570 30664 6690
rect 30182 6433 30188 6570
rect 30142 6421 30188 6433
rect 30400 6467 30446 6479
rect 30020 6150 30066 6162
rect 30400 6179 30406 6467
rect 30440 6179 30446 6467
rect 30658 6433 30664 6570
rect 30698 6433 30704 6721
rect 30760 6721 30828 6733
rect 30760 6590 30788 6721
rect 30658 6421 30704 6433
rect 30782 6433 30788 6590
rect 30822 6710 30828 6721
rect 31298 6721 31344 6733
rect 31298 6710 31304 6721
rect 30822 6590 31304 6710
rect 30822 6433 30828 6590
rect 30782 6421 30828 6433
rect 31040 6467 31086 6479
rect 30400 6167 30446 6179
rect 31040 6179 31046 6467
rect 31080 6330 31086 6467
rect 31298 6433 31304 6590
rect 31338 6710 31344 6721
rect 31660 6721 31728 6733
rect 31338 6590 31360 6710
rect 31660 6610 31688 6721
rect 31338 6433 31344 6590
rect 31298 6421 31344 6433
rect 31556 6467 31602 6479
rect 31556 6330 31562 6467
rect 31080 6290 31562 6330
rect 31080 6210 31260 6290
rect 31340 6210 31562 6290
rect 31080 6179 31562 6210
rect 31596 6179 31602 6467
rect 31682 6433 31688 6610
rect 31722 6710 31728 6721
rect 32198 6721 32244 6733
rect 32198 6710 32204 6721
rect 31722 6610 32204 6710
rect 31722 6433 31728 6610
rect 31682 6421 31728 6433
rect 31940 6467 31986 6479
rect 31940 6300 31946 6467
rect 31920 6190 31946 6300
rect 31040 6170 31602 6179
rect 31040 6167 31086 6170
rect 31556 6167 31602 6170
rect 31940 6179 31946 6190
rect 31980 6300 31986 6467
rect 32198 6433 32204 6610
rect 32238 6710 32244 6721
rect 32714 6721 32760 6733
rect 32714 6710 32720 6721
rect 32238 6610 32720 6710
rect 32238 6433 32244 6610
rect 32198 6421 32244 6433
rect 32456 6467 32502 6479
rect 32456 6300 32462 6467
rect 31980 6190 32462 6300
rect 31980 6179 31986 6190
rect 31940 6167 31986 6179
rect 32456 6179 32462 6190
rect 32496 6300 32502 6467
rect 32714 6433 32720 6610
rect 32754 6710 32760 6721
rect 33230 6721 33276 6733
rect 33230 6710 33236 6721
rect 32754 6610 33236 6710
rect 32754 6433 32760 6610
rect 32714 6421 32760 6433
rect 32972 6467 33018 6479
rect 32972 6300 32978 6467
rect 32496 6190 32978 6300
rect 32496 6179 32502 6190
rect 32456 6167 32502 6179
rect 32972 6179 32978 6190
rect 33012 6300 33018 6467
rect 33230 6433 33236 6610
rect 33270 6710 33276 6721
rect 33746 6721 33792 6733
rect 33746 6710 33752 6721
rect 33270 6610 33752 6710
rect 33270 6433 33276 6610
rect 33230 6421 33276 6433
rect 33488 6467 33534 6479
rect 33488 6300 33494 6467
rect 33012 6190 33494 6300
rect 33012 6179 33018 6190
rect 32972 6167 33018 6179
rect 33488 6179 33494 6190
rect 33528 6300 33534 6467
rect 33746 6433 33752 6610
rect 33786 6710 33792 6721
rect 34262 6721 34308 6733
rect 34262 6710 34268 6721
rect 33786 6610 34268 6710
rect 33786 6433 33792 6610
rect 33746 6421 33792 6433
rect 34004 6467 34050 6479
rect 33830 6360 33960 6380
rect 33830 6300 33850 6360
rect 33528 6200 33850 6300
rect 33950 6300 33960 6360
rect 34004 6300 34010 6467
rect 33950 6200 34010 6300
rect 33528 6190 34010 6200
rect 33528 6179 33534 6190
rect 33488 6167 33534 6179
rect 34004 6179 34010 6190
rect 34044 6179 34050 6467
rect 34262 6433 34268 6610
rect 34302 6433 34308 6721
rect 34380 6630 34388 6738
rect 34262 6421 34308 6433
rect 34004 6167 34050 6179
rect 30400 6110 30440 6167
rect 34382 6162 34388 6630
rect 34422 6630 34646 6738
rect 34422 6162 34428 6630
rect 34382 6150 34428 6162
rect 34640 6162 34646 6630
rect 34680 6630 34690 6738
rect 34680 6162 34686 6630
rect 34640 6150 34686 6162
rect 29200 6050 29770 6110
rect 29818 6103 30010 6109
rect 29818 6069 29830 6103
rect 29998 6069 30010 6103
rect 29818 6063 30010 6069
rect 30070 6103 34280 6110
rect 30070 6069 30210 6103
rect 30378 6069 30468 6103
rect 30636 6069 30850 6103
rect 31018 6069 31108 6103
rect 31276 6069 31366 6103
rect 31534 6069 31750 6103
rect 31918 6069 32008 6103
rect 32176 6069 32266 6103
rect 32434 6069 32524 6103
rect 32692 6069 32782 6103
rect 32950 6069 33040 6103
rect 33208 6069 33298 6103
rect 33466 6069 33556 6103
rect 33724 6069 33814 6103
rect 33982 6069 34072 6103
rect 34240 6069 34280 6103
rect 29200 5990 29400 6050
rect 29710 6030 29770 6050
rect 30070 6050 34280 6069
rect 34438 6103 34630 6109
rect 34438 6069 34450 6103
rect 34618 6069 34630 6103
rect 34438 6063 34630 6069
rect 30070 6030 30130 6050
rect 29710 5970 30130 6030
rect 35030 5990 35230 6000
rect 29470 5870 30440 5940
rect 28700 5690 29410 5760
rect 29470 5690 29520 5870
rect 30060 5820 30120 5830
rect 28700 5620 29520 5690
rect 30020 5811 30150 5820
rect 30020 5777 30072 5811
rect 30106 5777 30150 5811
rect 30370 5811 30440 5870
rect 30370 5780 30392 5811
rect 30020 5713 30150 5777
rect 30380 5777 30392 5780
rect 30426 5777 30440 5811
rect 30380 5770 30440 5777
rect 30560 5930 30660 5950
rect 35030 5930 35630 5990
rect 30560 5850 30580 5930
rect 30640 5850 30660 5930
rect 30020 5701 30156 5713
rect 30020 5660 30028 5701
rect 28700 5560 29410 5620
rect 30022 5413 30028 5660
rect 30062 5660 30116 5701
rect 30062 5413 30068 5660
rect 30022 5401 30068 5413
rect 30110 5413 30116 5660
rect 30150 5670 30156 5701
rect 30242 5701 30288 5713
rect 30242 5670 30248 5701
rect 30150 5550 30248 5670
rect 30150 5413 30156 5550
rect 30110 5401 30156 5413
rect 30242 5413 30248 5550
rect 30282 5690 30288 5701
rect 30434 5701 30480 5713
rect 30434 5690 30440 5701
rect 30282 5530 30440 5690
rect 30282 5413 30288 5530
rect 30242 5401 30288 5413
rect 30338 5447 30384 5459
rect 25125 5233 25870 5240
rect 25125 5221 25876 5233
rect 25125 4824 25832 5221
rect 25870 4824 25876 5221
rect 25125 4812 25876 4824
rect 26144 5221 26194 5233
rect 26144 4824 26150 5221
rect 26188 5190 26194 5221
rect 26462 5221 26512 5233
rect 26462 5190 26468 5221
rect 26188 4830 26468 5190
rect 26188 4824 26194 4830
rect 26144 4812 26194 4824
rect 26462 4824 26468 4830
rect 26506 4824 26512 5221
rect 26462 4812 26512 4824
rect 26780 5221 26830 5233
rect 26780 4824 26786 5221
rect 26824 5190 26830 5221
rect 27098 5221 27148 5233
rect 27098 5190 27104 5221
rect 26824 4830 27104 5190
rect 26824 4824 26830 4830
rect 26780 4812 26830 4824
rect 27098 4824 27104 4830
rect 27142 4824 27148 5221
rect 27098 4812 27148 4824
rect 27416 5221 27466 5233
rect 27416 4824 27422 5221
rect 27460 5220 27466 5221
rect 27734 5221 27784 5233
rect 27734 5220 27740 5221
rect 27460 4824 27740 5220
rect 27778 4824 27784 5221
rect 28052 5221 28102 5233
rect 28052 4940 28058 5221
rect 27416 4820 27784 4824
rect 27416 4812 27466 4820
rect 27734 4812 27784 4820
rect 27950 4824 28058 4940
rect 28096 4940 28102 5221
rect 30338 5159 30344 5447
rect 30378 5290 30384 5447
rect 30434 5413 30440 5530
rect 30474 5690 30480 5701
rect 30560 5690 30660 5850
rect 34905 5910 35630 5930
rect 34905 5830 34920 5910
rect 35010 5830 35630 5910
rect 30780 5811 30840 5830
rect 30780 5777 30792 5811
rect 30826 5777 30840 5811
rect 31080 5811 31140 5830
rect 34905 5820 35630 5830
rect 31080 5810 31092 5811
rect 30780 5770 30840 5777
rect 31070 5777 31092 5810
rect 31126 5810 31140 5811
rect 31126 5777 31150 5810
rect 35030 5800 35630 5820
rect 35430 5790 35630 5800
rect 31070 5713 31150 5777
rect 30738 5701 30784 5713
rect 30738 5690 30744 5701
rect 30474 5530 30744 5690
rect 30474 5413 30480 5530
rect 30434 5401 30480 5413
rect 30530 5447 30576 5459
rect 30530 5290 30536 5447
rect 30378 5159 30536 5290
rect 30570 5159 30576 5447
rect 30338 5150 30576 5159
rect 30338 5147 30420 5150
rect 30530 5147 30576 5150
rect 30642 5447 30688 5459
rect 30642 5159 30648 5447
rect 30682 5290 30688 5447
rect 30738 5413 30744 5530
rect 30778 5690 30784 5701
rect 30930 5701 30976 5713
rect 30930 5690 30936 5701
rect 30778 5530 30936 5690
rect 30778 5413 30784 5530
rect 30738 5401 30784 5413
rect 30834 5447 30880 5459
rect 30834 5290 30840 5447
rect 30682 5159 30840 5290
rect 30874 5159 30880 5447
rect 30930 5413 30936 5530
rect 30970 5680 30976 5701
rect 31042 5701 31176 5713
rect 31042 5680 31048 5701
rect 30970 5530 31048 5680
rect 30970 5413 30976 5530
rect 30930 5401 30976 5413
rect 31042 5413 31048 5530
rect 31082 5530 31136 5701
rect 31082 5413 31088 5530
rect 31042 5401 31088 5413
rect 31130 5413 31136 5530
rect 31170 5680 31176 5701
rect 31170 5530 31180 5680
rect 31170 5413 31176 5530
rect 31130 5401 31176 5413
rect 30642 5147 30880 5159
rect 30060 5083 30120 5090
rect 30060 5049 30072 5083
rect 30106 5049 30120 5083
rect 30060 5030 30120 5049
rect 30280 5089 30340 5090
rect 30280 5083 30342 5089
rect 30280 5049 30296 5083
rect 30330 5049 30342 5083
rect 30280 5043 30342 5049
rect 30280 5030 30340 5043
rect 28096 4824 28150 4940
rect 25125 4810 25870 4812
rect 25970 4311 26030 4330
rect 25970 4310 25982 4311
rect 25950 4277 25982 4310
rect 26016 4310 26030 4311
rect 26016 4277 26070 4310
rect 25950 4213 26070 4277
rect 25932 4201 26070 4213
rect 25932 3713 25938 4201
rect 25972 4180 26026 4201
rect 25972 3713 25978 4180
rect 25932 3701 25978 3713
rect 26020 3713 26026 4180
rect 26060 4180 26070 4201
rect 26260 4304 27510 4330
rect 26260 4270 26495 4304
rect 26529 4270 26687 4304
rect 26721 4270 26879 4304
rect 26913 4270 27071 4304
rect 27105 4270 27263 4304
rect 27297 4270 27455 4304
rect 27489 4270 27510 4304
rect 27670 4311 27730 4330
rect 27670 4277 27682 4311
rect 27716 4277 27730 4311
rect 27670 4270 27730 4277
rect 26060 3820 26066 4180
rect 26170 3911 26230 3930
rect 26170 3877 26182 3911
rect 26216 3877 26230 3911
rect 26170 3870 26230 3877
rect 26260 3830 26300 4270
rect 26483 4264 26541 4270
rect 26675 4264 26733 4270
rect 26867 4264 26925 4270
rect 27059 4264 27117 4270
rect 27251 4264 27309 4270
rect 27443 4264 27501 4270
rect 27632 4218 27678 4230
rect 26132 3820 26178 3830
rect 26060 3818 26178 3820
rect 26060 3713 26138 3818
rect 25540 3630 25760 3640
rect 25540 3450 25560 3630
rect 25740 3590 25760 3630
rect 26020 3590 26138 3713
rect 25740 3580 26138 3590
rect 25740 3490 25810 3580
rect 25860 3490 26138 3580
rect 25740 3480 26138 3490
rect 25740 3450 25760 3480
rect 25540 3440 25760 3450
rect 26020 3250 26138 3480
rect 26132 3242 26138 3250
rect 26172 3242 26178 3818
rect 26132 3230 26178 3242
rect 26220 3818 26300 3830
rect 26220 3242 26226 3818
rect 26260 3720 26300 3818
rect 26345 4200 26391 4206
rect 26537 4200 26583 4206
rect 26729 4200 26775 4206
rect 26921 4200 26967 4206
rect 27113 4200 27159 4206
rect 27305 4200 27351 4206
rect 27497 4200 27543 4206
rect 26345 4194 27543 4200
rect 26260 3380 26266 3720
rect 26345 3706 26351 4194
rect 26385 4050 26543 4194
rect 26385 3950 26390 4050
rect 26530 3950 26543 4050
rect 26385 3820 26543 3950
rect 26385 3706 26391 3820
rect 26345 3694 26391 3706
rect 26441 3740 26487 3752
rect 26441 3550 26447 3740
rect 26260 3242 26290 3380
rect 26430 3270 26447 3550
rect 26220 3230 26290 3242
rect 26441 3252 26447 3270
rect 26481 3550 26487 3740
rect 26537 3706 26543 3820
rect 26577 3820 26735 4194
rect 26577 3706 26583 3820
rect 26537 3694 26583 3706
rect 26633 3740 26679 3752
rect 26633 3550 26639 3740
rect 26481 3270 26639 3550
rect 26481 3252 26487 3270
rect 26441 3240 26487 3252
rect 26633 3252 26639 3270
rect 26673 3550 26679 3740
rect 26729 3706 26735 3820
rect 26769 3820 26927 4194
rect 26769 3706 26775 3820
rect 26729 3694 26775 3706
rect 26825 3740 26871 3752
rect 26825 3550 26831 3740
rect 26673 3270 26831 3550
rect 26673 3252 26679 3270
rect 26633 3240 26679 3252
rect 26825 3252 26831 3270
rect 26865 3550 26871 3740
rect 26921 3706 26927 3820
rect 26961 3820 27119 4194
rect 26961 3706 26967 3820
rect 26921 3694 26967 3706
rect 27017 3740 27063 3752
rect 27017 3550 27023 3740
rect 26865 3270 27023 3550
rect 26865 3252 26871 3270
rect 26825 3240 26871 3252
rect 27017 3252 27023 3270
rect 27057 3550 27063 3740
rect 27113 3706 27119 3820
rect 27153 3820 27311 4194
rect 27153 3706 27159 3820
rect 27113 3694 27159 3706
rect 27209 3740 27255 3752
rect 27209 3550 27215 3740
rect 27057 3270 27215 3550
rect 27057 3252 27063 3270
rect 27017 3240 27063 3252
rect 27209 3252 27215 3270
rect 27249 3550 27255 3740
rect 27305 3706 27311 3820
rect 27345 3820 27503 4194
rect 27345 3706 27351 3820
rect 27305 3694 27351 3706
rect 27401 3740 27447 3752
rect 27401 3550 27407 3740
rect 27249 3270 27407 3550
rect 27249 3252 27255 3270
rect 27209 3240 27255 3252
rect 27401 3252 27407 3270
rect 27441 3550 27447 3740
rect 27497 3706 27503 3820
rect 27537 3706 27543 4194
rect 27497 3694 27543 3706
rect 27441 3340 27580 3550
rect 27632 3340 27638 4218
rect 27441 3270 27638 3340
rect 27441 3252 27447 3270
rect 27480 3260 27638 3270
rect 27401 3240 27447 3252
rect 27550 3242 27638 3260
rect 27672 3340 27678 4218
rect 27720 4218 27766 4230
rect 27720 3340 27726 4218
rect 27672 3242 27726 3340
rect 27760 3340 27766 4218
rect 27760 3242 27790 3340
rect 25950 3183 26030 3190
rect 25950 3149 25982 3183
rect 26016 3149 26030 3183
rect 25950 3130 26030 3149
rect 26170 3183 26230 3190
rect 26170 3149 26182 3183
rect 26216 3149 26230 3183
rect 25940 2780 26060 2800
rect 25940 2746 25986 2780
rect 26020 2746 26060 2780
rect 25540 2690 25760 2700
rect 25940 2691 26060 2746
rect 26170 2786 26230 3149
rect 26170 2780 26232 2786
rect 26170 2746 26186 2780
rect 26220 2746 26232 2780
rect 26170 2740 26232 2746
rect 26260 2708 26290 3230
rect 26400 3182 27410 3190
rect 26387 3176 27410 3182
rect 26387 3142 26399 3176
rect 26433 3142 26591 3176
rect 26625 3142 26783 3176
rect 26817 3142 26975 3176
rect 27009 3142 27167 3176
rect 27201 3142 27359 3176
rect 27393 3142 27410 3176
rect 26387 3136 27410 3142
rect 26400 3130 27410 3136
rect 27550 3183 27790 3242
rect 27550 3149 27682 3183
rect 27716 3149 27790 3183
rect 27550 3100 27790 3149
rect 27950 3100 28150 4824
rect 27550 3000 28150 3100
rect 28700 4870 29410 4920
rect 29480 4870 29560 4880
rect 28700 4820 29490 4870
rect 28700 4720 29410 4820
rect 29480 4810 29490 4820
rect 29550 4810 29560 4870
rect 30380 4830 30420 5147
rect 30660 5130 30880 5147
rect 30480 5089 30540 5090
rect 30476 5083 30540 5089
rect 30476 5049 30488 5083
rect 30522 5049 30540 5083
rect 30476 5043 30540 5049
rect 30480 5030 30540 5043
rect 30670 5083 30750 5090
rect 30670 5080 30696 5083
rect 30730 5080 30750 5083
rect 30670 5020 30680 5080
rect 30740 5020 30750 5080
rect 30670 5010 30750 5020
rect 29480 4800 29560 4810
rect 30220 4790 30420 4830
rect 30780 4830 30820 5130
rect 30880 5089 30940 5090
rect 30876 5083 30940 5089
rect 30876 5049 30888 5083
rect 30922 5049 30940 5083
rect 30876 5043 30940 5049
rect 30880 5030 30940 5043
rect 31080 5083 31140 5090
rect 31080 5049 31092 5083
rect 31126 5049 31140 5083
rect 31080 5030 31140 5049
rect 30780 4790 30980 4830
rect 26490 2779 27510 2800
rect 26487 2773 27510 2779
rect 26487 2739 26499 2773
rect 26533 2740 26691 2773
rect 26533 2739 26545 2740
rect 26487 2733 26545 2739
rect 26679 2739 26691 2740
rect 26725 2740 26883 2773
rect 26725 2739 26737 2740
rect 26679 2733 26737 2739
rect 26871 2739 26883 2740
rect 26917 2740 27075 2773
rect 26917 2739 26929 2740
rect 26871 2733 26929 2739
rect 27063 2739 27075 2740
rect 27109 2740 27267 2773
rect 27109 2739 27121 2740
rect 27063 2733 27121 2739
rect 27255 2739 27267 2740
rect 27301 2740 27459 2773
rect 27301 2739 27313 2740
rect 27255 2733 27313 2739
rect 27447 2739 27459 2740
rect 27493 2740 27510 2773
rect 27493 2739 27505 2740
rect 27447 2733 27505 2739
rect 26136 2696 26182 2708
rect 25540 2510 25560 2690
rect 25740 2680 25760 2690
rect 25936 2680 26070 2691
rect 26136 2680 26142 2696
rect 25740 2679 26142 2680
rect 25740 2670 25942 2679
rect 25740 2540 25800 2670
rect 25860 2540 25942 2670
rect 25740 2530 25942 2540
rect 25740 2510 25760 2530
rect 25920 2520 25942 2530
rect 25540 2500 25760 2510
rect 25936 2191 25942 2520
rect 25976 2520 26030 2679
rect 25976 2191 25982 2520
rect 25936 2179 25982 2191
rect 26024 2191 26030 2520
rect 26064 2530 26142 2679
rect 26064 2191 26070 2530
rect 26136 2520 26142 2530
rect 26176 2520 26182 2696
rect 26136 2508 26182 2520
rect 26224 2696 26290 2708
rect 26224 2520 26230 2696
rect 26264 2600 26290 2696
rect 27550 2690 27580 3000
rect 27650 2780 27720 2800
rect 27650 2746 27666 2780
rect 27700 2746 27720 2780
rect 27650 2730 27720 2746
rect 27510 2684 27580 2690
rect 26349 2680 26395 2684
rect 26541 2680 26587 2684
rect 26733 2680 26779 2684
rect 26925 2680 26971 2684
rect 27117 2680 27163 2684
rect 27309 2680 27355 2684
rect 27501 2680 27580 2684
rect 26349 2672 27580 2680
rect 26264 2520 26270 2600
rect 26224 2508 26270 2520
rect 26170 2476 26230 2480
rect 26170 2470 26232 2476
rect 26170 2436 26186 2470
rect 26220 2436 26232 2470
rect 26170 2430 26232 2436
rect 26170 2420 26230 2430
rect 26024 2179 26070 2191
rect 24710 1975 25750 2060
rect 26180 1975 26230 2420
rect 26349 2184 26355 2672
rect 26389 2470 26547 2672
rect 26389 2184 26395 2470
rect 26349 2172 26395 2184
rect 26445 2218 26491 2230
rect 26445 2120 26451 2218
rect 24710 1925 26230 1975
rect 26420 2100 26451 2120
rect 26485 2120 26491 2218
rect 26541 2184 26547 2470
rect 26581 2470 26739 2672
rect 26581 2184 26587 2470
rect 26541 2172 26587 2184
rect 26637 2218 26683 2230
rect 26637 2120 26643 2218
rect 26485 2100 26643 2120
rect 26420 2000 26430 2100
rect 26540 2000 26643 2100
rect 26420 1980 26451 2000
rect 26485 1980 26643 2000
rect 24150 1870 24350 1920
rect 23944 1790 24350 1870
rect 24710 1860 25750 1925
rect 23944 1737 23950 1790
rect 22375 1669 22605 1675
rect 23810 1670 23950 1737
rect 22375 1663 22649 1669
rect 22375 1629 22603 1663
rect 22637 1660 22649 1663
rect 22783 1663 22841 1669
rect 22783 1660 22795 1663
rect 22637 1629 22795 1660
rect 22829 1660 22841 1663
rect 22975 1663 23033 1669
rect 22975 1660 22987 1663
rect 22829 1629 22987 1660
rect 23021 1660 23033 1663
rect 23167 1663 23225 1669
rect 23167 1660 23179 1663
rect 23021 1629 23179 1660
rect 23213 1660 23225 1663
rect 23359 1663 23417 1669
rect 23359 1660 23371 1663
rect 23213 1629 23371 1660
rect 23405 1660 23417 1663
rect 23551 1663 23609 1669
rect 23551 1660 23563 1663
rect 23405 1629 23563 1660
rect 23597 1660 23609 1663
rect 23597 1629 23610 1660
rect 23810 1636 23866 1670
rect 23900 1636 23950 1670
rect 23810 1630 23950 1636
rect 22375 1625 23610 1629
rect 22590 1600 23610 1625
rect 23850 1620 23910 1630
rect 24150 1250 24350 1790
rect 25970 1676 26030 1690
rect 25970 1670 26032 1676
rect 25970 1636 25986 1670
rect 26020 1636 26032 1670
rect 25970 1630 26032 1636
rect 26175 1675 26225 1925
rect 26420 1880 26430 1980
rect 26540 1880 26643 1980
rect 26420 1860 26451 1880
rect 26485 1860 26643 1880
rect 26420 1760 26430 1860
rect 26540 1760 26643 1860
rect 26420 1730 26451 1760
rect 26485 1730 26643 1760
rect 26677 2120 26683 2218
rect 26733 2184 26739 2470
rect 26773 2470 26931 2672
rect 26773 2184 26779 2470
rect 26733 2172 26779 2184
rect 26829 2218 26875 2230
rect 26829 2120 26835 2218
rect 26677 1730 26835 2120
rect 26869 2120 26875 2218
rect 26925 2184 26931 2470
rect 26965 2470 27123 2672
rect 26965 2184 26971 2470
rect 26925 2172 26971 2184
rect 27021 2218 27067 2230
rect 27021 2120 27027 2218
rect 26869 1730 27027 2120
rect 27061 2120 27067 2218
rect 27117 2184 27123 2470
rect 27157 2470 27315 2672
rect 27157 2184 27163 2470
rect 27117 2172 27163 2184
rect 27213 2218 27259 2230
rect 27213 2120 27219 2218
rect 27061 1730 27219 2120
rect 27253 2120 27259 2218
rect 27309 2184 27315 2470
rect 27349 2470 27507 2672
rect 27349 2184 27355 2470
rect 27309 2172 27355 2184
rect 27405 2218 27451 2230
rect 27405 2120 27411 2218
rect 27253 1730 27411 2120
rect 27445 1870 27451 2218
rect 27501 2184 27507 2470
rect 27541 2470 27580 2672
rect 27541 2184 27547 2470
rect 27501 2172 27547 2184
rect 27616 2225 27662 2237
rect 27616 1870 27622 2225
rect 27445 1790 27622 1870
rect 27445 1730 27451 1790
rect 26445 1718 26491 1730
rect 26637 1718 26683 1730
rect 26829 1718 26875 1730
rect 27021 1718 27067 1730
rect 27213 1718 27259 1730
rect 27405 1718 27451 1730
rect 27610 1737 27622 1790
rect 27656 1870 27662 2225
rect 27704 2225 27750 2237
rect 27704 1870 27710 2225
rect 27656 1737 27710 1870
rect 27744 1870 27750 2225
rect 27950 1870 28150 1920
rect 27744 1790 28150 1870
rect 27744 1737 27750 1790
rect 26175 1669 26405 1675
rect 27610 1670 27750 1737
rect 26175 1663 26449 1669
rect 26175 1629 26403 1663
rect 26437 1660 26449 1663
rect 26583 1663 26641 1669
rect 26583 1660 26595 1663
rect 26437 1629 26595 1660
rect 26629 1660 26641 1663
rect 26775 1663 26833 1669
rect 26775 1660 26787 1663
rect 26629 1629 26787 1660
rect 26821 1660 26833 1663
rect 26967 1663 27025 1669
rect 26967 1660 26979 1663
rect 26821 1629 26979 1660
rect 27013 1660 27025 1663
rect 27159 1663 27217 1669
rect 27159 1660 27171 1663
rect 27013 1629 27171 1660
rect 27205 1660 27217 1663
rect 27351 1663 27409 1669
rect 27351 1660 27363 1663
rect 27205 1629 27363 1660
rect 27397 1660 27409 1663
rect 27397 1629 27410 1660
rect 27610 1636 27666 1670
rect 27700 1636 27750 1670
rect 27610 1630 27750 1636
rect 26175 1625 27410 1629
rect 26390 1600 27410 1625
rect 27650 1620 27710 1630
rect 27950 1250 28150 1790
rect 3450 1050 28150 1250
rect 14050 -160 14250 1050
rect 28700 -200 28900 4720
rect 29922 4630 30114 4636
rect 29922 4596 29934 4630
rect 30102 4596 30114 4630
rect 29922 4590 30114 4596
rect 30220 4630 30260 4790
rect 30940 4640 30980 4790
rect 30302 4630 30494 4636
rect 30702 4630 30894 4636
rect 30940 4630 33340 4640
rect 30220 4596 30314 4630
rect 30482 4596 30714 4630
rect 30882 4596 30900 4630
rect 30220 4590 30900 4596
rect 30940 4600 31094 4630
rect 30220 4558 30260 4590
rect 30940 4560 30980 4600
rect 31082 4596 31094 4600
rect 31262 4600 31352 4630
rect 31262 4596 31274 4600
rect 31082 4590 31274 4596
rect 31340 4596 31352 4600
rect 31520 4600 31610 4630
rect 31520 4596 31532 4600
rect 31340 4590 31532 4596
rect 31598 4596 31610 4600
rect 31778 4600 31868 4630
rect 31778 4596 31790 4600
rect 31598 4590 31790 4596
rect 31856 4596 31868 4600
rect 32036 4600 32126 4630
rect 32036 4596 32048 4600
rect 31856 4590 32048 4596
rect 32114 4596 32126 4600
rect 32294 4600 32384 4630
rect 32294 4596 32306 4600
rect 32114 4590 32306 4596
rect 32372 4596 32384 4600
rect 32552 4600 32642 4630
rect 32552 4596 32564 4600
rect 32372 4590 32564 4596
rect 32630 4596 32642 4600
rect 32810 4600 32900 4630
rect 32810 4596 32822 4600
rect 32630 4590 32822 4596
rect 32888 4596 32900 4600
rect 33068 4600 33158 4630
rect 33068 4596 33080 4600
rect 32888 4590 33080 4596
rect 33146 4596 33158 4600
rect 33326 4600 33340 4630
rect 33522 4630 33714 4636
rect 33326 4596 33338 4600
rect 33146 4590 33338 4596
rect 33522 4596 33534 4630
rect 33702 4596 33714 4630
rect 33522 4590 33714 4596
rect 30930 4558 30990 4560
rect 29866 4546 29912 4558
rect 29866 4370 29872 4546
rect 29906 4450 29912 4546
rect 30124 4546 30170 4558
rect 30124 4450 30130 4546
rect 29906 4370 30130 4450
rect 30164 4370 30170 4546
rect 30220 4546 30292 4558
rect 30220 4530 30252 4546
rect 30240 4390 30252 4530
rect 29866 4358 30170 4370
rect 30246 4370 30252 4390
rect 30286 4370 30292 4546
rect 30504 4550 30550 4558
rect 30646 4550 30692 4558
rect 30504 4546 30692 4550
rect 30504 4450 30510 4546
rect 30500 4410 30510 4450
rect 30246 4358 30292 4370
rect 30504 4370 30510 4410
rect 30544 4370 30652 4546
rect 30686 4370 30692 4546
rect 30504 4358 30692 4370
rect 30904 4546 30990 4558
rect 30904 4370 30910 4546
rect 30944 4370 30990 4546
rect 31040 4541 33140 4560
rect 31026 4540 33140 4541
rect 31026 4529 32950 4540
rect 31026 4441 31032 4529
rect 31066 4520 31548 4529
rect 31066 4441 31072 4520
rect 31026 4429 31072 4441
rect 31284 4475 31330 4487
rect 31284 4400 31290 4475
rect 30904 4358 30990 4370
rect 31280 4387 31290 4400
rect 31324 4400 31330 4475
rect 31542 4441 31548 4520
rect 31582 4520 32064 4529
rect 31582 4441 31588 4520
rect 31542 4429 31588 4441
rect 31800 4475 31846 4487
rect 31800 4400 31806 4475
rect 31324 4387 31806 4400
rect 31840 4400 31846 4475
rect 32058 4441 32064 4520
rect 32098 4520 32580 4529
rect 32098 4441 32104 4520
rect 32058 4429 32104 4441
rect 32316 4475 32362 4487
rect 32316 4400 32322 4475
rect 31840 4387 32322 4400
rect 32356 4400 32362 4475
rect 32574 4441 32580 4520
rect 32614 4520 32950 4529
rect 32614 4441 32620 4520
rect 32574 4429 32620 4441
rect 32832 4475 32878 4487
rect 32832 4400 32838 4475
rect 32356 4387 32838 4400
rect 32872 4400 32878 4475
rect 32940 4460 32950 4520
rect 33030 4529 33140 4540
rect 33030 4520 33096 4529
rect 33030 4460 33040 4520
rect 32940 4450 33040 4460
rect 33090 4441 33096 4520
rect 33130 4520 33140 4529
rect 33466 4546 33512 4558
rect 33130 4441 33136 4520
rect 33090 4429 33136 4441
rect 33348 4475 33394 4487
rect 33348 4400 33354 4475
rect 32872 4387 33354 4400
rect 33388 4400 33394 4475
rect 33388 4387 33400 4400
rect 31280 4360 33400 4387
rect 29870 4320 30170 4358
rect 30520 4350 30680 4358
rect 29870 4286 29934 4320
rect 30102 4286 30170 4320
rect 29870 4090 30170 4286
rect 30302 4320 30494 4326
rect 30302 4286 30314 4320
rect 30482 4286 30494 4320
rect 30302 4280 30494 4286
rect 29090 3890 29100 4090
rect 29400 4040 29410 4090
rect 29870 4050 29900 4090
rect 30160 4050 30170 4090
rect 29870 4040 30170 4050
rect 30580 4040 30620 4350
rect 30702 4320 30894 4326
rect 30702 4286 30714 4320
rect 30882 4286 30894 4320
rect 30702 4280 30894 4286
rect 30930 4220 30990 4358
rect 31082 4320 31274 4326
rect 31082 4286 31094 4320
rect 31262 4286 31274 4320
rect 31082 4280 31274 4286
rect 31340 4320 31532 4326
rect 31340 4286 31352 4320
rect 31520 4286 31532 4320
rect 31340 4280 31532 4286
rect 31598 4320 31790 4326
rect 31598 4286 31610 4320
rect 31778 4286 31790 4320
rect 31598 4280 31790 4286
rect 31856 4320 32048 4326
rect 31856 4286 31868 4320
rect 32036 4286 32048 4320
rect 31856 4280 32048 4286
rect 32114 4320 32306 4326
rect 32114 4286 32126 4320
rect 32294 4286 32306 4320
rect 32114 4280 32306 4286
rect 32372 4320 32564 4326
rect 32372 4286 32384 4320
rect 32552 4286 32564 4320
rect 32372 4280 32564 4286
rect 32630 4320 32822 4326
rect 32630 4286 32642 4320
rect 32810 4286 32822 4320
rect 32630 4280 32822 4286
rect 32888 4320 33080 4326
rect 32888 4286 32900 4320
rect 33068 4286 33080 4320
rect 32888 4280 33080 4286
rect 33146 4320 33338 4326
rect 33146 4286 33158 4320
rect 33326 4286 33338 4320
rect 33146 4280 33338 4286
rect 30900 4210 31050 4220
rect 30900 4090 30920 4210
rect 31040 4090 31050 4210
rect 30900 4080 31050 4090
rect 33370 4040 33400 4360
rect 33466 4370 33472 4546
rect 33506 4400 33512 4546
rect 33724 4546 33770 4558
rect 33724 4400 33730 4546
rect 33506 4370 33730 4400
rect 33764 4370 33770 4546
rect 33466 4358 33770 4370
rect 33470 4320 33760 4358
rect 33470 4286 33534 4320
rect 33702 4286 33760 4320
rect 33470 4250 33760 4286
rect 33450 4170 33760 4250
rect 33450 4040 33750 4170
rect 29400 3920 33750 4040
rect 29400 3890 29410 3920
rect 29200 3880 29400 3890
<< rmetal1 >>
rect 290 19750 320 19840
<< via1 >>
rect 6043 27425 6095 27434
rect 6107 27425 6159 27434
rect 6043 27391 6081 27425
rect 6081 27391 6095 27425
rect 6107 27391 6115 27425
rect 6115 27391 6159 27425
rect 6043 27382 6095 27391
rect 6107 27382 6159 27391
rect 6171 27425 6223 27434
rect 6171 27391 6173 27425
rect 6173 27391 6207 27425
rect 6207 27391 6223 27425
rect 6171 27382 6223 27391
rect 6235 27425 6287 27434
rect 6235 27391 6265 27425
rect 6265 27391 6287 27425
rect 6235 27382 6287 27391
rect 6299 27382 6351 27434
rect 9861 27425 9913 27434
rect 9861 27391 9887 27425
rect 9887 27391 9913 27425
rect 9861 27382 9913 27391
rect 9925 27425 9977 27434
rect 9989 27425 10041 27434
rect 10053 27425 10105 27434
rect 9925 27391 9945 27425
rect 9945 27391 9977 27425
rect 9989 27391 10037 27425
rect 10037 27391 10041 27425
rect 10053 27391 10071 27425
rect 10071 27391 10105 27425
rect 9925 27382 9977 27391
rect 9989 27382 10041 27391
rect 10053 27382 10105 27391
rect 10117 27425 10169 27434
rect 13679 27425 13731 27434
rect 13743 27425 13795 27434
rect 10117 27391 10129 27425
rect 10129 27391 10163 27425
rect 10163 27391 10169 27425
rect 13679 27391 13717 27425
rect 13717 27391 13731 27425
rect 13743 27391 13751 27425
rect 13751 27391 13795 27425
rect 10117 27382 10169 27391
rect 13679 27382 13731 27391
rect 13743 27382 13795 27391
rect 13807 27425 13859 27434
rect 13807 27391 13809 27425
rect 13809 27391 13843 27425
rect 13843 27391 13859 27425
rect 13807 27382 13859 27391
rect 13871 27425 13923 27434
rect 13871 27391 13901 27425
rect 13901 27391 13923 27425
rect 13871 27382 13923 27391
rect 13935 27382 13987 27434
rect 17497 27425 17549 27434
rect 17497 27391 17523 27425
rect 17523 27391 17549 27425
rect 17497 27382 17549 27391
rect 17561 27425 17613 27434
rect 17625 27425 17677 27434
rect 17689 27425 17741 27434
rect 17561 27391 17581 27425
rect 17581 27391 17613 27425
rect 17625 27391 17673 27425
rect 17673 27391 17677 27425
rect 17689 27391 17707 27425
rect 17707 27391 17741 27425
rect 17561 27382 17613 27391
rect 17625 27382 17677 27391
rect 17689 27382 17741 27391
rect 17753 27425 17805 27434
rect 17753 27391 17765 27425
rect 17765 27391 17799 27425
rect 17799 27391 17805 27425
rect 17753 27382 17805 27391
rect 10212 27280 10264 27332
rect 5888 27255 5940 27264
rect 5888 27221 5897 27255
rect 5897 27221 5931 27255
rect 5931 27221 5940 27255
rect 5888 27212 5940 27221
rect 19044 27212 19096 27264
rect 5796 26983 5848 26992
rect 5796 26949 5805 26983
rect 5805 26949 5839 26983
rect 5839 26949 5848 26983
rect 5796 26940 5848 26949
rect 11040 26940 11092 26992
rect 18768 26983 18820 26992
rect 18768 26949 18777 26983
rect 18777 26949 18811 26983
rect 18811 26949 18820 26983
rect 18768 26940 18820 26949
rect 6703 26881 6755 26890
rect 6767 26881 6819 26890
rect 6831 26881 6883 26890
rect 6703 26847 6725 26881
rect 6725 26847 6755 26881
rect 6767 26847 6817 26881
rect 6817 26847 6819 26881
rect 6831 26847 6851 26881
rect 6851 26847 6883 26881
rect 6703 26838 6755 26847
rect 6767 26838 6819 26847
rect 6831 26838 6883 26847
rect 6895 26881 6947 26890
rect 6895 26847 6909 26881
rect 6909 26847 6943 26881
rect 6943 26847 6947 26881
rect 6895 26838 6947 26847
rect 6959 26881 7011 26890
rect 10521 26881 10573 26890
rect 6959 26847 7001 26881
rect 7001 26847 7011 26881
rect 10521 26847 10531 26881
rect 10531 26847 10573 26881
rect 6959 26838 7011 26847
rect 10521 26838 10573 26847
rect 10585 26881 10637 26890
rect 10585 26847 10589 26881
rect 10589 26847 10623 26881
rect 10623 26847 10637 26881
rect 10585 26838 10637 26847
rect 10649 26881 10701 26890
rect 10713 26881 10765 26890
rect 10777 26881 10829 26890
rect 14339 26881 14391 26890
rect 14403 26881 14455 26890
rect 14467 26881 14519 26890
rect 10649 26847 10681 26881
rect 10681 26847 10701 26881
rect 10713 26847 10715 26881
rect 10715 26847 10765 26881
rect 10777 26847 10807 26881
rect 10807 26847 10829 26881
rect 14339 26847 14361 26881
rect 14361 26847 14391 26881
rect 14403 26847 14453 26881
rect 14453 26847 14455 26881
rect 14467 26847 14487 26881
rect 14487 26847 14519 26881
rect 10649 26838 10701 26847
rect 10713 26838 10765 26847
rect 10777 26838 10829 26847
rect 14339 26838 14391 26847
rect 14403 26838 14455 26847
rect 14467 26838 14519 26847
rect 14531 26881 14583 26890
rect 14531 26847 14545 26881
rect 14545 26847 14579 26881
rect 14579 26847 14583 26881
rect 14531 26838 14583 26847
rect 14595 26881 14647 26890
rect 18157 26881 18209 26890
rect 14595 26847 14637 26881
rect 14637 26847 14647 26881
rect 18157 26847 18167 26881
rect 18167 26847 18209 26881
rect 14595 26838 14647 26847
rect 18157 26838 18209 26847
rect 18221 26881 18273 26890
rect 18221 26847 18225 26881
rect 18225 26847 18259 26881
rect 18259 26847 18273 26881
rect 18221 26838 18273 26847
rect 18285 26881 18337 26890
rect 18349 26881 18401 26890
rect 18413 26881 18465 26890
rect 18285 26847 18317 26881
rect 18317 26847 18337 26881
rect 18349 26847 18351 26881
rect 18351 26847 18401 26881
rect 18413 26847 18443 26881
rect 18443 26847 18465 26881
rect 18285 26838 18337 26847
rect 18349 26838 18401 26847
rect 18413 26838 18465 26847
rect 6043 26337 6095 26346
rect 6107 26337 6159 26346
rect 6043 26303 6081 26337
rect 6081 26303 6095 26337
rect 6107 26303 6115 26337
rect 6115 26303 6159 26337
rect 6043 26294 6095 26303
rect 6107 26294 6159 26303
rect 6171 26337 6223 26346
rect 6171 26303 6173 26337
rect 6173 26303 6207 26337
rect 6207 26303 6223 26337
rect 6171 26294 6223 26303
rect 6235 26337 6287 26346
rect 6235 26303 6265 26337
rect 6265 26303 6287 26337
rect 6235 26294 6287 26303
rect 6299 26294 6351 26346
rect 9861 26337 9913 26346
rect 9861 26303 9887 26337
rect 9887 26303 9913 26337
rect 9861 26294 9913 26303
rect 9925 26337 9977 26346
rect 9989 26337 10041 26346
rect 10053 26337 10105 26346
rect 9925 26303 9945 26337
rect 9945 26303 9977 26337
rect 9989 26303 10037 26337
rect 10037 26303 10041 26337
rect 10053 26303 10071 26337
rect 10071 26303 10105 26337
rect 9925 26294 9977 26303
rect 9989 26294 10041 26303
rect 10053 26294 10105 26303
rect 10117 26337 10169 26346
rect 13679 26337 13731 26346
rect 13743 26337 13795 26346
rect 10117 26303 10129 26337
rect 10129 26303 10163 26337
rect 10163 26303 10169 26337
rect 13679 26303 13717 26337
rect 13717 26303 13731 26337
rect 13743 26303 13751 26337
rect 13751 26303 13795 26337
rect 10117 26294 10169 26303
rect 13679 26294 13731 26303
rect 13743 26294 13795 26303
rect 13807 26337 13859 26346
rect 13807 26303 13809 26337
rect 13809 26303 13843 26337
rect 13843 26303 13859 26337
rect 13807 26294 13859 26303
rect 13871 26337 13923 26346
rect 13871 26303 13901 26337
rect 13901 26303 13923 26337
rect 13871 26294 13923 26303
rect 13935 26294 13987 26346
rect 17497 26337 17549 26346
rect 17497 26303 17523 26337
rect 17523 26303 17549 26337
rect 17497 26294 17549 26303
rect 17561 26337 17613 26346
rect 17625 26337 17677 26346
rect 17689 26337 17741 26346
rect 17561 26303 17581 26337
rect 17581 26303 17613 26337
rect 17625 26303 17673 26337
rect 17673 26303 17677 26337
rect 17689 26303 17707 26337
rect 17707 26303 17741 26337
rect 17561 26294 17613 26303
rect 17625 26294 17677 26303
rect 17689 26294 17741 26303
rect 17753 26337 17805 26346
rect 17753 26303 17765 26337
rect 17765 26303 17799 26337
rect 17799 26303 17805 26337
rect 17753 26294 17805 26303
rect 6703 25793 6755 25802
rect 6767 25793 6819 25802
rect 6831 25793 6883 25802
rect 6703 25759 6725 25793
rect 6725 25759 6755 25793
rect 6767 25759 6817 25793
rect 6817 25759 6819 25793
rect 6831 25759 6851 25793
rect 6851 25759 6883 25793
rect 6703 25750 6755 25759
rect 6767 25750 6819 25759
rect 6831 25750 6883 25759
rect 6895 25793 6947 25802
rect 6895 25759 6909 25793
rect 6909 25759 6943 25793
rect 6943 25759 6947 25793
rect 6895 25750 6947 25759
rect 6959 25793 7011 25802
rect 10521 25793 10573 25802
rect 6959 25759 7001 25793
rect 7001 25759 7011 25793
rect 10521 25759 10531 25793
rect 10531 25759 10573 25793
rect 6959 25750 7011 25759
rect 10521 25750 10573 25759
rect 10585 25793 10637 25802
rect 10585 25759 10589 25793
rect 10589 25759 10623 25793
rect 10623 25759 10637 25793
rect 10585 25750 10637 25759
rect 10649 25793 10701 25802
rect 10713 25793 10765 25802
rect 10777 25793 10829 25802
rect 14339 25793 14391 25802
rect 14403 25793 14455 25802
rect 14467 25793 14519 25802
rect 10649 25759 10681 25793
rect 10681 25759 10701 25793
rect 10713 25759 10715 25793
rect 10715 25759 10765 25793
rect 10777 25759 10807 25793
rect 10807 25759 10829 25793
rect 14339 25759 14361 25793
rect 14361 25759 14391 25793
rect 14403 25759 14453 25793
rect 14453 25759 14455 25793
rect 14467 25759 14487 25793
rect 14487 25759 14519 25793
rect 10649 25750 10701 25759
rect 10713 25750 10765 25759
rect 10777 25750 10829 25759
rect 14339 25750 14391 25759
rect 14403 25750 14455 25759
rect 14467 25750 14519 25759
rect 14531 25793 14583 25802
rect 14531 25759 14545 25793
rect 14545 25759 14579 25793
rect 14579 25759 14583 25793
rect 14531 25750 14583 25759
rect 14595 25793 14647 25802
rect 18157 25793 18209 25802
rect 14595 25759 14637 25793
rect 14637 25759 14647 25793
rect 18157 25759 18167 25793
rect 18167 25759 18209 25793
rect 14595 25750 14647 25759
rect 18157 25750 18209 25759
rect 18221 25793 18273 25802
rect 18221 25759 18225 25793
rect 18225 25759 18259 25793
rect 18259 25759 18273 25793
rect 18221 25750 18273 25759
rect 18285 25793 18337 25802
rect 18349 25793 18401 25802
rect 18413 25793 18465 25802
rect 18285 25759 18317 25793
rect 18317 25759 18337 25793
rect 18349 25759 18351 25793
rect 18351 25759 18401 25793
rect 18413 25759 18443 25793
rect 18443 25759 18465 25793
rect 18285 25750 18337 25759
rect 18349 25750 18401 25759
rect 18413 25750 18465 25759
rect 14076 25308 14128 25360
rect 14720 25308 14772 25360
rect 6043 25249 6095 25258
rect 6107 25249 6159 25258
rect 6043 25215 6081 25249
rect 6081 25215 6095 25249
rect 6107 25215 6115 25249
rect 6115 25215 6159 25249
rect 6043 25206 6095 25215
rect 6107 25206 6159 25215
rect 6171 25249 6223 25258
rect 6171 25215 6173 25249
rect 6173 25215 6207 25249
rect 6207 25215 6223 25249
rect 6171 25206 6223 25215
rect 6235 25249 6287 25258
rect 6235 25215 6265 25249
rect 6265 25215 6287 25249
rect 6235 25206 6287 25215
rect 6299 25206 6351 25258
rect 9861 25249 9913 25258
rect 9861 25215 9887 25249
rect 9887 25215 9913 25249
rect 9861 25206 9913 25215
rect 9925 25249 9977 25258
rect 9989 25249 10041 25258
rect 10053 25249 10105 25258
rect 9925 25215 9945 25249
rect 9945 25215 9977 25249
rect 9989 25215 10037 25249
rect 10037 25215 10041 25249
rect 10053 25215 10071 25249
rect 10071 25215 10105 25249
rect 9925 25206 9977 25215
rect 9989 25206 10041 25215
rect 10053 25206 10105 25215
rect 10117 25249 10169 25258
rect 13679 25249 13731 25258
rect 13743 25249 13795 25258
rect 10117 25215 10129 25249
rect 10129 25215 10163 25249
rect 10163 25215 10169 25249
rect 13679 25215 13717 25249
rect 13717 25215 13731 25249
rect 13743 25215 13751 25249
rect 13751 25215 13795 25249
rect 10117 25206 10169 25215
rect 13679 25206 13731 25215
rect 13743 25206 13795 25215
rect 13807 25249 13859 25258
rect 13807 25215 13809 25249
rect 13809 25215 13843 25249
rect 13843 25215 13859 25249
rect 13807 25206 13859 25215
rect 13871 25249 13923 25258
rect 13871 25215 13901 25249
rect 13901 25215 13923 25249
rect 13871 25206 13923 25215
rect 13935 25206 13987 25258
rect 17497 25249 17549 25258
rect 17497 25215 17523 25249
rect 17523 25215 17549 25249
rect 17497 25206 17549 25215
rect 17561 25249 17613 25258
rect 17625 25249 17677 25258
rect 17689 25249 17741 25258
rect 17561 25215 17581 25249
rect 17581 25215 17613 25249
rect 17625 25215 17673 25249
rect 17673 25215 17677 25249
rect 17689 25215 17707 25249
rect 17707 25215 17741 25249
rect 17561 25206 17613 25215
rect 17625 25206 17677 25215
rect 17689 25206 17741 25215
rect 17753 25249 17805 25258
rect 17753 25215 17765 25249
rect 17765 25215 17799 25249
rect 17799 25215 17805 25249
rect 17753 25206 17805 25215
rect 6703 24705 6755 24714
rect 6767 24705 6819 24714
rect 6831 24705 6883 24714
rect 6703 24671 6725 24705
rect 6725 24671 6755 24705
rect 6767 24671 6817 24705
rect 6817 24671 6819 24705
rect 6831 24671 6851 24705
rect 6851 24671 6883 24705
rect 6703 24662 6755 24671
rect 6767 24662 6819 24671
rect 6831 24662 6883 24671
rect 6895 24705 6947 24714
rect 6895 24671 6909 24705
rect 6909 24671 6943 24705
rect 6943 24671 6947 24705
rect 6895 24662 6947 24671
rect 6959 24705 7011 24714
rect 10521 24705 10573 24714
rect 6959 24671 7001 24705
rect 7001 24671 7011 24705
rect 10521 24671 10531 24705
rect 10531 24671 10573 24705
rect 6959 24662 7011 24671
rect 10521 24662 10573 24671
rect 10585 24705 10637 24714
rect 10585 24671 10589 24705
rect 10589 24671 10623 24705
rect 10623 24671 10637 24705
rect 10585 24662 10637 24671
rect 10649 24705 10701 24714
rect 10713 24705 10765 24714
rect 10777 24705 10829 24714
rect 14339 24705 14391 24714
rect 14403 24705 14455 24714
rect 14467 24705 14519 24714
rect 10649 24671 10681 24705
rect 10681 24671 10701 24705
rect 10713 24671 10715 24705
rect 10715 24671 10765 24705
rect 10777 24671 10807 24705
rect 10807 24671 10829 24705
rect 14339 24671 14361 24705
rect 14361 24671 14391 24705
rect 14403 24671 14453 24705
rect 14453 24671 14455 24705
rect 14467 24671 14487 24705
rect 14487 24671 14519 24705
rect 10649 24662 10701 24671
rect 10713 24662 10765 24671
rect 10777 24662 10829 24671
rect 14339 24662 14391 24671
rect 14403 24662 14455 24671
rect 14467 24662 14519 24671
rect 14531 24705 14583 24714
rect 14531 24671 14545 24705
rect 14545 24671 14579 24705
rect 14579 24671 14583 24705
rect 14531 24662 14583 24671
rect 14595 24705 14647 24714
rect 18157 24705 18209 24714
rect 14595 24671 14637 24705
rect 14637 24671 14647 24705
rect 18157 24671 18167 24705
rect 18167 24671 18209 24705
rect 14595 24662 14647 24671
rect 18157 24662 18209 24671
rect 18221 24705 18273 24714
rect 18221 24671 18225 24705
rect 18225 24671 18259 24705
rect 18259 24671 18273 24705
rect 18221 24662 18273 24671
rect 18285 24705 18337 24714
rect 18349 24705 18401 24714
rect 18413 24705 18465 24714
rect 18285 24671 18317 24705
rect 18317 24671 18337 24705
rect 18349 24671 18351 24705
rect 18351 24671 18401 24705
rect 18413 24671 18443 24705
rect 18443 24671 18465 24705
rect 18285 24662 18337 24671
rect 18349 24662 18401 24671
rect 18413 24662 18465 24671
rect 6043 24161 6095 24170
rect 6107 24161 6159 24170
rect 6043 24127 6081 24161
rect 6081 24127 6095 24161
rect 6107 24127 6115 24161
rect 6115 24127 6159 24161
rect 6043 24118 6095 24127
rect 6107 24118 6159 24127
rect 6171 24161 6223 24170
rect 6171 24127 6173 24161
rect 6173 24127 6207 24161
rect 6207 24127 6223 24161
rect 6171 24118 6223 24127
rect 6235 24161 6287 24170
rect 6235 24127 6265 24161
rect 6265 24127 6287 24161
rect 6235 24118 6287 24127
rect 6299 24118 6351 24170
rect 9861 24161 9913 24170
rect 9861 24127 9887 24161
rect 9887 24127 9913 24161
rect 9861 24118 9913 24127
rect 9925 24161 9977 24170
rect 9989 24161 10041 24170
rect 10053 24161 10105 24170
rect 9925 24127 9945 24161
rect 9945 24127 9977 24161
rect 9989 24127 10037 24161
rect 10037 24127 10041 24161
rect 10053 24127 10071 24161
rect 10071 24127 10105 24161
rect 9925 24118 9977 24127
rect 9989 24118 10041 24127
rect 10053 24118 10105 24127
rect 10117 24161 10169 24170
rect 13679 24161 13731 24170
rect 13743 24161 13795 24170
rect 10117 24127 10129 24161
rect 10129 24127 10163 24161
rect 10163 24127 10169 24161
rect 13679 24127 13717 24161
rect 13717 24127 13731 24161
rect 13743 24127 13751 24161
rect 13751 24127 13795 24161
rect 10117 24118 10169 24127
rect 13679 24118 13731 24127
rect 13743 24118 13795 24127
rect 13807 24161 13859 24170
rect 13807 24127 13809 24161
rect 13809 24127 13843 24161
rect 13843 24127 13859 24161
rect 13807 24118 13859 24127
rect 13871 24161 13923 24170
rect 13871 24127 13901 24161
rect 13901 24127 13923 24161
rect 13871 24118 13923 24127
rect 13935 24118 13987 24170
rect 17497 24161 17549 24170
rect 17497 24127 17523 24161
rect 17523 24127 17549 24161
rect 17497 24118 17549 24127
rect 17561 24161 17613 24170
rect 17625 24161 17677 24170
rect 17689 24161 17741 24170
rect 17561 24127 17581 24161
rect 17581 24127 17613 24161
rect 17625 24127 17673 24161
rect 17673 24127 17677 24161
rect 17689 24127 17707 24161
rect 17707 24127 17741 24161
rect 17561 24118 17613 24127
rect 17625 24118 17677 24127
rect 17689 24118 17741 24127
rect 17753 24161 17805 24170
rect 17753 24127 17765 24161
rect 17765 24127 17799 24161
rect 17799 24127 17805 24161
rect 17753 24118 17805 24127
rect 6703 23617 6755 23626
rect 6767 23617 6819 23626
rect 6831 23617 6883 23626
rect 6703 23583 6725 23617
rect 6725 23583 6755 23617
rect 6767 23583 6817 23617
rect 6817 23583 6819 23617
rect 6831 23583 6851 23617
rect 6851 23583 6883 23617
rect 6703 23574 6755 23583
rect 6767 23574 6819 23583
rect 6831 23574 6883 23583
rect 6895 23617 6947 23626
rect 6895 23583 6909 23617
rect 6909 23583 6943 23617
rect 6943 23583 6947 23617
rect 6895 23574 6947 23583
rect 6959 23617 7011 23626
rect 10521 23617 10573 23626
rect 6959 23583 7001 23617
rect 7001 23583 7011 23617
rect 10521 23583 10531 23617
rect 10531 23583 10573 23617
rect 6959 23574 7011 23583
rect 10521 23574 10573 23583
rect 10585 23617 10637 23626
rect 10585 23583 10589 23617
rect 10589 23583 10623 23617
rect 10623 23583 10637 23617
rect 10585 23574 10637 23583
rect 10649 23617 10701 23626
rect 10713 23617 10765 23626
rect 10777 23617 10829 23626
rect 14339 23617 14391 23626
rect 14403 23617 14455 23626
rect 14467 23617 14519 23626
rect 10649 23583 10681 23617
rect 10681 23583 10701 23617
rect 10713 23583 10715 23617
rect 10715 23583 10765 23617
rect 10777 23583 10807 23617
rect 10807 23583 10829 23617
rect 14339 23583 14361 23617
rect 14361 23583 14391 23617
rect 14403 23583 14453 23617
rect 14453 23583 14455 23617
rect 14467 23583 14487 23617
rect 14487 23583 14519 23617
rect 10649 23574 10701 23583
rect 10713 23574 10765 23583
rect 10777 23574 10829 23583
rect 14339 23574 14391 23583
rect 14403 23574 14455 23583
rect 14467 23574 14519 23583
rect 14531 23617 14583 23626
rect 14531 23583 14545 23617
rect 14545 23583 14579 23617
rect 14579 23583 14583 23617
rect 14531 23574 14583 23583
rect 14595 23617 14647 23626
rect 18157 23617 18209 23626
rect 14595 23583 14637 23617
rect 14637 23583 14647 23617
rect 18157 23583 18167 23617
rect 18167 23583 18209 23617
rect 14595 23574 14647 23583
rect 18157 23574 18209 23583
rect 18221 23617 18273 23626
rect 18221 23583 18225 23617
rect 18225 23583 18259 23617
rect 18259 23583 18273 23617
rect 18221 23574 18273 23583
rect 18285 23617 18337 23626
rect 18349 23617 18401 23626
rect 18413 23617 18465 23626
rect 18285 23583 18317 23617
rect 18317 23583 18337 23617
rect 18349 23583 18351 23617
rect 18351 23583 18401 23617
rect 18413 23583 18443 23617
rect 18443 23583 18465 23617
rect 18285 23574 18337 23583
rect 18349 23574 18401 23583
rect 18413 23574 18465 23583
rect 6043 23073 6095 23082
rect 6107 23073 6159 23082
rect 6043 23039 6081 23073
rect 6081 23039 6095 23073
rect 6107 23039 6115 23073
rect 6115 23039 6159 23073
rect 6043 23030 6095 23039
rect 6107 23030 6159 23039
rect 6171 23073 6223 23082
rect 6171 23039 6173 23073
rect 6173 23039 6207 23073
rect 6207 23039 6223 23073
rect 6171 23030 6223 23039
rect 6235 23073 6287 23082
rect 6235 23039 6265 23073
rect 6265 23039 6287 23073
rect 6235 23030 6287 23039
rect 6299 23030 6351 23082
rect 9861 23073 9913 23082
rect 9861 23039 9887 23073
rect 9887 23039 9913 23073
rect 9861 23030 9913 23039
rect 9925 23073 9977 23082
rect 9989 23073 10041 23082
rect 10053 23073 10105 23082
rect 9925 23039 9945 23073
rect 9945 23039 9977 23073
rect 9989 23039 10037 23073
rect 10037 23039 10041 23073
rect 10053 23039 10071 23073
rect 10071 23039 10105 23073
rect 9925 23030 9977 23039
rect 9989 23030 10041 23039
rect 10053 23030 10105 23039
rect 10117 23073 10169 23082
rect 13679 23073 13731 23082
rect 13743 23073 13795 23082
rect 10117 23039 10129 23073
rect 10129 23039 10163 23073
rect 10163 23039 10169 23073
rect 13679 23039 13717 23073
rect 13717 23039 13731 23073
rect 13743 23039 13751 23073
rect 13751 23039 13795 23073
rect 10117 23030 10169 23039
rect 13679 23030 13731 23039
rect 13743 23030 13795 23039
rect 13807 23073 13859 23082
rect 13807 23039 13809 23073
rect 13809 23039 13843 23073
rect 13843 23039 13859 23073
rect 13807 23030 13859 23039
rect 13871 23073 13923 23082
rect 13871 23039 13901 23073
rect 13901 23039 13923 23073
rect 13871 23030 13923 23039
rect 13935 23030 13987 23082
rect 17497 23073 17549 23082
rect 17497 23039 17523 23073
rect 17523 23039 17549 23073
rect 17497 23030 17549 23039
rect 17561 23073 17613 23082
rect 17625 23073 17677 23082
rect 17689 23073 17741 23082
rect 17561 23039 17581 23073
rect 17581 23039 17613 23073
rect 17625 23039 17673 23073
rect 17673 23039 17677 23073
rect 17689 23039 17707 23073
rect 17707 23039 17741 23073
rect 17561 23030 17613 23039
rect 17625 23030 17677 23039
rect 17689 23030 17741 23039
rect 17753 23073 17805 23082
rect 17753 23039 17765 23073
rect 17765 23039 17799 23073
rect 17799 23039 17805 23073
rect 17753 23030 17805 23039
rect 6703 22529 6755 22538
rect 6767 22529 6819 22538
rect 6831 22529 6883 22538
rect 6703 22495 6725 22529
rect 6725 22495 6755 22529
rect 6767 22495 6817 22529
rect 6817 22495 6819 22529
rect 6831 22495 6851 22529
rect 6851 22495 6883 22529
rect 6703 22486 6755 22495
rect 6767 22486 6819 22495
rect 6831 22486 6883 22495
rect 6895 22529 6947 22538
rect 6895 22495 6909 22529
rect 6909 22495 6943 22529
rect 6943 22495 6947 22529
rect 6895 22486 6947 22495
rect 6959 22529 7011 22538
rect 10521 22529 10573 22538
rect 6959 22495 7001 22529
rect 7001 22495 7011 22529
rect 10521 22495 10531 22529
rect 10531 22495 10573 22529
rect 6959 22486 7011 22495
rect 10521 22486 10573 22495
rect 10585 22529 10637 22538
rect 10585 22495 10589 22529
rect 10589 22495 10623 22529
rect 10623 22495 10637 22529
rect 10585 22486 10637 22495
rect 10649 22529 10701 22538
rect 10713 22529 10765 22538
rect 10777 22529 10829 22538
rect 14339 22529 14391 22538
rect 14403 22529 14455 22538
rect 14467 22529 14519 22538
rect 10649 22495 10681 22529
rect 10681 22495 10701 22529
rect 10713 22495 10715 22529
rect 10715 22495 10765 22529
rect 10777 22495 10807 22529
rect 10807 22495 10829 22529
rect 14339 22495 14361 22529
rect 14361 22495 14391 22529
rect 14403 22495 14453 22529
rect 14453 22495 14455 22529
rect 14467 22495 14487 22529
rect 14487 22495 14519 22529
rect 10649 22486 10701 22495
rect 10713 22486 10765 22495
rect 10777 22486 10829 22495
rect 14339 22486 14391 22495
rect 14403 22486 14455 22495
rect 14467 22486 14519 22495
rect 14531 22529 14583 22538
rect 14531 22495 14545 22529
rect 14545 22495 14579 22529
rect 14579 22495 14583 22529
rect 14531 22486 14583 22495
rect 14595 22529 14647 22538
rect 18157 22529 18209 22538
rect 14595 22495 14637 22529
rect 14637 22495 14647 22529
rect 18157 22495 18167 22529
rect 18167 22495 18209 22529
rect 14595 22486 14647 22495
rect 18157 22486 18209 22495
rect 18221 22529 18273 22538
rect 18221 22495 18225 22529
rect 18225 22495 18259 22529
rect 18259 22495 18273 22529
rect 18221 22486 18273 22495
rect 18285 22529 18337 22538
rect 18349 22529 18401 22538
rect 18413 22529 18465 22538
rect 18285 22495 18317 22529
rect 18317 22495 18337 22529
rect 18349 22495 18351 22529
rect 18351 22495 18401 22529
rect 18413 22495 18443 22529
rect 18443 22495 18465 22529
rect 18285 22486 18337 22495
rect 18349 22486 18401 22495
rect 18413 22486 18465 22495
rect 6043 21985 6095 21994
rect 6107 21985 6159 21994
rect 6043 21951 6081 21985
rect 6081 21951 6095 21985
rect 6107 21951 6115 21985
rect 6115 21951 6159 21985
rect 6043 21942 6095 21951
rect 6107 21942 6159 21951
rect 6171 21985 6223 21994
rect 6171 21951 6173 21985
rect 6173 21951 6207 21985
rect 6207 21951 6223 21985
rect 6171 21942 6223 21951
rect 6235 21985 6287 21994
rect 6235 21951 6265 21985
rect 6265 21951 6287 21985
rect 6235 21942 6287 21951
rect 6299 21942 6351 21994
rect 9861 21985 9913 21994
rect 9861 21951 9887 21985
rect 9887 21951 9913 21985
rect 9861 21942 9913 21951
rect 9925 21985 9977 21994
rect 9989 21985 10041 21994
rect 10053 21985 10105 21994
rect 9925 21951 9945 21985
rect 9945 21951 9977 21985
rect 9989 21951 10037 21985
rect 10037 21951 10041 21985
rect 10053 21951 10071 21985
rect 10071 21951 10105 21985
rect 9925 21942 9977 21951
rect 9989 21942 10041 21951
rect 10053 21942 10105 21951
rect 10117 21985 10169 21994
rect 13679 21985 13731 21994
rect 13743 21985 13795 21994
rect 10117 21951 10129 21985
rect 10129 21951 10163 21985
rect 10163 21951 10169 21985
rect 13679 21951 13717 21985
rect 13717 21951 13731 21985
rect 13743 21951 13751 21985
rect 13751 21951 13795 21985
rect 10117 21942 10169 21951
rect 13679 21942 13731 21951
rect 13743 21942 13795 21951
rect 13807 21985 13859 21994
rect 13807 21951 13809 21985
rect 13809 21951 13843 21985
rect 13843 21951 13859 21985
rect 13807 21942 13859 21951
rect 13871 21985 13923 21994
rect 13871 21951 13901 21985
rect 13901 21951 13923 21985
rect 13871 21942 13923 21951
rect 13935 21942 13987 21994
rect 17497 21985 17549 21994
rect 17497 21951 17523 21985
rect 17523 21951 17549 21985
rect 17497 21942 17549 21951
rect 17561 21985 17613 21994
rect 17625 21985 17677 21994
rect 17689 21985 17741 21994
rect 17561 21951 17581 21985
rect 17581 21951 17613 21985
rect 17625 21951 17673 21985
rect 17673 21951 17677 21985
rect 17689 21951 17707 21985
rect 17707 21951 17741 21985
rect 17561 21942 17613 21951
rect 17625 21942 17677 21951
rect 17689 21942 17741 21951
rect 17753 21985 17805 21994
rect 17753 21951 17765 21985
rect 17765 21951 17799 21985
rect 17799 21951 17805 21985
rect 17753 21942 17805 21951
rect 6703 21441 6755 21450
rect 6767 21441 6819 21450
rect 6831 21441 6883 21450
rect 6703 21407 6725 21441
rect 6725 21407 6755 21441
rect 6767 21407 6817 21441
rect 6817 21407 6819 21441
rect 6831 21407 6851 21441
rect 6851 21407 6883 21441
rect 6703 21398 6755 21407
rect 6767 21398 6819 21407
rect 6831 21398 6883 21407
rect 6895 21441 6947 21450
rect 6895 21407 6909 21441
rect 6909 21407 6943 21441
rect 6943 21407 6947 21441
rect 6895 21398 6947 21407
rect 6959 21441 7011 21450
rect 10521 21441 10573 21450
rect 6959 21407 7001 21441
rect 7001 21407 7011 21441
rect 10521 21407 10531 21441
rect 10531 21407 10573 21441
rect 6959 21398 7011 21407
rect 10521 21398 10573 21407
rect 10585 21441 10637 21450
rect 10585 21407 10589 21441
rect 10589 21407 10623 21441
rect 10623 21407 10637 21441
rect 10585 21398 10637 21407
rect 10649 21441 10701 21450
rect 10713 21441 10765 21450
rect 10777 21441 10829 21450
rect 14339 21441 14391 21450
rect 14403 21441 14455 21450
rect 14467 21441 14519 21450
rect 10649 21407 10681 21441
rect 10681 21407 10701 21441
rect 10713 21407 10715 21441
rect 10715 21407 10765 21441
rect 10777 21407 10807 21441
rect 10807 21407 10829 21441
rect 14339 21407 14361 21441
rect 14361 21407 14391 21441
rect 14403 21407 14453 21441
rect 14453 21407 14455 21441
rect 14467 21407 14487 21441
rect 14487 21407 14519 21441
rect 10649 21398 10701 21407
rect 10713 21398 10765 21407
rect 10777 21398 10829 21407
rect 14339 21398 14391 21407
rect 14403 21398 14455 21407
rect 14467 21398 14519 21407
rect 14531 21441 14583 21450
rect 14531 21407 14545 21441
rect 14545 21407 14579 21441
rect 14579 21407 14583 21441
rect 14531 21398 14583 21407
rect 14595 21441 14647 21450
rect 18157 21441 18209 21450
rect 14595 21407 14637 21441
rect 14637 21407 14647 21441
rect 18157 21407 18167 21441
rect 18167 21407 18209 21441
rect 14595 21398 14647 21407
rect 18157 21398 18209 21407
rect 18221 21441 18273 21450
rect 18221 21407 18225 21441
rect 18225 21407 18259 21441
rect 18259 21407 18273 21441
rect 18221 21398 18273 21407
rect 18285 21441 18337 21450
rect 18349 21441 18401 21450
rect 18413 21441 18465 21450
rect 18285 21407 18317 21441
rect 18317 21407 18337 21441
rect 18349 21407 18351 21441
rect 18351 21407 18401 21441
rect 18413 21407 18443 21441
rect 18443 21407 18465 21441
rect 18285 21398 18337 21407
rect 18349 21398 18401 21407
rect 18413 21398 18465 21407
rect 6043 20897 6095 20906
rect 6107 20897 6159 20906
rect 6043 20863 6081 20897
rect 6081 20863 6095 20897
rect 6107 20863 6115 20897
rect 6115 20863 6159 20897
rect 6043 20854 6095 20863
rect 6107 20854 6159 20863
rect 6171 20897 6223 20906
rect 6171 20863 6173 20897
rect 6173 20863 6207 20897
rect 6207 20863 6223 20897
rect 6171 20854 6223 20863
rect 6235 20897 6287 20906
rect 6235 20863 6265 20897
rect 6265 20863 6287 20897
rect 6235 20854 6287 20863
rect 6299 20854 6351 20906
rect 9861 20897 9913 20906
rect 9861 20863 9887 20897
rect 9887 20863 9913 20897
rect 9861 20854 9913 20863
rect 9925 20897 9977 20906
rect 9989 20897 10041 20906
rect 10053 20897 10105 20906
rect 9925 20863 9945 20897
rect 9945 20863 9977 20897
rect 9989 20863 10037 20897
rect 10037 20863 10041 20897
rect 10053 20863 10071 20897
rect 10071 20863 10105 20897
rect 9925 20854 9977 20863
rect 9989 20854 10041 20863
rect 10053 20854 10105 20863
rect 10117 20897 10169 20906
rect 13679 20897 13731 20906
rect 13743 20897 13795 20906
rect 10117 20863 10129 20897
rect 10129 20863 10163 20897
rect 10163 20863 10169 20897
rect 13679 20863 13717 20897
rect 13717 20863 13731 20897
rect 13743 20863 13751 20897
rect 13751 20863 13795 20897
rect 10117 20854 10169 20863
rect 13679 20854 13731 20863
rect 13743 20854 13795 20863
rect 13807 20897 13859 20906
rect 13807 20863 13809 20897
rect 13809 20863 13843 20897
rect 13843 20863 13859 20897
rect 13807 20854 13859 20863
rect 13871 20897 13923 20906
rect 13871 20863 13901 20897
rect 13901 20863 13923 20897
rect 13871 20854 13923 20863
rect 13935 20854 13987 20906
rect 17497 20897 17549 20906
rect 17497 20863 17523 20897
rect 17523 20863 17549 20897
rect 17497 20854 17549 20863
rect 17561 20897 17613 20906
rect 17625 20897 17677 20906
rect 17689 20897 17741 20906
rect 17561 20863 17581 20897
rect 17581 20863 17613 20897
rect 17625 20863 17673 20897
rect 17673 20863 17677 20897
rect 17689 20863 17707 20897
rect 17707 20863 17741 20897
rect 17561 20854 17613 20863
rect 17625 20854 17677 20863
rect 17689 20854 17741 20863
rect 17753 20897 17805 20906
rect 17753 20863 17765 20897
rect 17765 20863 17799 20897
rect 17799 20863 17805 20897
rect 17753 20854 17805 20863
rect 6703 20353 6755 20362
rect 6767 20353 6819 20362
rect 6831 20353 6883 20362
rect 6703 20319 6725 20353
rect 6725 20319 6755 20353
rect 6767 20319 6817 20353
rect 6817 20319 6819 20353
rect 6831 20319 6851 20353
rect 6851 20319 6883 20353
rect 6703 20310 6755 20319
rect 6767 20310 6819 20319
rect 6831 20310 6883 20319
rect 6895 20353 6947 20362
rect 6895 20319 6909 20353
rect 6909 20319 6943 20353
rect 6943 20319 6947 20353
rect 6895 20310 6947 20319
rect 6959 20353 7011 20362
rect 10521 20353 10573 20362
rect 6959 20319 7001 20353
rect 7001 20319 7011 20353
rect 10521 20319 10531 20353
rect 10531 20319 10573 20353
rect 6959 20310 7011 20319
rect 10521 20310 10573 20319
rect 10585 20353 10637 20362
rect 10585 20319 10589 20353
rect 10589 20319 10623 20353
rect 10623 20319 10637 20353
rect 10585 20310 10637 20319
rect 10649 20353 10701 20362
rect 10713 20353 10765 20362
rect 10777 20353 10829 20362
rect 14339 20353 14391 20362
rect 14403 20353 14455 20362
rect 14467 20353 14519 20362
rect 10649 20319 10681 20353
rect 10681 20319 10701 20353
rect 10713 20319 10715 20353
rect 10715 20319 10765 20353
rect 10777 20319 10807 20353
rect 10807 20319 10829 20353
rect 14339 20319 14361 20353
rect 14361 20319 14391 20353
rect 14403 20319 14453 20353
rect 14453 20319 14455 20353
rect 14467 20319 14487 20353
rect 14487 20319 14519 20353
rect 10649 20310 10701 20319
rect 10713 20310 10765 20319
rect 10777 20310 10829 20319
rect 14339 20310 14391 20319
rect 14403 20310 14455 20319
rect 14467 20310 14519 20319
rect 14531 20353 14583 20362
rect 14531 20319 14545 20353
rect 14545 20319 14579 20353
rect 14579 20319 14583 20353
rect 14531 20310 14583 20319
rect 14595 20353 14647 20362
rect 18157 20353 18209 20362
rect 14595 20319 14637 20353
rect 14637 20319 14647 20353
rect 18157 20319 18167 20353
rect 18167 20319 18209 20353
rect 14595 20310 14647 20319
rect 18157 20310 18209 20319
rect 18221 20353 18273 20362
rect 18221 20319 18225 20353
rect 18225 20319 18259 20353
rect 18259 20319 18273 20353
rect 18221 20310 18273 20319
rect 18285 20353 18337 20362
rect 18349 20353 18401 20362
rect 18413 20353 18465 20362
rect 18285 20319 18317 20353
rect 18317 20319 18337 20353
rect 18349 20319 18351 20353
rect 18351 20319 18401 20353
rect 18413 20319 18443 20353
rect 18443 20319 18465 20353
rect 18285 20310 18337 20319
rect 18349 20310 18401 20319
rect 18413 20310 18465 20319
rect 6043 19809 6095 19818
rect 6107 19809 6159 19818
rect 6043 19775 6081 19809
rect 6081 19775 6095 19809
rect 6107 19775 6115 19809
rect 6115 19775 6159 19809
rect 6043 19766 6095 19775
rect 6107 19766 6159 19775
rect 6171 19809 6223 19818
rect 6171 19775 6173 19809
rect 6173 19775 6207 19809
rect 6207 19775 6223 19809
rect 6171 19766 6223 19775
rect 6235 19809 6287 19818
rect 6235 19775 6265 19809
rect 6265 19775 6287 19809
rect 6235 19766 6287 19775
rect 6299 19766 6351 19818
rect 9861 19809 9913 19818
rect 9861 19775 9887 19809
rect 9887 19775 9913 19809
rect 9861 19766 9913 19775
rect 9925 19809 9977 19818
rect 9989 19809 10041 19818
rect 10053 19809 10105 19818
rect 9925 19775 9945 19809
rect 9945 19775 9977 19809
rect 9989 19775 10037 19809
rect 10037 19775 10041 19809
rect 10053 19775 10071 19809
rect 10071 19775 10105 19809
rect 9925 19766 9977 19775
rect 9989 19766 10041 19775
rect 10053 19766 10105 19775
rect 10117 19809 10169 19818
rect 13679 19809 13731 19818
rect 13743 19809 13795 19818
rect 10117 19775 10129 19809
rect 10129 19775 10163 19809
rect 10163 19775 10169 19809
rect 13679 19775 13717 19809
rect 13717 19775 13731 19809
rect 13743 19775 13751 19809
rect 13751 19775 13795 19809
rect 10117 19766 10169 19775
rect 13679 19766 13731 19775
rect 13743 19766 13795 19775
rect 13807 19809 13859 19818
rect 13807 19775 13809 19809
rect 13809 19775 13843 19809
rect 13843 19775 13859 19809
rect 13807 19766 13859 19775
rect 13871 19809 13923 19818
rect 13871 19775 13901 19809
rect 13901 19775 13923 19809
rect 13871 19766 13923 19775
rect 13935 19766 13987 19818
rect 17497 19809 17549 19818
rect 17497 19775 17523 19809
rect 17523 19775 17549 19809
rect 17497 19766 17549 19775
rect 17561 19809 17613 19818
rect 17625 19809 17677 19818
rect 17689 19809 17741 19818
rect 17561 19775 17581 19809
rect 17581 19775 17613 19809
rect 17625 19775 17673 19809
rect 17673 19775 17677 19809
rect 17689 19775 17707 19809
rect 17707 19775 17741 19809
rect 17561 19766 17613 19775
rect 17625 19766 17677 19775
rect 17689 19766 17741 19775
rect 17753 19809 17805 19818
rect 17753 19775 17765 19809
rect 17765 19775 17799 19809
rect 17799 19775 17805 19809
rect 17753 19766 17805 19775
rect 6703 19265 6755 19274
rect 6767 19265 6819 19274
rect 6831 19265 6883 19274
rect 6703 19231 6725 19265
rect 6725 19231 6755 19265
rect 6767 19231 6817 19265
rect 6817 19231 6819 19265
rect 6831 19231 6851 19265
rect 6851 19231 6883 19265
rect 6703 19222 6755 19231
rect 6767 19222 6819 19231
rect 6831 19222 6883 19231
rect 6895 19265 6947 19274
rect 6895 19231 6909 19265
rect 6909 19231 6943 19265
rect 6943 19231 6947 19265
rect 6895 19222 6947 19231
rect 6959 19265 7011 19274
rect 10521 19265 10573 19274
rect 6959 19231 7001 19265
rect 7001 19231 7011 19265
rect 10521 19231 10531 19265
rect 10531 19231 10573 19265
rect 6959 19222 7011 19231
rect 10521 19222 10573 19231
rect 10585 19265 10637 19274
rect 10585 19231 10589 19265
rect 10589 19231 10623 19265
rect 10623 19231 10637 19265
rect 10585 19222 10637 19231
rect 10649 19265 10701 19274
rect 10713 19265 10765 19274
rect 10777 19265 10829 19274
rect 14339 19265 14391 19274
rect 14403 19265 14455 19274
rect 14467 19265 14519 19274
rect 10649 19231 10681 19265
rect 10681 19231 10701 19265
rect 10713 19231 10715 19265
rect 10715 19231 10765 19265
rect 10777 19231 10807 19265
rect 10807 19231 10829 19265
rect 14339 19231 14361 19265
rect 14361 19231 14391 19265
rect 14403 19231 14453 19265
rect 14453 19231 14455 19265
rect 14467 19231 14487 19265
rect 14487 19231 14519 19265
rect 10649 19222 10701 19231
rect 10713 19222 10765 19231
rect 10777 19222 10829 19231
rect 14339 19222 14391 19231
rect 14403 19222 14455 19231
rect 14467 19222 14519 19231
rect 14531 19265 14583 19274
rect 14531 19231 14545 19265
rect 14545 19231 14579 19265
rect 14579 19231 14583 19265
rect 14531 19222 14583 19231
rect 14595 19265 14647 19274
rect 18157 19265 18209 19274
rect 14595 19231 14637 19265
rect 14637 19231 14647 19265
rect 18157 19231 18167 19265
rect 18167 19231 18209 19265
rect 14595 19222 14647 19231
rect 18157 19222 18209 19231
rect 18221 19265 18273 19274
rect 18221 19231 18225 19265
rect 18225 19231 18259 19265
rect 18259 19231 18273 19265
rect 18221 19222 18273 19231
rect 18285 19265 18337 19274
rect 18349 19265 18401 19274
rect 18413 19265 18465 19274
rect 18285 19231 18317 19265
rect 18317 19231 18337 19265
rect 18349 19231 18351 19265
rect 18351 19231 18401 19265
rect 18413 19231 18443 19265
rect 18443 19231 18465 19265
rect 18285 19222 18337 19231
rect 18349 19222 18401 19231
rect 18413 19222 18465 19231
rect 6043 18721 6095 18730
rect 6107 18721 6159 18730
rect 6043 18687 6081 18721
rect 6081 18687 6095 18721
rect 6107 18687 6115 18721
rect 6115 18687 6159 18721
rect 6043 18678 6095 18687
rect 6107 18678 6159 18687
rect 6171 18721 6223 18730
rect 6171 18687 6173 18721
rect 6173 18687 6207 18721
rect 6207 18687 6223 18721
rect 6171 18678 6223 18687
rect 6235 18721 6287 18730
rect 6235 18687 6265 18721
rect 6265 18687 6287 18721
rect 6235 18678 6287 18687
rect 6299 18678 6351 18730
rect 9861 18721 9913 18730
rect 9861 18687 9887 18721
rect 9887 18687 9913 18721
rect 9861 18678 9913 18687
rect 9925 18721 9977 18730
rect 9989 18721 10041 18730
rect 10053 18721 10105 18730
rect 9925 18687 9945 18721
rect 9945 18687 9977 18721
rect 9989 18687 10037 18721
rect 10037 18687 10041 18721
rect 10053 18687 10071 18721
rect 10071 18687 10105 18721
rect 9925 18678 9977 18687
rect 9989 18678 10041 18687
rect 10053 18678 10105 18687
rect 10117 18721 10169 18730
rect 13679 18721 13731 18730
rect 13743 18721 13795 18730
rect 10117 18687 10129 18721
rect 10129 18687 10163 18721
rect 10163 18687 10169 18721
rect 13679 18687 13717 18721
rect 13717 18687 13731 18721
rect 13743 18687 13751 18721
rect 13751 18687 13795 18721
rect 10117 18678 10169 18687
rect 13679 18678 13731 18687
rect 13743 18678 13795 18687
rect 13807 18721 13859 18730
rect 13807 18687 13809 18721
rect 13809 18687 13843 18721
rect 13843 18687 13859 18721
rect 13807 18678 13859 18687
rect 13871 18721 13923 18730
rect 13871 18687 13901 18721
rect 13901 18687 13923 18721
rect 13871 18678 13923 18687
rect 13935 18678 13987 18730
rect 17497 18721 17549 18730
rect 17497 18687 17523 18721
rect 17523 18687 17549 18721
rect 17497 18678 17549 18687
rect 17561 18721 17613 18730
rect 17625 18721 17677 18730
rect 17689 18721 17741 18730
rect 17561 18687 17581 18721
rect 17581 18687 17613 18721
rect 17625 18687 17673 18721
rect 17673 18687 17677 18721
rect 17689 18687 17707 18721
rect 17707 18687 17741 18721
rect 17561 18678 17613 18687
rect 17625 18678 17677 18687
rect 17689 18678 17741 18687
rect 17753 18721 17805 18730
rect 17753 18687 17765 18721
rect 17765 18687 17799 18721
rect 17799 18687 17805 18721
rect 17753 18678 17805 18687
rect 6703 18177 6755 18186
rect 6767 18177 6819 18186
rect 6831 18177 6883 18186
rect 6703 18143 6725 18177
rect 6725 18143 6755 18177
rect 6767 18143 6817 18177
rect 6817 18143 6819 18177
rect 6831 18143 6851 18177
rect 6851 18143 6883 18177
rect 6703 18134 6755 18143
rect 6767 18134 6819 18143
rect 6831 18134 6883 18143
rect 6895 18177 6947 18186
rect 6895 18143 6909 18177
rect 6909 18143 6943 18177
rect 6943 18143 6947 18177
rect 6895 18134 6947 18143
rect 6959 18177 7011 18186
rect 10521 18177 10573 18186
rect 6959 18143 7001 18177
rect 7001 18143 7011 18177
rect 10521 18143 10531 18177
rect 10531 18143 10573 18177
rect 6959 18134 7011 18143
rect 10521 18134 10573 18143
rect 10585 18177 10637 18186
rect 10585 18143 10589 18177
rect 10589 18143 10623 18177
rect 10623 18143 10637 18177
rect 10585 18134 10637 18143
rect 10649 18177 10701 18186
rect 10713 18177 10765 18186
rect 10777 18177 10829 18186
rect 14339 18177 14391 18186
rect 14403 18177 14455 18186
rect 14467 18177 14519 18186
rect 10649 18143 10681 18177
rect 10681 18143 10701 18177
rect 10713 18143 10715 18177
rect 10715 18143 10765 18177
rect 10777 18143 10807 18177
rect 10807 18143 10829 18177
rect 14339 18143 14361 18177
rect 14361 18143 14391 18177
rect 14403 18143 14453 18177
rect 14453 18143 14455 18177
rect 14467 18143 14487 18177
rect 14487 18143 14519 18177
rect 10649 18134 10701 18143
rect 10713 18134 10765 18143
rect 10777 18134 10829 18143
rect 14339 18134 14391 18143
rect 14403 18134 14455 18143
rect 14467 18134 14519 18143
rect 14531 18177 14583 18186
rect 14531 18143 14545 18177
rect 14545 18143 14579 18177
rect 14579 18143 14583 18177
rect 14531 18134 14583 18143
rect 14595 18177 14647 18186
rect 18157 18177 18209 18186
rect 14595 18143 14637 18177
rect 14637 18143 14647 18177
rect 18157 18143 18167 18177
rect 18167 18143 18209 18177
rect 14595 18134 14647 18143
rect 18157 18134 18209 18143
rect 18221 18177 18273 18186
rect 18221 18143 18225 18177
rect 18225 18143 18259 18177
rect 18259 18143 18273 18177
rect 18221 18134 18273 18143
rect 18285 18177 18337 18186
rect 18349 18177 18401 18186
rect 18413 18177 18465 18186
rect 18285 18143 18317 18177
rect 18317 18143 18337 18177
rect 18349 18143 18351 18177
rect 18351 18143 18401 18177
rect 18413 18143 18443 18177
rect 18443 18143 18465 18177
rect 18285 18134 18337 18143
rect 18349 18134 18401 18143
rect 18413 18134 18465 18143
rect 6043 17633 6095 17642
rect 6107 17633 6159 17642
rect 6043 17599 6081 17633
rect 6081 17599 6095 17633
rect 6107 17599 6115 17633
rect 6115 17599 6159 17633
rect 6043 17590 6095 17599
rect 6107 17590 6159 17599
rect 6171 17633 6223 17642
rect 6171 17599 6173 17633
rect 6173 17599 6207 17633
rect 6207 17599 6223 17633
rect 6171 17590 6223 17599
rect 6235 17633 6287 17642
rect 6235 17599 6265 17633
rect 6265 17599 6287 17633
rect 6235 17590 6287 17599
rect 6299 17590 6351 17642
rect 9861 17633 9913 17642
rect 9861 17599 9887 17633
rect 9887 17599 9913 17633
rect 9861 17590 9913 17599
rect 9925 17633 9977 17642
rect 9989 17633 10041 17642
rect 10053 17633 10105 17642
rect 9925 17599 9945 17633
rect 9945 17599 9977 17633
rect 9989 17599 10037 17633
rect 10037 17599 10041 17633
rect 10053 17599 10071 17633
rect 10071 17599 10105 17633
rect 9925 17590 9977 17599
rect 9989 17590 10041 17599
rect 10053 17590 10105 17599
rect 10117 17633 10169 17642
rect 13679 17633 13731 17642
rect 13743 17633 13795 17642
rect 10117 17599 10129 17633
rect 10129 17599 10163 17633
rect 10163 17599 10169 17633
rect 13679 17599 13717 17633
rect 13717 17599 13731 17633
rect 13743 17599 13751 17633
rect 13751 17599 13795 17633
rect 10117 17590 10169 17599
rect 13679 17590 13731 17599
rect 13743 17590 13795 17599
rect 13807 17633 13859 17642
rect 13807 17599 13809 17633
rect 13809 17599 13843 17633
rect 13843 17599 13859 17633
rect 13807 17590 13859 17599
rect 13871 17633 13923 17642
rect 13871 17599 13901 17633
rect 13901 17599 13923 17633
rect 13871 17590 13923 17599
rect 13935 17590 13987 17642
rect 17497 17633 17549 17642
rect 17497 17599 17523 17633
rect 17523 17599 17549 17633
rect 17497 17590 17549 17599
rect 17561 17633 17613 17642
rect 17625 17633 17677 17642
rect 17689 17633 17741 17642
rect 17561 17599 17581 17633
rect 17581 17599 17613 17633
rect 17625 17599 17673 17633
rect 17673 17599 17677 17633
rect 17689 17599 17707 17633
rect 17707 17599 17741 17633
rect 17561 17590 17613 17599
rect 17625 17590 17677 17599
rect 17689 17590 17741 17599
rect 17753 17633 17805 17642
rect 17753 17599 17765 17633
rect 17765 17599 17799 17633
rect 17799 17599 17805 17633
rect 17753 17590 17805 17599
rect 6703 17089 6755 17098
rect 6767 17089 6819 17098
rect 6831 17089 6883 17098
rect 6703 17055 6725 17089
rect 6725 17055 6755 17089
rect 6767 17055 6817 17089
rect 6817 17055 6819 17089
rect 6831 17055 6851 17089
rect 6851 17055 6883 17089
rect 6703 17046 6755 17055
rect 6767 17046 6819 17055
rect 6831 17046 6883 17055
rect 6895 17089 6947 17098
rect 6895 17055 6909 17089
rect 6909 17055 6943 17089
rect 6943 17055 6947 17089
rect 6895 17046 6947 17055
rect 6959 17089 7011 17098
rect 10521 17089 10573 17098
rect 6959 17055 7001 17089
rect 7001 17055 7011 17089
rect 10521 17055 10531 17089
rect 10531 17055 10573 17089
rect 6959 17046 7011 17055
rect 10521 17046 10573 17055
rect 10585 17089 10637 17098
rect 10585 17055 10589 17089
rect 10589 17055 10623 17089
rect 10623 17055 10637 17089
rect 10585 17046 10637 17055
rect 10649 17089 10701 17098
rect 10713 17089 10765 17098
rect 10777 17089 10829 17098
rect 14339 17089 14391 17098
rect 14403 17089 14455 17098
rect 14467 17089 14519 17098
rect 10649 17055 10681 17089
rect 10681 17055 10701 17089
rect 10713 17055 10715 17089
rect 10715 17055 10765 17089
rect 10777 17055 10807 17089
rect 10807 17055 10829 17089
rect 14339 17055 14361 17089
rect 14361 17055 14391 17089
rect 14403 17055 14453 17089
rect 14453 17055 14455 17089
rect 14467 17055 14487 17089
rect 14487 17055 14519 17089
rect 10649 17046 10701 17055
rect 10713 17046 10765 17055
rect 10777 17046 10829 17055
rect 14339 17046 14391 17055
rect 14403 17046 14455 17055
rect 14467 17046 14519 17055
rect 14531 17089 14583 17098
rect 14531 17055 14545 17089
rect 14545 17055 14579 17089
rect 14579 17055 14583 17089
rect 14531 17046 14583 17055
rect 14595 17089 14647 17098
rect 18157 17089 18209 17098
rect 14595 17055 14637 17089
rect 14637 17055 14647 17089
rect 18157 17055 18167 17089
rect 18167 17055 18209 17089
rect 14595 17046 14647 17055
rect 18157 17046 18209 17055
rect 18221 17089 18273 17098
rect 18221 17055 18225 17089
rect 18225 17055 18259 17089
rect 18259 17055 18273 17089
rect 18221 17046 18273 17055
rect 18285 17089 18337 17098
rect 18349 17089 18401 17098
rect 18413 17089 18465 17098
rect 18285 17055 18317 17089
rect 18317 17055 18337 17089
rect 18349 17055 18351 17089
rect 18351 17055 18401 17089
rect 18413 17055 18443 17089
rect 18443 17055 18465 17089
rect 18285 17046 18337 17055
rect 18349 17046 18401 17055
rect 18413 17046 18465 17055
rect 6043 16545 6095 16554
rect 6107 16545 6159 16554
rect 6043 16511 6081 16545
rect 6081 16511 6095 16545
rect 6107 16511 6115 16545
rect 6115 16511 6159 16545
rect 6043 16502 6095 16511
rect 6107 16502 6159 16511
rect 6171 16545 6223 16554
rect 6171 16511 6173 16545
rect 6173 16511 6207 16545
rect 6207 16511 6223 16545
rect 6171 16502 6223 16511
rect 6235 16545 6287 16554
rect 6235 16511 6265 16545
rect 6265 16511 6287 16545
rect 6235 16502 6287 16511
rect 6299 16502 6351 16554
rect 9861 16545 9913 16554
rect 9861 16511 9887 16545
rect 9887 16511 9913 16545
rect 9861 16502 9913 16511
rect 9925 16545 9977 16554
rect 9989 16545 10041 16554
rect 10053 16545 10105 16554
rect 9925 16511 9945 16545
rect 9945 16511 9977 16545
rect 9989 16511 10037 16545
rect 10037 16511 10041 16545
rect 10053 16511 10071 16545
rect 10071 16511 10105 16545
rect 9925 16502 9977 16511
rect 9989 16502 10041 16511
rect 10053 16502 10105 16511
rect 10117 16545 10169 16554
rect 13679 16545 13731 16554
rect 13743 16545 13795 16554
rect 10117 16511 10129 16545
rect 10129 16511 10163 16545
rect 10163 16511 10169 16545
rect 13679 16511 13717 16545
rect 13717 16511 13731 16545
rect 13743 16511 13751 16545
rect 13751 16511 13795 16545
rect 10117 16502 10169 16511
rect 13679 16502 13731 16511
rect 13743 16502 13795 16511
rect 13807 16545 13859 16554
rect 13807 16511 13809 16545
rect 13809 16511 13843 16545
rect 13843 16511 13859 16545
rect 13807 16502 13859 16511
rect 13871 16545 13923 16554
rect 13871 16511 13901 16545
rect 13901 16511 13923 16545
rect 13871 16502 13923 16511
rect 13935 16502 13987 16554
rect 17497 16545 17549 16554
rect 17497 16511 17523 16545
rect 17523 16511 17549 16545
rect 17497 16502 17549 16511
rect 17561 16545 17613 16554
rect 17625 16545 17677 16554
rect 17689 16545 17741 16554
rect 17561 16511 17581 16545
rect 17581 16511 17613 16545
rect 17625 16511 17673 16545
rect 17673 16511 17677 16545
rect 17689 16511 17707 16545
rect 17707 16511 17741 16545
rect 17561 16502 17613 16511
rect 17625 16502 17677 16511
rect 17689 16502 17741 16511
rect 17753 16545 17805 16554
rect 17753 16511 17765 16545
rect 17765 16511 17799 16545
rect 17799 16511 17805 16545
rect 17753 16502 17805 16511
rect 6703 16001 6755 16010
rect 6767 16001 6819 16010
rect 6831 16001 6883 16010
rect 6703 15967 6725 16001
rect 6725 15967 6755 16001
rect 6767 15967 6817 16001
rect 6817 15967 6819 16001
rect 6831 15967 6851 16001
rect 6851 15967 6883 16001
rect 6703 15958 6755 15967
rect 6767 15958 6819 15967
rect 6831 15958 6883 15967
rect 6895 16001 6947 16010
rect 6895 15967 6909 16001
rect 6909 15967 6943 16001
rect 6943 15967 6947 16001
rect 6895 15958 6947 15967
rect 6959 16001 7011 16010
rect 10521 16001 10573 16010
rect 6959 15967 7001 16001
rect 7001 15967 7011 16001
rect 10521 15967 10531 16001
rect 10531 15967 10573 16001
rect 6959 15958 7011 15967
rect 10521 15958 10573 15967
rect 10585 16001 10637 16010
rect 10585 15967 10589 16001
rect 10589 15967 10623 16001
rect 10623 15967 10637 16001
rect 10585 15958 10637 15967
rect 10649 16001 10701 16010
rect 10713 16001 10765 16010
rect 10777 16001 10829 16010
rect 14339 16001 14391 16010
rect 14403 16001 14455 16010
rect 14467 16001 14519 16010
rect 10649 15967 10681 16001
rect 10681 15967 10701 16001
rect 10713 15967 10715 16001
rect 10715 15967 10765 16001
rect 10777 15967 10807 16001
rect 10807 15967 10829 16001
rect 14339 15967 14361 16001
rect 14361 15967 14391 16001
rect 14403 15967 14453 16001
rect 14453 15967 14455 16001
rect 14467 15967 14487 16001
rect 14487 15967 14519 16001
rect 10649 15958 10701 15967
rect 10713 15958 10765 15967
rect 10777 15958 10829 15967
rect 14339 15958 14391 15967
rect 14403 15958 14455 15967
rect 14467 15958 14519 15967
rect 14531 16001 14583 16010
rect 14531 15967 14545 16001
rect 14545 15967 14579 16001
rect 14579 15967 14583 16001
rect 14531 15958 14583 15967
rect 14595 16001 14647 16010
rect 18157 16001 18209 16010
rect 14595 15967 14637 16001
rect 14637 15967 14647 16001
rect 18157 15967 18167 16001
rect 18167 15967 18209 16001
rect 14595 15958 14647 15967
rect 18157 15958 18209 15967
rect 18221 16001 18273 16010
rect 18221 15967 18225 16001
rect 18225 15967 18259 16001
rect 18259 15967 18273 16001
rect 18221 15958 18273 15967
rect 18285 16001 18337 16010
rect 18349 16001 18401 16010
rect 18413 16001 18465 16010
rect 18285 15967 18317 16001
rect 18317 15967 18337 16001
rect 18349 15967 18351 16001
rect 18351 15967 18401 16001
rect 18413 15967 18443 16001
rect 18443 15967 18465 16001
rect 18285 15958 18337 15967
rect 18349 15958 18401 15967
rect 18413 15958 18465 15967
rect 6043 15457 6095 15466
rect 6107 15457 6159 15466
rect 6043 15423 6081 15457
rect 6081 15423 6095 15457
rect 6107 15423 6115 15457
rect 6115 15423 6159 15457
rect 6043 15414 6095 15423
rect 6107 15414 6159 15423
rect 6171 15457 6223 15466
rect 6171 15423 6173 15457
rect 6173 15423 6207 15457
rect 6207 15423 6223 15457
rect 6171 15414 6223 15423
rect 6235 15457 6287 15466
rect 6235 15423 6265 15457
rect 6265 15423 6287 15457
rect 6235 15414 6287 15423
rect 6299 15414 6351 15466
rect 9861 15457 9913 15466
rect 9861 15423 9887 15457
rect 9887 15423 9913 15457
rect 9861 15414 9913 15423
rect 9925 15457 9977 15466
rect 9989 15457 10041 15466
rect 10053 15457 10105 15466
rect 9925 15423 9945 15457
rect 9945 15423 9977 15457
rect 9989 15423 10037 15457
rect 10037 15423 10041 15457
rect 10053 15423 10071 15457
rect 10071 15423 10105 15457
rect 9925 15414 9977 15423
rect 9989 15414 10041 15423
rect 10053 15414 10105 15423
rect 10117 15457 10169 15466
rect 13679 15457 13731 15466
rect 13743 15457 13795 15466
rect 10117 15423 10129 15457
rect 10129 15423 10163 15457
rect 10163 15423 10169 15457
rect 13679 15423 13717 15457
rect 13717 15423 13731 15457
rect 13743 15423 13751 15457
rect 13751 15423 13795 15457
rect 10117 15414 10169 15423
rect 13679 15414 13731 15423
rect 13743 15414 13795 15423
rect 13807 15457 13859 15466
rect 13807 15423 13809 15457
rect 13809 15423 13843 15457
rect 13843 15423 13859 15457
rect 13807 15414 13859 15423
rect 13871 15457 13923 15466
rect 13871 15423 13901 15457
rect 13901 15423 13923 15457
rect 13871 15414 13923 15423
rect 13935 15414 13987 15466
rect 17497 15457 17549 15466
rect 17497 15423 17523 15457
rect 17523 15423 17549 15457
rect 17497 15414 17549 15423
rect 17561 15457 17613 15466
rect 17625 15457 17677 15466
rect 17689 15457 17741 15466
rect 17561 15423 17581 15457
rect 17581 15423 17613 15457
rect 17625 15423 17673 15457
rect 17673 15423 17677 15457
rect 17689 15423 17707 15457
rect 17707 15423 17741 15457
rect 17561 15414 17613 15423
rect 17625 15414 17677 15423
rect 17689 15414 17741 15423
rect 17753 15457 17805 15466
rect 17753 15423 17765 15457
rect 17765 15423 17799 15457
rect 17799 15423 17805 15457
rect 17753 15414 17805 15423
rect 12880 15151 12932 15160
rect 12880 15117 12889 15151
rect 12889 15117 12923 15151
rect 12923 15117 12932 15151
rect 12880 15108 12932 15117
rect 15364 15151 15416 15160
rect 15364 15117 15373 15151
rect 15373 15117 15407 15151
rect 15407 15117 15416 15151
rect 15364 15108 15416 15117
rect 13432 15015 13484 15024
rect 13432 14981 13441 15015
rect 13441 14981 13475 15015
rect 13475 14981 13484 15015
rect 13432 14972 13484 14981
rect 16100 14972 16152 15024
rect 6703 14913 6755 14922
rect 6767 14913 6819 14922
rect 6831 14913 6883 14922
rect 6703 14879 6725 14913
rect 6725 14879 6755 14913
rect 6767 14879 6817 14913
rect 6817 14879 6819 14913
rect 6831 14879 6851 14913
rect 6851 14879 6883 14913
rect 6703 14870 6755 14879
rect 6767 14870 6819 14879
rect 6831 14870 6883 14879
rect 6895 14913 6947 14922
rect 6895 14879 6909 14913
rect 6909 14879 6943 14913
rect 6943 14879 6947 14913
rect 6895 14870 6947 14879
rect 6959 14913 7011 14922
rect 10521 14913 10573 14922
rect 6959 14879 7001 14913
rect 7001 14879 7011 14913
rect 10521 14879 10531 14913
rect 10531 14879 10573 14913
rect 6959 14870 7011 14879
rect 10521 14870 10573 14879
rect 10585 14913 10637 14922
rect 10585 14879 10589 14913
rect 10589 14879 10623 14913
rect 10623 14879 10637 14913
rect 10585 14870 10637 14879
rect 10649 14913 10701 14922
rect 10713 14913 10765 14922
rect 10777 14913 10829 14922
rect 14339 14913 14391 14922
rect 14403 14913 14455 14922
rect 14467 14913 14519 14922
rect 10649 14879 10681 14913
rect 10681 14879 10701 14913
rect 10713 14879 10715 14913
rect 10715 14879 10765 14913
rect 10777 14879 10807 14913
rect 10807 14879 10829 14913
rect 14339 14879 14361 14913
rect 14361 14879 14391 14913
rect 14403 14879 14453 14913
rect 14453 14879 14455 14913
rect 14467 14879 14487 14913
rect 14487 14879 14519 14913
rect 10649 14870 10701 14879
rect 10713 14870 10765 14879
rect 10777 14870 10829 14879
rect 14339 14870 14391 14879
rect 14403 14870 14455 14879
rect 14467 14870 14519 14879
rect 14531 14913 14583 14922
rect 14531 14879 14545 14913
rect 14545 14879 14579 14913
rect 14579 14879 14583 14913
rect 14531 14870 14583 14879
rect 14595 14913 14647 14922
rect 18157 14913 18209 14922
rect 14595 14879 14637 14913
rect 14637 14879 14647 14913
rect 18157 14879 18167 14913
rect 18167 14879 18209 14913
rect 14595 14870 14647 14879
rect 18157 14870 18209 14879
rect 18221 14913 18273 14922
rect 18221 14879 18225 14913
rect 18225 14879 18259 14913
rect 18259 14879 18273 14913
rect 18221 14870 18273 14879
rect 18285 14913 18337 14922
rect 18349 14913 18401 14922
rect 18413 14913 18465 14922
rect 18285 14879 18317 14913
rect 18317 14879 18337 14913
rect 18349 14879 18351 14913
rect 18351 14879 18401 14913
rect 18413 14879 18443 14913
rect 18443 14879 18465 14913
rect 18285 14870 18337 14879
rect 18349 14870 18401 14879
rect 18413 14870 18465 14879
rect 11684 14632 11736 14684
rect 11040 14607 11092 14616
rect 11040 14573 11049 14607
rect 11049 14573 11083 14607
rect 11083 14573 11092 14607
rect 11040 14564 11092 14573
rect 13432 14768 13484 14820
rect 14996 14700 15048 14752
rect 14260 14607 14312 14616
rect 14260 14573 14269 14607
rect 14269 14573 14303 14607
rect 14303 14573 14312 14607
rect 14260 14564 14312 14573
rect 16284 14607 16336 14616
rect 16284 14573 16293 14607
rect 16293 14573 16327 14607
rect 16327 14573 16336 14607
rect 16284 14564 16336 14573
rect 15548 14539 15600 14548
rect 15548 14505 15561 14539
rect 15561 14505 15595 14539
rect 15595 14505 15600 14539
rect 15548 14496 15600 14505
rect 16008 14539 16060 14548
rect 16008 14505 16017 14539
rect 16017 14505 16051 14539
rect 16051 14505 16060 14539
rect 16008 14496 16060 14505
rect 10212 14428 10264 14480
rect 11408 14471 11460 14480
rect 11408 14437 11417 14471
rect 11417 14437 11451 14471
rect 11451 14437 11460 14471
rect 11408 14428 11460 14437
rect 13064 14428 13116 14480
rect 13432 14471 13484 14480
rect 13432 14437 13441 14471
rect 13441 14437 13475 14471
rect 13475 14437 13484 14471
rect 13432 14428 13484 14437
rect 14352 14428 14404 14480
rect 15640 14428 15692 14480
rect 6043 14369 6095 14378
rect 6107 14369 6159 14378
rect 6043 14335 6081 14369
rect 6081 14335 6095 14369
rect 6107 14335 6115 14369
rect 6115 14335 6159 14369
rect 6043 14326 6095 14335
rect 6107 14326 6159 14335
rect 6171 14369 6223 14378
rect 6171 14335 6173 14369
rect 6173 14335 6207 14369
rect 6207 14335 6223 14369
rect 6171 14326 6223 14335
rect 6235 14369 6287 14378
rect 6235 14335 6265 14369
rect 6265 14335 6287 14369
rect 6235 14326 6287 14335
rect 6299 14326 6351 14378
rect 9861 14369 9913 14378
rect 9861 14335 9887 14369
rect 9887 14335 9913 14369
rect 9861 14326 9913 14335
rect 9925 14369 9977 14378
rect 9989 14369 10041 14378
rect 10053 14369 10105 14378
rect 9925 14335 9945 14369
rect 9945 14335 9977 14369
rect 9989 14335 10037 14369
rect 10037 14335 10041 14369
rect 10053 14335 10071 14369
rect 10071 14335 10105 14369
rect 9925 14326 9977 14335
rect 9989 14326 10041 14335
rect 10053 14326 10105 14335
rect 10117 14369 10169 14378
rect 13679 14369 13731 14378
rect 13743 14369 13795 14378
rect 10117 14335 10129 14369
rect 10129 14335 10163 14369
rect 10163 14335 10169 14369
rect 13679 14335 13717 14369
rect 13717 14335 13731 14369
rect 13743 14335 13751 14369
rect 13751 14335 13795 14369
rect 10117 14326 10169 14335
rect 13679 14326 13731 14335
rect 13743 14326 13795 14335
rect 13807 14369 13859 14378
rect 13807 14335 13809 14369
rect 13809 14335 13843 14369
rect 13843 14335 13859 14369
rect 13807 14326 13859 14335
rect 13871 14369 13923 14378
rect 13871 14335 13901 14369
rect 13901 14335 13923 14369
rect 13871 14326 13923 14335
rect 13935 14326 13987 14378
rect 17497 14369 17549 14378
rect 17497 14335 17523 14369
rect 17523 14335 17549 14369
rect 17497 14326 17549 14335
rect 17561 14369 17613 14378
rect 17625 14369 17677 14378
rect 17689 14369 17741 14378
rect 17561 14335 17581 14369
rect 17581 14335 17613 14369
rect 17625 14335 17673 14369
rect 17673 14335 17677 14369
rect 17689 14335 17707 14369
rect 17707 14335 17741 14369
rect 17561 14326 17613 14335
rect 17625 14326 17677 14335
rect 17689 14326 17741 14335
rect 17753 14369 17805 14378
rect 17753 14335 17765 14369
rect 17765 14335 17799 14369
rect 17799 14335 17805 14369
rect 17753 14326 17805 14335
rect 11408 14224 11460 14276
rect 15364 14224 15416 14276
rect 15640 14267 15692 14276
rect 15640 14233 15649 14267
rect 15649 14233 15683 14267
rect 15683 14233 15692 14267
rect 15640 14224 15692 14233
rect 16008 14267 16060 14276
rect 16008 14233 16017 14267
rect 16017 14233 16051 14267
rect 16051 14233 16060 14267
rect 16008 14224 16060 14233
rect 16100 14224 16152 14276
rect 5796 14156 5848 14208
rect 13984 14199 14036 14208
rect 13984 14165 13993 14199
rect 13993 14165 14027 14199
rect 14027 14165 14036 14199
rect 13984 14156 14036 14165
rect 16468 14131 16520 14140
rect 16468 14097 16477 14131
rect 16477 14097 16511 14131
rect 16511 14097 16520 14131
rect 16468 14088 16520 14097
rect 10856 14020 10908 14072
rect 10212 13884 10264 13936
rect 11868 14063 11920 14072
rect 11868 14029 11877 14063
rect 11877 14029 11911 14063
rect 11911 14029 11920 14063
rect 11868 14020 11920 14029
rect 14168 14020 14220 14072
rect 14352 14020 14404 14072
rect 14812 14020 14864 14072
rect 12696 13927 12748 13936
rect 12696 13893 12705 13927
rect 12705 13893 12739 13927
rect 12739 13893 12748 13927
rect 12696 13884 12748 13893
rect 14720 13884 14772 13936
rect 15732 13884 15784 13936
rect 17112 13884 17164 13936
rect 6703 13825 6755 13834
rect 6767 13825 6819 13834
rect 6831 13825 6883 13834
rect 6703 13791 6725 13825
rect 6725 13791 6755 13825
rect 6767 13791 6817 13825
rect 6817 13791 6819 13825
rect 6831 13791 6851 13825
rect 6851 13791 6883 13825
rect 6703 13782 6755 13791
rect 6767 13782 6819 13791
rect 6831 13782 6883 13791
rect 6895 13825 6947 13834
rect 6895 13791 6909 13825
rect 6909 13791 6943 13825
rect 6943 13791 6947 13825
rect 6895 13782 6947 13791
rect 6959 13825 7011 13834
rect 10521 13825 10573 13834
rect 6959 13791 7001 13825
rect 7001 13791 7011 13825
rect 10521 13791 10531 13825
rect 10531 13791 10573 13825
rect 6959 13782 7011 13791
rect 10521 13782 10573 13791
rect 10585 13825 10637 13834
rect 10585 13791 10589 13825
rect 10589 13791 10623 13825
rect 10623 13791 10637 13825
rect 10585 13782 10637 13791
rect 10649 13825 10701 13834
rect 10713 13825 10765 13834
rect 10777 13825 10829 13834
rect 14339 13825 14391 13834
rect 14403 13825 14455 13834
rect 14467 13825 14519 13834
rect 10649 13791 10681 13825
rect 10681 13791 10701 13825
rect 10713 13791 10715 13825
rect 10715 13791 10765 13825
rect 10777 13791 10807 13825
rect 10807 13791 10829 13825
rect 14339 13791 14361 13825
rect 14361 13791 14391 13825
rect 14403 13791 14453 13825
rect 14453 13791 14455 13825
rect 14467 13791 14487 13825
rect 14487 13791 14519 13825
rect 10649 13782 10701 13791
rect 10713 13782 10765 13791
rect 10777 13782 10829 13791
rect 14339 13782 14391 13791
rect 14403 13782 14455 13791
rect 14467 13782 14519 13791
rect 14531 13825 14583 13834
rect 14531 13791 14545 13825
rect 14545 13791 14579 13825
rect 14579 13791 14583 13825
rect 14531 13782 14583 13791
rect 14595 13825 14647 13834
rect 18157 13825 18209 13834
rect 14595 13791 14637 13825
rect 14637 13791 14647 13825
rect 18157 13791 18167 13825
rect 18167 13791 18209 13825
rect 14595 13782 14647 13791
rect 18157 13782 18209 13791
rect 18221 13825 18273 13834
rect 18221 13791 18225 13825
rect 18225 13791 18259 13825
rect 18259 13791 18273 13825
rect 18221 13782 18273 13791
rect 18285 13825 18337 13834
rect 18349 13825 18401 13834
rect 18413 13825 18465 13834
rect 18285 13791 18317 13825
rect 18317 13791 18337 13825
rect 18349 13791 18351 13825
rect 18351 13791 18401 13825
rect 18413 13791 18443 13825
rect 18443 13791 18465 13825
rect 18285 13782 18337 13791
rect 18349 13782 18401 13791
rect 18413 13782 18465 13791
rect 11868 13680 11920 13732
rect 12696 13680 12748 13732
rect 13064 13680 13116 13732
rect 9660 13519 9712 13528
rect 9660 13485 9669 13519
rect 9669 13485 9703 13519
rect 9703 13485 9712 13519
rect 9660 13476 9712 13485
rect 10856 13476 10908 13528
rect 15088 13544 15140 13596
rect 16284 13680 16336 13732
rect 16468 13680 16520 13732
rect 17112 13587 17164 13596
rect 17112 13553 17121 13587
rect 17121 13553 17155 13587
rect 17155 13553 17164 13587
rect 17112 13544 17164 13553
rect 18768 13544 18820 13596
rect 12696 13519 12748 13528
rect 12696 13485 12705 13519
rect 12705 13485 12739 13519
rect 12739 13485 12748 13519
rect 12696 13476 12748 13485
rect 14720 13519 14772 13528
rect 14720 13485 14729 13519
rect 14729 13485 14763 13519
rect 14763 13485 14772 13519
rect 14720 13476 14772 13485
rect 15640 13476 15692 13528
rect 16928 13519 16980 13528
rect 16928 13485 16937 13519
rect 16937 13485 16971 13519
rect 16971 13485 16980 13519
rect 16928 13476 16980 13485
rect 10580 13340 10632 13392
rect 12512 13383 12564 13392
rect 12512 13349 12521 13383
rect 12521 13349 12555 13383
rect 12555 13349 12564 13383
rect 12512 13340 12564 13349
rect 14076 13408 14128 13460
rect 14444 13340 14496 13392
rect 17020 13383 17072 13392
rect 17020 13349 17029 13383
rect 17029 13349 17063 13383
rect 17063 13349 17072 13383
rect 17020 13340 17072 13349
rect 6043 13281 6095 13290
rect 6107 13281 6159 13290
rect 6043 13247 6081 13281
rect 6081 13247 6095 13281
rect 6107 13247 6115 13281
rect 6115 13247 6159 13281
rect 6043 13238 6095 13247
rect 6107 13238 6159 13247
rect 6171 13281 6223 13290
rect 6171 13247 6173 13281
rect 6173 13247 6207 13281
rect 6207 13247 6223 13281
rect 6171 13238 6223 13247
rect 6235 13281 6287 13290
rect 6235 13247 6265 13281
rect 6265 13247 6287 13281
rect 6235 13238 6287 13247
rect 6299 13238 6351 13290
rect 9861 13281 9913 13290
rect 9861 13247 9887 13281
rect 9887 13247 9913 13281
rect 9861 13238 9913 13247
rect 9925 13281 9977 13290
rect 9989 13281 10041 13290
rect 10053 13281 10105 13290
rect 9925 13247 9945 13281
rect 9945 13247 9977 13281
rect 9989 13247 10037 13281
rect 10037 13247 10041 13281
rect 10053 13247 10071 13281
rect 10071 13247 10105 13281
rect 9925 13238 9977 13247
rect 9989 13238 10041 13247
rect 10053 13238 10105 13247
rect 10117 13281 10169 13290
rect 13679 13281 13731 13290
rect 13743 13281 13795 13290
rect 10117 13247 10129 13281
rect 10129 13247 10163 13281
rect 10163 13247 10169 13281
rect 13679 13247 13717 13281
rect 13717 13247 13731 13281
rect 13743 13247 13751 13281
rect 13751 13247 13795 13281
rect 10117 13238 10169 13247
rect 13679 13238 13731 13247
rect 13743 13238 13795 13247
rect 13807 13281 13859 13290
rect 13807 13247 13809 13281
rect 13809 13247 13843 13281
rect 13843 13247 13859 13281
rect 13807 13238 13859 13247
rect 13871 13281 13923 13290
rect 13871 13247 13901 13281
rect 13901 13247 13923 13281
rect 13871 13238 13923 13247
rect 13935 13238 13987 13290
rect 17497 13281 17549 13290
rect 17497 13247 17523 13281
rect 17523 13247 17549 13281
rect 17497 13238 17549 13247
rect 17561 13281 17613 13290
rect 17625 13281 17677 13290
rect 17689 13281 17741 13290
rect 17561 13247 17581 13281
rect 17581 13247 17613 13281
rect 17625 13247 17673 13281
rect 17673 13247 17677 13281
rect 17689 13247 17707 13281
rect 17707 13247 17741 13281
rect 17561 13238 17613 13247
rect 17625 13238 17677 13247
rect 17689 13238 17741 13247
rect 17753 13281 17805 13290
rect 17753 13247 17765 13281
rect 17765 13247 17799 13281
rect 17799 13247 17805 13281
rect 17753 13238 17805 13247
rect 10580 13136 10632 13188
rect 11868 13136 11920 13188
rect 9200 12975 9252 12984
rect 9200 12941 9209 12975
rect 9209 12941 9243 12975
rect 9243 12941 9252 12975
rect 9200 12932 9252 12941
rect 10856 13068 10908 13120
rect 14444 13136 14496 13188
rect 14720 13068 14772 13120
rect 14812 13068 14864 13120
rect 14996 13068 15048 13120
rect 16284 13136 16336 13188
rect 17020 13136 17072 13188
rect 12512 12975 12564 12984
rect 12512 12941 12521 12975
rect 12521 12941 12555 12975
rect 12555 12941 12564 12975
rect 12512 12932 12564 12941
rect 13064 12932 13116 12984
rect 15548 13000 15600 13052
rect 17572 12975 17624 12984
rect 17572 12941 17581 12975
rect 17581 12941 17615 12975
rect 17615 12941 17624 12975
rect 17572 12932 17624 12941
rect 14260 12864 14312 12916
rect 9752 12839 9804 12848
rect 9752 12805 9761 12839
rect 9761 12805 9795 12839
rect 9795 12805 9804 12839
rect 9752 12796 9804 12805
rect 10212 12796 10264 12848
rect 11500 12796 11552 12848
rect 12880 12796 12932 12848
rect 14168 12796 14220 12848
rect 6703 12737 6755 12746
rect 6767 12737 6819 12746
rect 6831 12737 6883 12746
rect 6703 12703 6725 12737
rect 6725 12703 6755 12737
rect 6767 12703 6817 12737
rect 6817 12703 6819 12737
rect 6831 12703 6851 12737
rect 6851 12703 6883 12737
rect 6703 12694 6755 12703
rect 6767 12694 6819 12703
rect 6831 12694 6883 12703
rect 6895 12737 6947 12746
rect 6895 12703 6909 12737
rect 6909 12703 6943 12737
rect 6943 12703 6947 12737
rect 6895 12694 6947 12703
rect 6959 12737 7011 12746
rect 10521 12737 10573 12746
rect 6959 12703 7001 12737
rect 7001 12703 7011 12737
rect 10521 12703 10531 12737
rect 10531 12703 10573 12737
rect 6959 12694 7011 12703
rect 10521 12694 10573 12703
rect 10585 12737 10637 12746
rect 10585 12703 10589 12737
rect 10589 12703 10623 12737
rect 10623 12703 10637 12737
rect 10585 12694 10637 12703
rect 10649 12737 10701 12746
rect 10713 12737 10765 12746
rect 10777 12737 10829 12746
rect 14339 12737 14391 12746
rect 14403 12737 14455 12746
rect 14467 12737 14519 12746
rect 10649 12703 10681 12737
rect 10681 12703 10701 12737
rect 10713 12703 10715 12737
rect 10715 12703 10765 12737
rect 10777 12703 10807 12737
rect 10807 12703 10829 12737
rect 14339 12703 14361 12737
rect 14361 12703 14391 12737
rect 14403 12703 14453 12737
rect 14453 12703 14455 12737
rect 14467 12703 14487 12737
rect 14487 12703 14519 12737
rect 10649 12694 10701 12703
rect 10713 12694 10765 12703
rect 10777 12694 10829 12703
rect 14339 12694 14391 12703
rect 14403 12694 14455 12703
rect 14467 12694 14519 12703
rect 14531 12737 14583 12746
rect 14531 12703 14545 12737
rect 14545 12703 14579 12737
rect 14579 12703 14583 12737
rect 14531 12694 14583 12703
rect 14595 12737 14647 12746
rect 18157 12737 18209 12746
rect 14595 12703 14637 12737
rect 14637 12703 14647 12737
rect 18157 12703 18167 12737
rect 18167 12703 18209 12737
rect 14595 12694 14647 12703
rect 18157 12694 18209 12703
rect 18221 12737 18273 12746
rect 18221 12703 18225 12737
rect 18225 12703 18259 12737
rect 18259 12703 18273 12737
rect 18221 12694 18273 12703
rect 18285 12737 18337 12746
rect 18349 12737 18401 12746
rect 18413 12737 18465 12746
rect 18285 12703 18317 12737
rect 18317 12703 18337 12737
rect 18349 12703 18351 12737
rect 18351 12703 18401 12737
rect 18413 12703 18443 12737
rect 18443 12703 18465 12737
rect 18285 12694 18337 12703
rect 18349 12694 18401 12703
rect 18413 12694 18465 12703
rect 9660 12592 9712 12644
rect 10212 12635 10264 12644
rect 10212 12601 10221 12635
rect 10221 12601 10255 12635
rect 10255 12601 10264 12635
rect 10212 12592 10264 12601
rect 12696 12592 12748 12644
rect 14076 12592 14128 12644
rect 14720 12635 14772 12644
rect 14720 12601 14729 12635
rect 14729 12601 14763 12635
rect 14763 12601 14772 12635
rect 14720 12592 14772 12601
rect 9752 12456 9804 12508
rect 5244 12431 5296 12440
rect 5244 12397 5253 12431
rect 5253 12397 5287 12431
rect 5287 12397 5296 12431
rect 5244 12388 5296 12397
rect 9200 12431 9252 12440
rect 9200 12397 9209 12431
rect 9209 12397 9243 12431
rect 9243 12397 9252 12431
rect 9200 12388 9252 12397
rect 10120 12388 10172 12440
rect 11684 12456 11736 12508
rect 14168 12499 14220 12508
rect 14168 12465 14177 12499
rect 14177 12465 14211 12499
rect 14211 12465 14220 12499
rect 14168 12456 14220 12465
rect 15088 12499 15140 12508
rect 15088 12465 15097 12499
rect 15097 12465 15131 12499
rect 15131 12465 15140 12499
rect 15088 12456 15140 12465
rect 15732 12456 15784 12508
rect 13156 12388 13208 12440
rect 13432 12388 13484 12440
rect 7268 12252 7320 12304
rect 9384 12252 9436 12304
rect 12880 12252 12932 12304
rect 15640 12320 15692 12372
rect 16928 12388 16980 12440
rect 17572 12388 17624 12440
rect 13616 12295 13668 12304
rect 13616 12261 13625 12295
rect 13625 12261 13659 12295
rect 13659 12261 13668 12295
rect 13616 12252 13668 12261
rect 15548 12252 15600 12304
rect 17848 12320 17900 12372
rect 19964 12320 20016 12372
rect 6043 12193 6095 12202
rect 6107 12193 6159 12202
rect 6043 12159 6081 12193
rect 6081 12159 6095 12193
rect 6107 12159 6115 12193
rect 6115 12159 6159 12193
rect 6043 12150 6095 12159
rect 6107 12150 6159 12159
rect 6171 12193 6223 12202
rect 6171 12159 6173 12193
rect 6173 12159 6207 12193
rect 6207 12159 6223 12193
rect 6171 12150 6223 12159
rect 6235 12193 6287 12202
rect 6235 12159 6265 12193
rect 6265 12159 6287 12193
rect 6235 12150 6287 12159
rect 6299 12150 6351 12202
rect 9861 12193 9913 12202
rect 9861 12159 9887 12193
rect 9887 12159 9913 12193
rect 9861 12150 9913 12159
rect 9925 12193 9977 12202
rect 9989 12193 10041 12202
rect 10053 12193 10105 12202
rect 9925 12159 9945 12193
rect 9945 12159 9977 12193
rect 9989 12159 10037 12193
rect 10037 12159 10041 12193
rect 10053 12159 10071 12193
rect 10071 12159 10105 12193
rect 9925 12150 9977 12159
rect 9989 12150 10041 12159
rect 10053 12150 10105 12159
rect 10117 12193 10169 12202
rect 13679 12193 13731 12202
rect 13743 12193 13795 12202
rect 10117 12159 10129 12193
rect 10129 12159 10163 12193
rect 10163 12159 10169 12193
rect 13679 12159 13717 12193
rect 13717 12159 13731 12193
rect 13743 12159 13751 12193
rect 13751 12159 13795 12193
rect 10117 12150 10169 12159
rect 13679 12150 13731 12159
rect 13743 12150 13795 12159
rect 13807 12193 13859 12202
rect 13807 12159 13809 12193
rect 13809 12159 13843 12193
rect 13843 12159 13859 12193
rect 13807 12150 13859 12159
rect 13871 12193 13923 12202
rect 13871 12159 13901 12193
rect 13901 12159 13923 12193
rect 13871 12150 13923 12159
rect 13935 12150 13987 12202
rect 17497 12193 17549 12202
rect 17497 12159 17523 12193
rect 17523 12159 17549 12193
rect 17497 12150 17549 12159
rect 17561 12193 17613 12202
rect 17625 12193 17677 12202
rect 17689 12193 17741 12202
rect 17561 12159 17581 12193
rect 17581 12159 17613 12193
rect 17625 12159 17673 12193
rect 17673 12159 17677 12193
rect 17689 12159 17707 12193
rect 17707 12159 17741 12193
rect 17561 12150 17613 12159
rect 17625 12150 17677 12159
rect 17689 12150 17741 12159
rect 17753 12193 17805 12202
rect 17753 12159 17765 12193
rect 17765 12159 17799 12193
rect 17799 12159 17805 12193
rect 17753 12150 17805 12159
rect 5160 10020 5260 10160
rect 430 3450 610 3630
rect 440 2510 620 2690
rect 7240 9980 7370 10150
rect 9340 10020 9470 10190
rect 3430 6480 3650 6720
rect 1050 3440 1230 3620
rect 1890 3950 2030 4050
rect 1060 2510 1240 2690
rect 1930 2000 1951 2100
rect 1951 2000 1985 2100
rect 1985 2000 2040 2100
rect 1930 1880 1951 1980
rect 1951 1880 1985 1980
rect 1985 1880 2040 1980
rect 1930 1760 1951 1860
rect 1951 1760 1985 1860
rect 1985 1760 2040 1860
rect 11430 10020 11560 10190
rect 13600 10020 13730 10190
rect 6730 6490 6940 6610
rect 4360 3450 4540 3630
rect 5190 3950 5330 4050
rect 4350 2510 4530 2690
rect 5230 2000 5251 2100
rect 5251 2000 5285 2100
rect 5285 2000 5340 2100
rect 5230 1880 5251 1980
rect 5251 1880 5285 1980
rect 5285 1880 5340 1980
rect 5230 1760 5251 1860
rect 5251 1760 5285 1860
rect 5285 1760 5340 1860
rect 10040 6470 10240 6730
rect 7660 3450 7840 3630
rect 8490 3950 8630 4050
rect 7660 2510 7840 2690
rect 8530 2000 8551 2100
rect 8551 2000 8585 2100
rect 8585 2000 8640 2100
rect 8530 1880 8551 1980
rect 8551 1880 8585 1980
rect 8585 1880 8640 1980
rect 8530 1760 8551 1860
rect 8551 1760 8585 1860
rect 8585 1760 8640 1860
rect 13360 6480 13560 6790
rect 10960 3450 11140 3630
rect 11790 3950 11930 4050
rect 10960 2510 11140 2690
rect 11830 2000 11851 2100
rect 11851 2000 11885 2100
rect 11885 2000 11940 2100
rect 11830 1880 11851 1980
rect 11851 1880 11885 1980
rect 11885 1880 11940 1980
rect 11830 1760 11851 1860
rect 11851 1760 11885 1860
rect 11885 1760 11940 1860
rect 15720 10020 15850 10190
rect 17810 10010 17940 10180
rect 19940 10020 20070 10190
rect 16930 6736 17150 6810
rect 16930 6500 17032 6736
rect 17032 6500 17070 6736
rect 17070 6500 17150 6736
rect 14560 3450 14740 3630
rect 15390 3950 15530 4050
rect 14550 2510 14730 2690
rect 15430 2000 15451 2100
rect 15451 2000 15485 2100
rect 15485 2000 15540 2100
rect 15430 1880 15451 1980
rect 15451 1880 15485 1980
rect 15485 1880 15540 1980
rect 15430 1760 15451 1860
rect 15451 1760 15485 1860
rect 15485 1760 15540 1860
rect 19490 6490 19820 6780
rect 18060 3450 18240 3630
rect 18890 3950 19030 4050
rect 18060 2500 18240 2680
rect 18930 2000 18951 2100
rect 18951 2000 18985 2100
rect 18985 2000 19040 2100
rect 18930 1880 18951 1980
rect 18951 1880 18985 1980
rect 18985 1880 19040 1980
rect 18930 1760 18951 1860
rect 18951 1760 18985 1860
rect 18985 1760 19040 1860
rect 22560 6500 22860 6780
rect 21760 3450 21940 3630
rect 22590 3950 22730 4050
rect 21760 2510 21940 2690
rect 22630 2000 22651 2100
rect 22651 2000 22685 2100
rect 22685 2000 22740 2100
rect 22630 1880 22651 1980
rect 22651 1880 22685 1980
rect 22685 1880 22740 1980
rect 22630 1760 22651 1860
rect 22651 1760 22685 1860
rect 22685 1760 22740 1860
rect 25210 7410 25340 7540
rect 25410 7400 25540 7530
rect 25600 7390 25730 7520
rect 25220 7230 25350 7360
rect 25400 7210 25530 7340
rect 25580 7200 25710 7330
rect 25170 6490 25500 6710
rect 28380 6520 28590 6850
rect 32080 7180 32230 7320
rect 31260 6210 31340 6290
rect 33850 6200 33950 6360
rect 30580 5850 30640 5930
rect 34920 5830 35010 5910
rect 25560 3450 25740 3630
rect 26390 3950 26530 4050
rect 29490 4810 29550 4870
rect 30680 5049 30696 5080
rect 30696 5049 30730 5080
rect 30730 5049 30740 5080
rect 30680 5020 30740 5049
rect 25560 2510 25740 2690
rect 26430 2000 26451 2100
rect 26451 2000 26485 2100
rect 26485 2000 26540 2100
rect 26430 1880 26451 1980
rect 26451 1880 26485 1980
rect 26485 1880 26540 1980
rect 26430 1760 26451 1860
rect 26451 1760 26485 1860
rect 26485 1760 26540 1860
rect 32950 4460 33030 4540
rect 29100 3890 29400 4090
rect 30920 4090 31040 4210
<< metal2 >>
rect 6000 29510 6200 29700
rect 6070 28986 6126 29510
rect 10320 29470 10520 29660
rect 14650 29470 14850 29660
rect 18980 29470 19180 29660
rect 10394 28986 10450 29470
rect 5900 28958 6126 28986
rect 5900 27270 5928 28958
rect 6070 28856 6126 28958
rect 10316 28958 10450 28986
rect 6043 27436 6351 27445
rect 6043 27434 6049 27436
rect 6105 27434 6129 27436
rect 6185 27434 6209 27436
rect 6265 27434 6289 27436
rect 6345 27434 6351 27436
rect 6105 27382 6107 27434
rect 6287 27382 6289 27434
rect 6043 27380 6049 27382
rect 6105 27380 6129 27382
rect 6185 27380 6209 27382
rect 6265 27380 6289 27382
rect 6345 27380 6351 27382
rect 6043 27371 6351 27380
rect 9861 27436 10169 27445
rect 9861 27434 9867 27436
rect 9923 27434 9947 27436
rect 10003 27434 10027 27436
rect 10083 27434 10107 27436
rect 10163 27434 10169 27436
rect 9923 27382 9925 27434
rect 10105 27382 10107 27434
rect 9861 27380 9867 27382
rect 9923 27380 9947 27382
rect 10003 27380 10027 27382
rect 10083 27380 10107 27382
rect 10163 27380 10169 27382
rect 9861 27371 10169 27380
rect 10316 27354 10344 28958
rect 10394 28856 10450 28958
rect 14718 28856 14774 29470
rect 19042 28856 19098 29470
rect 13679 27436 13987 27445
rect 13679 27434 13685 27436
rect 13741 27434 13765 27436
rect 13821 27434 13845 27436
rect 13901 27434 13925 27436
rect 13981 27434 13987 27436
rect 13741 27382 13743 27434
rect 13923 27382 13925 27434
rect 13679 27380 13685 27382
rect 13741 27380 13765 27382
rect 13821 27380 13845 27382
rect 13901 27380 13925 27382
rect 13981 27380 13987 27382
rect 13679 27371 13987 27380
rect 10224 27338 10344 27354
rect 10212 27332 10344 27338
rect 10264 27326 10344 27332
rect 10212 27274 10264 27280
rect 5888 27264 5940 27270
rect 5888 27206 5940 27212
rect 5796 26992 5848 26998
rect 5796 26934 5848 26940
rect 11040 26992 11092 26998
rect 11040 26934 11092 26940
rect 5808 14214 5836 26934
rect 6703 26892 7011 26901
rect 6703 26890 6709 26892
rect 6765 26890 6789 26892
rect 6845 26890 6869 26892
rect 6925 26890 6949 26892
rect 7005 26890 7011 26892
rect 6765 26838 6767 26890
rect 6947 26838 6949 26890
rect 6703 26836 6709 26838
rect 6765 26836 6789 26838
rect 6845 26836 6869 26838
rect 6925 26836 6949 26838
rect 7005 26836 7011 26838
rect 6703 26827 7011 26836
rect 10521 26892 10829 26901
rect 10521 26890 10527 26892
rect 10583 26890 10607 26892
rect 10663 26890 10687 26892
rect 10743 26890 10767 26892
rect 10823 26890 10829 26892
rect 10583 26838 10585 26890
rect 10765 26838 10767 26890
rect 10521 26836 10527 26838
rect 10583 26836 10607 26838
rect 10663 26836 10687 26838
rect 10743 26836 10767 26838
rect 10823 26836 10829 26838
rect 10521 26827 10829 26836
rect 6043 26348 6351 26357
rect 6043 26346 6049 26348
rect 6105 26346 6129 26348
rect 6185 26346 6209 26348
rect 6265 26346 6289 26348
rect 6345 26346 6351 26348
rect 6105 26294 6107 26346
rect 6287 26294 6289 26346
rect 6043 26292 6049 26294
rect 6105 26292 6129 26294
rect 6185 26292 6209 26294
rect 6265 26292 6289 26294
rect 6345 26292 6351 26294
rect 6043 26283 6351 26292
rect 9861 26348 10169 26357
rect 9861 26346 9867 26348
rect 9923 26346 9947 26348
rect 10003 26346 10027 26348
rect 10083 26346 10107 26348
rect 10163 26346 10169 26348
rect 9923 26294 9925 26346
rect 10105 26294 10107 26346
rect 9861 26292 9867 26294
rect 9923 26292 9947 26294
rect 10003 26292 10027 26294
rect 10083 26292 10107 26294
rect 10163 26292 10169 26294
rect 9861 26283 10169 26292
rect 6703 25804 7011 25813
rect 6703 25802 6709 25804
rect 6765 25802 6789 25804
rect 6845 25802 6869 25804
rect 6925 25802 6949 25804
rect 7005 25802 7011 25804
rect 6765 25750 6767 25802
rect 6947 25750 6949 25802
rect 6703 25748 6709 25750
rect 6765 25748 6789 25750
rect 6845 25748 6869 25750
rect 6925 25748 6949 25750
rect 7005 25748 7011 25750
rect 6703 25739 7011 25748
rect 10521 25804 10829 25813
rect 10521 25802 10527 25804
rect 10583 25802 10607 25804
rect 10663 25802 10687 25804
rect 10743 25802 10767 25804
rect 10823 25802 10829 25804
rect 10583 25750 10585 25802
rect 10765 25750 10767 25802
rect 10521 25748 10527 25750
rect 10583 25748 10607 25750
rect 10663 25748 10687 25750
rect 10743 25748 10767 25750
rect 10823 25748 10829 25750
rect 10521 25739 10829 25748
rect 6043 25260 6351 25269
rect 6043 25258 6049 25260
rect 6105 25258 6129 25260
rect 6185 25258 6209 25260
rect 6265 25258 6289 25260
rect 6345 25258 6351 25260
rect 6105 25206 6107 25258
rect 6287 25206 6289 25258
rect 6043 25204 6049 25206
rect 6105 25204 6129 25206
rect 6185 25204 6209 25206
rect 6265 25204 6289 25206
rect 6345 25204 6351 25206
rect 6043 25195 6351 25204
rect 9861 25260 10169 25269
rect 9861 25258 9867 25260
rect 9923 25258 9947 25260
rect 10003 25258 10027 25260
rect 10083 25258 10107 25260
rect 10163 25258 10169 25260
rect 9923 25206 9925 25258
rect 10105 25206 10107 25258
rect 9861 25204 9867 25206
rect 9923 25204 9947 25206
rect 10003 25204 10027 25206
rect 10083 25204 10107 25206
rect 10163 25204 10169 25206
rect 9861 25195 10169 25204
rect 6703 24716 7011 24725
rect 6703 24714 6709 24716
rect 6765 24714 6789 24716
rect 6845 24714 6869 24716
rect 6925 24714 6949 24716
rect 7005 24714 7011 24716
rect 6765 24662 6767 24714
rect 6947 24662 6949 24714
rect 6703 24660 6709 24662
rect 6765 24660 6789 24662
rect 6845 24660 6869 24662
rect 6925 24660 6949 24662
rect 7005 24660 7011 24662
rect 6703 24651 7011 24660
rect 10521 24716 10829 24725
rect 10521 24714 10527 24716
rect 10583 24714 10607 24716
rect 10663 24714 10687 24716
rect 10743 24714 10767 24716
rect 10823 24714 10829 24716
rect 10583 24662 10585 24714
rect 10765 24662 10767 24714
rect 10521 24660 10527 24662
rect 10583 24660 10607 24662
rect 10663 24660 10687 24662
rect 10743 24660 10767 24662
rect 10823 24660 10829 24662
rect 10521 24651 10829 24660
rect 6043 24172 6351 24181
rect 6043 24170 6049 24172
rect 6105 24170 6129 24172
rect 6185 24170 6209 24172
rect 6265 24170 6289 24172
rect 6345 24170 6351 24172
rect 6105 24118 6107 24170
rect 6287 24118 6289 24170
rect 6043 24116 6049 24118
rect 6105 24116 6129 24118
rect 6185 24116 6209 24118
rect 6265 24116 6289 24118
rect 6345 24116 6351 24118
rect 6043 24107 6351 24116
rect 9861 24172 10169 24181
rect 9861 24170 9867 24172
rect 9923 24170 9947 24172
rect 10003 24170 10027 24172
rect 10083 24170 10107 24172
rect 10163 24170 10169 24172
rect 9923 24118 9925 24170
rect 10105 24118 10107 24170
rect 9861 24116 9867 24118
rect 9923 24116 9947 24118
rect 10003 24116 10027 24118
rect 10083 24116 10107 24118
rect 10163 24116 10169 24118
rect 9861 24107 10169 24116
rect 6703 23628 7011 23637
rect 6703 23626 6709 23628
rect 6765 23626 6789 23628
rect 6845 23626 6869 23628
rect 6925 23626 6949 23628
rect 7005 23626 7011 23628
rect 6765 23574 6767 23626
rect 6947 23574 6949 23626
rect 6703 23572 6709 23574
rect 6765 23572 6789 23574
rect 6845 23572 6869 23574
rect 6925 23572 6949 23574
rect 7005 23572 7011 23574
rect 6703 23563 7011 23572
rect 10521 23628 10829 23637
rect 10521 23626 10527 23628
rect 10583 23626 10607 23628
rect 10663 23626 10687 23628
rect 10743 23626 10767 23628
rect 10823 23626 10829 23628
rect 10583 23574 10585 23626
rect 10765 23574 10767 23626
rect 10521 23572 10527 23574
rect 10583 23572 10607 23574
rect 10663 23572 10687 23574
rect 10743 23572 10767 23574
rect 10823 23572 10829 23574
rect 10521 23563 10829 23572
rect 6043 23084 6351 23093
rect 6043 23082 6049 23084
rect 6105 23082 6129 23084
rect 6185 23082 6209 23084
rect 6265 23082 6289 23084
rect 6345 23082 6351 23084
rect 6105 23030 6107 23082
rect 6287 23030 6289 23082
rect 6043 23028 6049 23030
rect 6105 23028 6129 23030
rect 6185 23028 6209 23030
rect 6265 23028 6289 23030
rect 6345 23028 6351 23030
rect 6043 23019 6351 23028
rect 9861 23084 10169 23093
rect 9861 23082 9867 23084
rect 9923 23082 9947 23084
rect 10003 23082 10027 23084
rect 10083 23082 10107 23084
rect 10163 23082 10169 23084
rect 9923 23030 9925 23082
rect 10105 23030 10107 23082
rect 9861 23028 9867 23030
rect 9923 23028 9947 23030
rect 10003 23028 10027 23030
rect 10083 23028 10107 23030
rect 10163 23028 10169 23030
rect 9861 23019 10169 23028
rect 6703 22540 7011 22549
rect 6703 22538 6709 22540
rect 6765 22538 6789 22540
rect 6845 22538 6869 22540
rect 6925 22538 6949 22540
rect 7005 22538 7011 22540
rect 6765 22486 6767 22538
rect 6947 22486 6949 22538
rect 6703 22484 6709 22486
rect 6765 22484 6789 22486
rect 6845 22484 6869 22486
rect 6925 22484 6949 22486
rect 7005 22484 7011 22486
rect 6703 22475 7011 22484
rect 10521 22540 10829 22549
rect 10521 22538 10527 22540
rect 10583 22538 10607 22540
rect 10663 22538 10687 22540
rect 10743 22538 10767 22540
rect 10823 22538 10829 22540
rect 10583 22486 10585 22538
rect 10765 22486 10767 22538
rect 10521 22484 10527 22486
rect 10583 22484 10607 22486
rect 10663 22484 10687 22486
rect 10743 22484 10767 22486
rect 10823 22484 10829 22486
rect 10521 22475 10829 22484
rect 6043 21996 6351 22005
rect 6043 21994 6049 21996
rect 6105 21994 6129 21996
rect 6185 21994 6209 21996
rect 6265 21994 6289 21996
rect 6345 21994 6351 21996
rect 6105 21942 6107 21994
rect 6287 21942 6289 21994
rect 6043 21940 6049 21942
rect 6105 21940 6129 21942
rect 6185 21940 6209 21942
rect 6265 21940 6289 21942
rect 6345 21940 6351 21942
rect 6043 21931 6351 21940
rect 9861 21996 10169 22005
rect 9861 21994 9867 21996
rect 9923 21994 9947 21996
rect 10003 21994 10027 21996
rect 10083 21994 10107 21996
rect 10163 21994 10169 21996
rect 9923 21942 9925 21994
rect 10105 21942 10107 21994
rect 9861 21940 9867 21942
rect 9923 21940 9947 21942
rect 10003 21940 10027 21942
rect 10083 21940 10107 21942
rect 10163 21940 10169 21942
rect 9861 21931 10169 21940
rect 6703 21452 7011 21461
rect 6703 21450 6709 21452
rect 6765 21450 6789 21452
rect 6845 21450 6869 21452
rect 6925 21450 6949 21452
rect 7005 21450 7011 21452
rect 6765 21398 6767 21450
rect 6947 21398 6949 21450
rect 6703 21396 6709 21398
rect 6765 21396 6789 21398
rect 6845 21396 6869 21398
rect 6925 21396 6949 21398
rect 7005 21396 7011 21398
rect 6703 21387 7011 21396
rect 10521 21452 10829 21461
rect 10521 21450 10527 21452
rect 10583 21450 10607 21452
rect 10663 21450 10687 21452
rect 10743 21450 10767 21452
rect 10823 21450 10829 21452
rect 10583 21398 10585 21450
rect 10765 21398 10767 21450
rect 10521 21396 10527 21398
rect 10583 21396 10607 21398
rect 10663 21396 10687 21398
rect 10743 21396 10767 21398
rect 10823 21396 10829 21398
rect 10521 21387 10829 21396
rect 6043 20908 6351 20917
rect 6043 20906 6049 20908
rect 6105 20906 6129 20908
rect 6185 20906 6209 20908
rect 6265 20906 6289 20908
rect 6345 20906 6351 20908
rect 6105 20854 6107 20906
rect 6287 20854 6289 20906
rect 6043 20852 6049 20854
rect 6105 20852 6129 20854
rect 6185 20852 6209 20854
rect 6265 20852 6289 20854
rect 6345 20852 6351 20854
rect 6043 20843 6351 20852
rect 9861 20908 10169 20917
rect 9861 20906 9867 20908
rect 9923 20906 9947 20908
rect 10003 20906 10027 20908
rect 10083 20906 10107 20908
rect 10163 20906 10169 20908
rect 9923 20854 9925 20906
rect 10105 20854 10107 20906
rect 9861 20852 9867 20854
rect 9923 20852 9947 20854
rect 10003 20852 10027 20854
rect 10083 20852 10107 20854
rect 10163 20852 10169 20854
rect 9861 20843 10169 20852
rect 6703 20364 7011 20373
rect 6703 20362 6709 20364
rect 6765 20362 6789 20364
rect 6845 20362 6869 20364
rect 6925 20362 6949 20364
rect 7005 20362 7011 20364
rect 6765 20310 6767 20362
rect 6947 20310 6949 20362
rect 6703 20308 6709 20310
rect 6765 20308 6789 20310
rect 6845 20308 6869 20310
rect 6925 20308 6949 20310
rect 7005 20308 7011 20310
rect 6703 20299 7011 20308
rect 10521 20364 10829 20373
rect 10521 20362 10527 20364
rect 10583 20362 10607 20364
rect 10663 20362 10687 20364
rect 10743 20362 10767 20364
rect 10823 20362 10829 20364
rect 10583 20310 10585 20362
rect 10765 20310 10767 20362
rect 10521 20308 10527 20310
rect 10583 20308 10607 20310
rect 10663 20308 10687 20310
rect 10743 20308 10767 20310
rect 10823 20308 10829 20310
rect 10521 20299 10829 20308
rect 6043 19820 6351 19829
rect 6043 19818 6049 19820
rect 6105 19818 6129 19820
rect 6185 19818 6209 19820
rect 6265 19818 6289 19820
rect 6345 19818 6351 19820
rect 6105 19766 6107 19818
rect 6287 19766 6289 19818
rect 6043 19764 6049 19766
rect 6105 19764 6129 19766
rect 6185 19764 6209 19766
rect 6265 19764 6289 19766
rect 6345 19764 6351 19766
rect 6043 19755 6351 19764
rect 9861 19820 10169 19829
rect 9861 19818 9867 19820
rect 9923 19818 9947 19820
rect 10003 19818 10027 19820
rect 10083 19818 10107 19820
rect 10163 19818 10169 19820
rect 9923 19766 9925 19818
rect 10105 19766 10107 19818
rect 9861 19764 9867 19766
rect 9923 19764 9947 19766
rect 10003 19764 10027 19766
rect 10083 19764 10107 19766
rect 10163 19764 10169 19766
rect 9861 19755 10169 19764
rect 6703 19276 7011 19285
rect 6703 19274 6709 19276
rect 6765 19274 6789 19276
rect 6845 19274 6869 19276
rect 6925 19274 6949 19276
rect 7005 19274 7011 19276
rect 6765 19222 6767 19274
rect 6947 19222 6949 19274
rect 6703 19220 6709 19222
rect 6765 19220 6789 19222
rect 6845 19220 6869 19222
rect 6925 19220 6949 19222
rect 7005 19220 7011 19222
rect 6703 19211 7011 19220
rect 10521 19276 10829 19285
rect 10521 19274 10527 19276
rect 10583 19274 10607 19276
rect 10663 19274 10687 19276
rect 10743 19274 10767 19276
rect 10823 19274 10829 19276
rect 10583 19222 10585 19274
rect 10765 19222 10767 19274
rect 10521 19220 10527 19222
rect 10583 19220 10607 19222
rect 10663 19220 10687 19222
rect 10743 19220 10767 19222
rect 10823 19220 10829 19222
rect 10521 19211 10829 19220
rect 6043 18732 6351 18741
rect 6043 18730 6049 18732
rect 6105 18730 6129 18732
rect 6185 18730 6209 18732
rect 6265 18730 6289 18732
rect 6345 18730 6351 18732
rect 6105 18678 6107 18730
rect 6287 18678 6289 18730
rect 6043 18676 6049 18678
rect 6105 18676 6129 18678
rect 6185 18676 6209 18678
rect 6265 18676 6289 18678
rect 6345 18676 6351 18678
rect 6043 18667 6351 18676
rect 9861 18732 10169 18741
rect 9861 18730 9867 18732
rect 9923 18730 9947 18732
rect 10003 18730 10027 18732
rect 10083 18730 10107 18732
rect 10163 18730 10169 18732
rect 9923 18678 9925 18730
rect 10105 18678 10107 18730
rect 9861 18676 9867 18678
rect 9923 18676 9947 18678
rect 10003 18676 10027 18678
rect 10083 18676 10107 18678
rect 10163 18676 10169 18678
rect 9861 18667 10169 18676
rect 6703 18188 7011 18197
rect 6703 18186 6709 18188
rect 6765 18186 6789 18188
rect 6845 18186 6869 18188
rect 6925 18186 6949 18188
rect 7005 18186 7011 18188
rect 6765 18134 6767 18186
rect 6947 18134 6949 18186
rect 6703 18132 6709 18134
rect 6765 18132 6789 18134
rect 6845 18132 6869 18134
rect 6925 18132 6949 18134
rect 7005 18132 7011 18134
rect 6703 18123 7011 18132
rect 10521 18188 10829 18197
rect 10521 18186 10527 18188
rect 10583 18186 10607 18188
rect 10663 18186 10687 18188
rect 10743 18186 10767 18188
rect 10823 18186 10829 18188
rect 10583 18134 10585 18186
rect 10765 18134 10767 18186
rect 10521 18132 10527 18134
rect 10583 18132 10607 18134
rect 10663 18132 10687 18134
rect 10743 18132 10767 18134
rect 10823 18132 10829 18134
rect 10521 18123 10829 18132
rect 6043 17644 6351 17653
rect 6043 17642 6049 17644
rect 6105 17642 6129 17644
rect 6185 17642 6209 17644
rect 6265 17642 6289 17644
rect 6345 17642 6351 17644
rect 6105 17590 6107 17642
rect 6287 17590 6289 17642
rect 6043 17588 6049 17590
rect 6105 17588 6129 17590
rect 6185 17588 6209 17590
rect 6265 17588 6289 17590
rect 6345 17588 6351 17590
rect 6043 17579 6351 17588
rect 9861 17644 10169 17653
rect 9861 17642 9867 17644
rect 9923 17642 9947 17644
rect 10003 17642 10027 17644
rect 10083 17642 10107 17644
rect 10163 17642 10169 17644
rect 9923 17590 9925 17642
rect 10105 17590 10107 17642
rect 9861 17588 9867 17590
rect 9923 17588 9947 17590
rect 10003 17588 10027 17590
rect 10083 17588 10107 17590
rect 10163 17588 10169 17590
rect 9861 17579 10169 17588
rect 6703 17100 7011 17109
rect 6703 17098 6709 17100
rect 6765 17098 6789 17100
rect 6845 17098 6869 17100
rect 6925 17098 6949 17100
rect 7005 17098 7011 17100
rect 6765 17046 6767 17098
rect 6947 17046 6949 17098
rect 6703 17044 6709 17046
rect 6765 17044 6789 17046
rect 6845 17044 6869 17046
rect 6925 17044 6949 17046
rect 7005 17044 7011 17046
rect 6703 17035 7011 17044
rect 10521 17100 10829 17109
rect 10521 17098 10527 17100
rect 10583 17098 10607 17100
rect 10663 17098 10687 17100
rect 10743 17098 10767 17100
rect 10823 17098 10829 17100
rect 10583 17046 10585 17098
rect 10765 17046 10767 17098
rect 10521 17044 10527 17046
rect 10583 17044 10607 17046
rect 10663 17044 10687 17046
rect 10743 17044 10767 17046
rect 10823 17044 10829 17046
rect 10521 17035 10829 17044
rect 6043 16556 6351 16565
rect 6043 16554 6049 16556
rect 6105 16554 6129 16556
rect 6185 16554 6209 16556
rect 6265 16554 6289 16556
rect 6345 16554 6351 16556
rect 6105 16502 6107 16554
rect 6287 16502 6289 16554
rect 6043 16500 6049 16502
rect 6105 16500 6129 16502
rect 6185 16500 6209 16502
rect 6265 16500 6289 16502
rect 6345 16500 6351 16502
rect 6043 16491 6351 16500
rect 9861 16556 10169 16565
rect 9861 16554 9867 16556
rect 9923 16554 9947 16556
rect 10003 16554 10027 16556
rect 10083 16554 10107 16556
rect 10163 16554 10169 16556
rect 9923 16502 9925 16554
rect 10105 16502 10107 16554
rect 9861 16500 9867 16502
rect 9923 16500 9947 16502
rect 10003 16500 10027 16502
rect 10083 16500 10107 16502
rect 10163 16500 10169 16502
rect 9861 16491 10169 16500
rect 6703 16012 7011 16021
rect 6703 16010 6709 16012
rect 6765 16010 6789 16012
rect 6845 16010 6869 16012
rect 6925 16010 6949 16012
rect 7005 16010 7011 16012
rect 6765 15958 6767 16010
rect 6947 15958 6949 16010
rect 6703 15956 6709 15958
rect 6765 15956 6789 15958
rect 6845 15956 6869 15958
rect 6925 15956 6949 15958
rect 7005 15956 7011 15958
rect 6703 15947 7011 15956
rect 10521 16012 10829 16021
rect 10521 16010 10527 16012
rect 10583 16010 10607 16012
rect 10663 16010 10687 16012
rect 10743 16010 10767 16012
rect 10823 16010 10829 16012
rect 10583 15958 10585 16010
rect 10765 15958 10767 16010
rect 10521 15956 10527 15958
rect 10583 15956 10607 15958
rect 10663 15956 10687 15958
rect 10743 15956 10767 15958
rect 10823 15956 10829 15958
rect 10521 15947 10829 15956
rect 6043 15468 6351 15477
rect 6043 15466 6049 15468
rect 6105 15466 6129 15468
rect 6185 15466 6209 15468
rect 6265 15466 6289 15468
rect 6345 15466 6351 15468
rect 6105 15414 6107 15466
rect 6287 15414 6289 15466
rect 6043 15412 6049 15414
rect 6105 15412 6129 15414
rect 6185 15412 6209 15414
rect 6265 15412 6289 15414
rect 6345 15412 6351 15414
rect 6043 15403 6351 15412
rect 9861 15468 10169 15477
rect 9861 15466 9867 15468
rect 9923 15466 9947 15468
rect 10003 15466 10027 15468
rect 10083 15466 10107 15468
rect 10163 15466 10169 15468
rect 9923 15414 9925 15466
rect 10105 15414 10107 15466
rect 9861 15412 9867 15414
rect 9923 15412 9947 15414
rect 10003 15412 10027 15414
rect 10083 15412 10107 15414
rect 10163 15412 10169 15414
rect 9861 15403 10169 15412
rect 6703 14924 7011 14933
rect 6703 14922 6709 14924
rect 6765 14922 6789 14924
rect 6845 14922 6869 14924
rect 6925 14922 6949 14924
rect 7005 14922 7011 14924
rect 6765 14870 6767 14922
rect 6947 14870 6949 14922
rect 6703 14868 6709 14870
rect 6765 14868 6789 14870
rect 6845 14868 6869 14870
rect 6925 14868 6949 14870
rect 7005 14868 7011 14870
rect 6703 14859 7011 14868
rect 10521 14924 10829 14933
rect 10521 14922 10527 14924
rect 10583 14922 10607 14924
rect 10663 14922 10687 14924
rect 10743 14922 10767 14924
rect 10823 14922 10829 14924
rect 10583 14870 10585 14922
rect 10765 14870 10767 14922
rect 10521 14868 10527 14870
rect 10583 14868 10607 14870
rect 10663 14868 10687 14870
rect 10743 14868 10767 14870
rect 10823 14868 10829 14870
rect 10521 14859 10829 14868
rect 11052 14622 11080 26934
rect 14339 26892 14647 26901
rect 14339 26890 14345 26892
rect 14401 26890 14425 26892
rect 14481 26890 14505 26892
rect 14561 26890 14585 26892
rect 14641 26890 14647 26892
rect 14401 26838 14403 26890
rect 14583 26838 14585 26890
rect 14339 26836 14345 26838
rect 14401 26836 14425 26838
rect 14481 26836 14505 26838
rect 14561 26836 14585 26838
rect 14641 26836 14647 26838
rect 14339 26827 14647 26836
rect 13679 26348 13987 26357
rect 13679 26346 13685 26348
rect 13741 26346 13765 26348
rect 13821 26346 13845 26348
rect 13901 26346 13925 26348
rect 13981 26346 13987 26348
rect 13741 26294 13743 26346
rect 13923 26294 13925 26346
rect 13679 26292 13685 26294
rect 13741 26292 13765 26294
rect 13821 26292 13845 26294
rect 13901 26292 13925 26294
rect 13981 26292 13987 26294
rect 13679 26283 13987 26292
rect 14339 25804 14647 25813
rect 14339 25802 14345 25804
rect 14401 25802 14425 25804
rect 14481 25802 14505 25804
rect 14561 25802 14585 25804
rect 14641 25802 14647 25804
rect 14401 25750 14403 25802
rect 14583 25750 14585 25802
rect 14339 25748 14345 25750
rect 14401 25748 14425 25750
rect 14481 25748 14505 25750
rect 14561 25748 14585 25750
rect 14641 25748 14647 25750
rect 14339 25739 14647 25748
rect 14732 25366 14760 28856
rect 17497 27436 17805 27445
rect 17497 27434 17503 27436
rect 17559 27434 17583 27436
rect 17639 27434 17663 27436
rect 17719 27434 17743 27436
rect 17799 27434 17805 27436
rect 17559 27382 17561 27434
rect 17741 27382 17743 27434
rect 17497 27380 17503 27382
rect 17559 27380 17583 27382
rect 17639 27380 17663 27382
rect 17719 27380 17743 27382
rect 17799 27380 17805 27382
rect 17497 27371 17805 27380
rect 19056 27270 19084 28856
rect 19044 27264 19096 27270
rect 19044 27206 19096 27212
rect 18768 26992 18820 26998
rect 18768 26934 18820 26940
rect 18157 26892 18465 26901
rect 18157 26890 18163 26892
rect 18219 26890 18243 26892
rect 18299 26890 18323 26892
rect 18379 26890 18403 26892
rect 18459 26890 18465 26892
rect 18219 26838 18221 26890
rect 18401 26838 18403 26890
rect 18157 26836 18163 26838
rect 18219 26836 18243 26838
rect 18299 26836 18323 26838
rect 18379 26836 18403 26838
rect 18459 26836 18465 26838
rect 18157 26827 18465 26836
rect 17497 26348 17805 26357
rect 17497 26346 17503 26348
rect 17559 26346 17583 26348
rect 17639 26346 17663 26348
rect 17719 26346 17743 26348
rect 17799 26346 17805 26348
rect 17559 26294 17561 26346
rect 17741 26294 17743 26346
rect 17497 26292 17503 26294
rect 17559 26292 17583 26294
rect 17639 26292 17663 26294
rect 17719 26292 17743 26294
rect 17799 26292 17805 26294
rect 17497 26283 17805 26292
rect 18157 25804 18465 25813
rect 18157 25802 18163 25804
rect 18219 25802 18243 25804
rect 18299 25802 18323 25804
rect 18379 25802 18403 25804
rect 18459 25802 18465 25804
rect 18219 25750 18221 25802
rect 18401 25750 18403 25802
rect 18157 25748 18163 25750
rect 18219 25748 18243 25750
rect 18299 25748 18323 25750
rect 18379 25748 18403 25750
rect 18459 25748 18465 25750
rect 18157 25739 18465 25748
rect 14076 25360 14128 25366
rect 14076 25302 14128 25308
rect 14720 25360 14772 25366
rect 14720 25302 14772 25308
rect 13679 25260 13987 25269
rect 13679 25258 13685 25260
rect 13741 25258 13765 25260
rect 13821 25258 13845 25260
rect 13901 25258 13925 25260
rect 13981 25258 13987 25260
rect 13741 25206 13743 25258
rect 13923 25206 13925 25258
rect 13679 25204 13685 25206
rect 13741 25204 13765 25206
rect 13821 25204 13845 25206
rect 13901 25204 13925 25206
rect 13981 25204 13987 25206
rect 13679 25195 13987 25204
rect 13679 24172 13987 24181
rect 13679 24170 13685 24172
rect 13741 24170 13765 24172
rect 13821 24170 13845 24172
rect 13901 24170 13925 24172
rect 13981 24170 13987 24172
rect 13741 24118 13743 24170
rect 13923 24118 13925 24170
rect 13679 24116 13685 24118
rect 13741 24116 13765 24118
rect 13821 24116 13845 24118
rect 13901 24116 13925 24118
rect 13981 24116 13987 24118
rect 13679 24107 13987 24116
rect 13679 23084 13987 23093
rect 13679 23082 13685 23084
rect 13741 23082 13765 23084
rect 13821 23082 13845 23084
rect 13901 23082 13925 23084
rect 13981 23082 13987 23084
rect 13741 23030 13743 23082
rect 13923 23030 13925 23082
rect 13679 23028 13685 23030
rect 13741 23028 13765 23030
rect 13821 23028 13845 23030
rect 13901 23028 13925 23030
rect 13981 23028 13987 23030
rect 13679 23019 13987 23028
rect 13679 21996 13987 22005
rect 13679 21994 13685 21996
rect 13741 21994 13765 21996
rect 13821 21994 13845 21996
rect 13901 21994 13925 21996
rect 13981 21994 13987 21996
rect 13741 21942 13743 21994
rect 13923 21942 13925 21994
rect 13679 21940 13685 21942
rect 13741 21940 13765 21942
rect 13821 21940 13845 21942
rect 13901 21940 13925 21942
rect 13981 21940 13987 21942
rect 13679 21931 13987 21940
rect 13679 20908 13987 20917
rect 13679 20906 13685 20908
rect 13741 20906 13765 20908
rect 13821 20906 13845 20908
rect 13901 20906 13925 20908
rect 13981 20906 13987 20908
rect 13741 20854 13743 20906
rect 13923 20854 13925 20906
rect 13679 20852 13685 20854
rect 13741 20852 13765 20854
rect 13821 20852 13845 20854
rect 13901 20852 13925 20854
rect 13981 20852 13987 20854
rect 13679 20843 13987 20852
rect 13679 19820 13987 19829
rect 13679 19818 13685 19820
rect 13741 19818 13765 19820
rect 13821 19818 13845 19820
rect 13901 19818 13925 19820
rect 13981 19818 13987 19820
rect 13741 19766 13743 19818
rect 13923 19766 13925 19818
rect 13679 19764 13685 19766
rect 13741 19764 13765 19766
rect 13821 19764 13845 19766
rect 13901 19764 13925 19766
rect 13981 19764 13987 19766
rect 13679 19755 13987 19764
rect 13679 18732 13987 18741
rect 13679 18730 13685 18732
rect 13741 18730 13765 18732
rect 13821 18730 13845 18732
rect 13901 18730 13925 18732
rect 13981 18730 13987 18732
rect 13741 18678 13743 18730
rect 13923 18678 13925 18730
rect 13679 18676 13685 18678
rect 13741 18676 13765 18678
rect 13821 18676 13845 18678
rect 13901 18676 13925 18678
rect 13981 18676 13987 18678
rect 13679 18667 13987 18676
rect 13679 17644 13987 17653
rect 13679 17642 13685 17644
rect 13741 17642 13765 17644
rect 13821 17642 13845 17644
rect 13901 17642 13925 17644
rect 13981 17642 13987 17644
rect 13741 17590 13743 17642
rect 13923 17590 13925 17642
rect 13679 17588 13685 17590
rect 13741 17588 13765 17590
rect 13821 17588 13845 17590
rect 13901 17588 13925 17590
rect 13981 17588 13987 17590
rect 13679 17579 13987 17588
rect 13679 16556 13987 16565
rect 13679 16554 13685 16556
rect 13741 16554 13765 16556
rect 13821 16554 13845 16556
rect 13901 16554 13925 16556
rect 13981 16554 13987 16556
rect 13741 16502 13743 16554
rect 13923 16502 13925 16554
rect 13679 16500 13685 16502
rect 13741 16500 13765 16502
rect 13821 16500 13845 16502
rect 13901 16500 13925 16502
rect 13981 16500 13987 16502
rect 13679 16491 13987 16500
rect 13679 15468 13987 15477
rect 13679 15466 13685 15468
rect 13741 15466 13765 15468
rect 13821 15466 13845 15468
rect 13901 15466 13925 15468
rect 13981 15466 13987 15468
rect 13741 15414 13743 15466
rect 13923 15414 13925 15466
rect 13679 15412 13685 15414
rect 13741 15412 13765 15414
rect 13821 15412 13845 15414
rect 13901 15412 13925 15414
rect 13981 15412 13987 15414
rect 13679 15403 13987 15412
rect 12880 15160 12932 15166
rect 12880 15102 12932 15108
rect 11684 14684 11736 14690
rect 11684 14626 11736 14632
rect 11040 14616 11092 14622
rect 11040 14558 11092 14564
rect 10212 14480 10264 14486
rect 10212 14422 10264 14428
rect 11408 14480 11460 14486
rect 11408 14422 11460 14428
rect 6043 14380 6351 14389
rect 6043 14378 6049 14380
rect 6105 14378 6129 14380
rect 6185 14378 6209 14380
rect 6265 14378 6289 14380
rect 6345 14378 6351 14380
rect 6105 14326 6107 14378
rect 6287 14326 6289 14378
rect 6043 14324 6049 14326
rect 6105 14324 6129 14326
rect 6185 14324 6209 14326
rect 6265 14324 6289 14326
rect 6345 14324 6351 14326
rect 6043 14315 6351 14324
rect 9861 14380 10169 14389
rect 9861 14378 9867 14380
rect 9923 14378 9947 14380
rect 10003 14378 10027 14380
rect 10083 14378 10107 14380
rect 10163 14378 10169 14380
rect 9923 14326 9925 14378
rect 10105 14326 10107 14378
rect 9861 14324 9867 14326
rect 9923 14324 9947 14326
rect 10003 14324 10027 14326
rect 10083 14324 10107 14326
rect 10163 14324 10169 14326
rect 9861 14315 10169 14324
rect 5796 14208 5848 14214
rect 5796 14150 5848 14156
rect 10224 13942 10252 14422
rect 11420 14282 11448 14422
rect 11408 14276 11460 14282
rect 11408 14218 11460 14224
rect 10856 14072 10908 14078
rect 10856 14014 10908 14020
rect 10212 13936 10264 13942
rect 10212 13878 10264 13884
rect 6703 13836 7011 13845
rect 6703 13834 6709 13836
rect 6765 13834 6789 13836
rect 6845 13834 6869 13836
rect 6925 13834 6949 13836
rect 7005 13834 7011 13836
rect 6765 13782 6767 13834
rect 6947 13782 6949 13834
rect 6703 13780 6709 13782
rect 6765 13780 6789 13782
rect 6845 13780 6869 13782
rect 6925 13780 6949 13782
rect 7005 13780 7011 13782
rect 6703 13771 7011 13780
rect 9660 13528 9712 13534
rect 9660 13470 9712 13476
rect 6043 13292 6351 13301
rect 6043 13290 6049 13292
rect 6105 13290 6129 13292
rect 6185 13290 6209 13292
rect 6265 13290 6289 13292
rect 6345 13290 6351 13292
rect 6105 13238 6107 13290
rect 6287 13238 6289 13290
rect 6043 13236 6049 13238
rect 6105 13236 6129 13238
rect 6185 13236 6209 13238
rect 6265 13236 6289 13238
rect 6345 13236 6351 13238
rect 6043 13227 6351 13236
rect 9200 12984 9252 12990
rect 9200 12926 9252 12932
rect 6703 12748 7011 12757
rect 6703 12746 6709 12748
rect 6765 12746 6789 12748
rect 6845 12746 6869 12748
rect 6925 12746 6949 12748
rect 7005 12746 7011 12748
rect 6765 12694 6767 12746
rect 6947 12694 6949 12746
rect 6703 12692 6709 12694
rect 6765 12692 6789 12694
rect 6845 12692 6869 12694
rect 6925 12692 6949 12694
rect 7005 12692 7011 12694
rect 6703 12683 7011 12692
rect 9212 12446 9240 12926
rect 9672 12650 9700 13470
rect 9861 13292 10169 13301
rect 9861 13290 9867 13292
rect 9923 13290 9947 13292
rect 10003 13290 10027 13292
rect 10083 13290 10107 13292
rect 10163 13290 10169 13292
rect 9923 13238 9925 13290
rect 10105 13238 10107 13290
rect 9861 13236 9867 13238
rect 9923 13236 9947 13238
rect 10003 13236 10027 13238
rect 10083 13236 10107 13238
rect 10163 13236 10169 13238
rect 9861 13227 10169 13236
rect 10224 13176 10252 13878
rect 10521 13836 10829 13845
rect 10521 13834 10527 13836
rect 10583 13834 10607 13836
rect 10663 13834 10687 13836
rect 10743 13834 10767 13836
rect 10823 13834 10829 13836
rect 10583 13782 10585 13834
rect 10765 13782 10767 13834
rect 10521 13780 10527 13782
rect 10583 13780 10607 13782
rect 10663 13780 10687 13782
rect 10743 13780 10767 13782
rect 10823 13780 10829 13782
rect 10521 13771 10829 13780
rect 10868 13534 10896 14014
rect 10856 13528 10908 13534
rect 10856 13470 10908 13476
rect 10580 13392 10632 13398
rect 10580 13334 10632 13340
rect 10592 13194 10620 13334
rect 10132 13148 10252 13176
rect 10580 13188 10632 13194
rect 9752 12848 9804 12854
rect 9752 12790 9804 12796
rect 9660 12644 9712 12650
rect 9660 12586 9712 12592
rect 9764 12514 9792 12790
rect 9752 12508 9804 12514
rect 9752 12450 9804 12456
rect 10132 12446 10160 13148
rect 10580 13130 10632 13136
rect 10868 13126 10896 13470
rect 10856 13120 10908 13126
rect 10856 13062 10908 13068
rect 10212 12848 10264 12854
rect 10212 12790 10264 12796
rect 11500 12848 11552 12854
rect 11500 12790 11552 12796
rect 10224 12650 10252 12790
rect 10521 12748 10829 12757
rect 10521 12746 10527 12748
rect 10583 12746 10607 12748
rect 10663 12746 10687 12748
rect 10743 12746 10767 12748
rect 10823 12746 10829 12748
rect 10583 12694 10585 12746
rect 10765 12694 10767 12746
rect 10521 12692 10527 12694
rect 10583 12692 10607 12694
rect 10663 12692 10687 12694
rect 10743 12692 10767 12694
rect 10823 12692 10829 12694
rect 10521 12683 10829 12692
rect 10212 12644 10264 12650
rect 10212 12586 10264 12592
rect 5244 12440 5296 12446
rect 5244 12382 5296 12388
rect 9200 12440 9252 12446
rect 9200 12382 9252 12388
rect 10120 12440 10172 12446
rect 10120 12382 10172 12388
rect 5256 11306 5284 12382
rect 7268 12304 7320 12310
rect 7268 12246 7320 12252
rect 9384 12304 9436 12310
rect 9384 12246 9436 12252
rect 6043 12204 6351 12213
rect 6043 12202 6049 12204
rect 6105 12202 6129 12204
rect 6185 12202 6209 12204
rect 6265 12202 6289 12204
rect 6345 12202 6351 12204
rect 6105 12150 6107 12202
rect 6287 12150 6289 12202
rect 6043 12148 6049 12150
rect 6105 12148 6129 12150
rect 6185 12148 6209 12150
rect 6265 12148 6289 12150
rect 6345 12148 6351 12150
rect 6043 12139 6351 12148
rect 5164 11278 5284 11306
rect 5164 10800 5192 11278
rect 7280 10800 7308 12246
rect 9396 10800 9424 12246
rect 9861 12204 10169 12213
rect 9861 12202 9867 12204
rect 9923 12202 9947 12204
rect 10003 12202 10027 12204
rect 10083 12202 10107 12204
rect 10163 12202 10169 12204
rect 9923 12150 9925 12202
rect 10105 12150 10107 12202
rect 9861 12148 9867 12150
rect 9923 12148 9947 12150
rect 10003 12148 10027 12150
rect 10083 12148 10107 12150
rect 10163 12148 10169 12150
rect 9861 12139 10169 12148
rect 11512 10800 11540 12790
rect 11696 12514 11724 14626
rect 11868 14072 11920 14078
rect 11868 14014 11920 14020
rect 11880 13738 11908 14014
rect 12696 13936 12748 13942
rect 12696 13878 12748 13884
rect 12708 13738 12736 13878
rect 11868 13732 11920 13738
rect 11868 13674 11920 13680
rect 12696 13732 12748 13738
rect 12696 13674 12748 13680
rect 11880 13194 11908 13674
rect 12696 13528 12748 13534
rect 12696 13470 12748 13476
rect 12512 13392 12564 13398
rect 12512 13334 12564 13340
rect 11868 13188 11920 13194
rect 11868 13130 11920 13136
rect 12524 12990 12552 13334
rect 12512 12984 12564 12990
rect 12512 12926 12564 12932
rect 12708 12650 12736 13470
rect 12892 12854 12920 15102
rect 13432 15024 13484 15030
rect 13432 14966 13484 14972
rect 13444 14826 13472 14966
rect 13432 14820 13484 14826
rect 13432 14762 13484 14768
rect 13064 14480 13116 14486
rect 13064 14422 13116 14428
rect 13432 14480 13484 14486
rect 13432 14422 13484 14428
rect 13076 13738 13104 14422
rect 13064 13732 13116 13738
rect 13064 13674 13116 13680
rect 13076 12990 13104 13674
rect 13064 12984 13116 12990
rect 13064 12926 13116 12932
rect 12880 12848 12932 12854
rect 12880 12790 12932 12796
rect 12696 12644 12748 12650
rect 12696 12586 12748 12592
rect 11684 12508 11736 12514
rect 11684 12450 11736 12456
rect 12892 12310 12920 12790
rect 13076 12530 13104 12926
rect 13076 12502 13196 12530
rect 13168 12446 13196 12502
rect 13444 12446 13472 14422
rect 13679 14380 13987 14389
rect 13679 14378 13685 14380
rect 13741 14378 13765 14380
rect 13821 14378 13845 14380
rect 13901 14378 13925 14380
rect 13981 14378 13987 14380
rect 13741 14326 13743 14378
rect 13923 14326 13925 14378
rect 13679 14324 13685 14326
rect 13741 14324 13765 14326
rect 13821 14324 13845 14326
rect 13901 14324 13925 14326
rect 13981 14324 13987 14326
rect 13679 14315 13987 14324
rect 13984 14208 14036 14214
rect 14088 14162 14116 25302
rect 17497 25260 17805 25269
rect 17497 25258 17503 25260
rect 17559 25258 17583 25260
rect 17639 25258 17663 25260
rect 17719 25258 17743 25260
rect 17799 25258 17805 25260
rect 17559 25206 17561 25258
rect 17741 25206 17743 25258
rect 17497 25204 17503 25206
rect 17559 25204 17583 25206
rect 17639 25204 17663 25206
rect 17719 25204 17743 25206
rect 17799 25204 17805 25206
rect 17497 25195 17805 25204
rect 14339 24716 14647 24725
rect 14339 24714 14345 24716
rect 14401 24714 14425 24716
rect 14481 24714 14505 24716
rect 14561 24714 14585 24716
rect 14641 24714 14647 24716
rect 14401 24662 14403 24714
rect 14583 24662 14585 24714
rect 14339 24660 14345 24662
rect 14401 24660 14425 24662
rect 14481 24660 14505 24662
rect 14561 24660 14585 24662
rect 14641 24660 14647 24662
rect 14339 24651 14647 24660
rect 18157 24716 18465 24725
rect 18157 24714 18163 24716
rect 18219 24714 18243 24716
rect 18299 24714 18323 24716
rect 18379 24714 18403 24716
rect 18459 24714 18465 24716
rect 18219 24662 18221 24714
rect 18401 24662 18403 24714
rect 18157 24660 18163 24662
rect 18219 24660 18243 24662
rect 18299 24660 18323 24662
rect 18379 24660 18403 24662
rect 18459 24660 18465 24662
rect 18157 24651 18465 24660
rect 17497 24172 17805 24181
rect 17497 24170 17503 24172
rect 17559 24170 17583 24172
rect 17639 24170 17663 24172
rect 17719 24170 17743 24172
rect 17799 24170 17805 24172
rect 17559 24118 17561 24170
rect 17741 24118 17743 24170
rect 17497 24116 17503 24118
rect 17559 24116 17583 24118
rect 17639 24116 17663 24118
rect 17719 24116 17743 24118
rect 17799 24116 17805 24118
rect 17497 24107 17805 24116
rect 14339 23628 14647 23637
rect 14339 23626 14345 23628
rect 14401 23626 14425 23628
rect 14481 23626 14505 23628
rect 14561 23626 14585 23628
rect 14641 23626 14647 23628
rect 14401 23574 14403 23626
rect 14583 23574 14585 23626
rect 14339 23572 14345 23574
rect 14401 23572 14425 23574
rect 14481 23572 14505 23574
rect 14561 23572 14585 23574
rect 14641 23572 14647 23574
rect 14339 23563 14647 23572
rect 18157 23628 18465 23637
rect 18157 23626 18163 23628
rect 18219 23626 18243 23628
rect 18299 23626 18323 23628
rect 18379 23626 18403 23628
rect 18459 23626 18465 23628
rect 18219 23574 18221 23626
rect 18401 23574 18403 23626
rect 18157 23572 18163 23574
rect 18219 23572 18243 23574
rect 18299 23572 18323 23574
rect 18379 23572 18403 23574
rect 18459 23572 18465 23574
rect 18157 23563 18465 23572
rect 17497 23084 17805 23093
rect 17497 23082 17503 23084
rect 17559 23082 17583 23084
rect 17639 23082 17663 23084
rect 17719 23082 17743 23084
rect 17799 23082 17805 23084
rect 17559 23030 17561 23082
rect 17741 23030 17743 23082
rect 17497 23028 17503 23030
rect 17559 23028 17583 23030
rect 17639 23028 17663 23030
rect 17719 23028 17743 23030
rect 17799 23028 17805 23030
rect 17497 23019 17805 23028
rect 14339 22540 14647 22549
rect 14339 22538 14345 22540
rect 14401 22538 14425 22540
rect 14481 22538 14505 22540
rect 14561 22538 14585 22540
rect 14641 22538 14647 22540
rect 14401 22486 14403 22538
rect 14583 22486 14585 22538
rect 14339 22484 14345 22486
rect 14401 22484 14425 22486
rect 14481 22484 14505 22486
rect 14561 22484 14585 22486
rect 14641 22484 14647 22486
rect 14339 22475 14647 22484
rect 18157 22540 18465 22549
rect 18157 22538 18163 22540
rect 18219 22538 18243 22540
rect 18299 22538 18323 22540
rect 18379 22538 18403 22540
rect 18459 22538 18465 22540
rect 18219 22486 18221 22538
rect 18401 22486 18403 22538
rect 18157 22484 18163 22486
rect 18219 22484 18243 22486
rect 18299 22484 18323 22486
rect 18379 22484 18403 22486
rect 18459 22484 18465 22486
rect 18157 22475 18465 22484
rect 17497 21996 17805 22005
rect 17497 21994 17503 21996
rect 17559 21994 17583 21996
rect 17639 21994 17663 21996
rect 17719 21994 17743 21996
rect 17799 21994 17805 21996
rect 17559 21942 17561 21994
rect 17741 21942 17743 21994
rect 17497 21940 17503 21942
rect 17559 21940 17583 21942
rect 17639 21940 17663 21942
rect 17719 21940 17743 21942
rect 17799 21940 17805 21942
rect 17497 21931 17805 21940
rect 14339 21452 14647 21461
rect 14339 21450 14345 21452
rect 14401 21450 14425 21452
rect 14481 21450 14505 21452
rect 14561 21450 14585 21452
rect 14641 21450 14647 21452
rect 14401 21398 14403 21450
rect 14583 21398 14585 21450
rect 14339 21396 14345 21398
rect 14401 21396 14425 21398
rect 14481 21396 14505 21398
rect 14561 21396 14585 21398
rect 14641 21396 14647 21398
rect 14339 21387 14647 21396
rect 18157 21452 18465 21461
rect 18157 21450 18163 21452
rect 18219 21450 18243 21452
rect 18299 21450 18323 21452
rect 18379 21450 18403 21452
rect 18459 21450 18465 21452
rect 18219 21398 18221 21450
rect 18401 21398 18403 21450
rect 18157 21396 18163 21398
rect 18219 21396 18243 21398
rect 18299 21396 18323 21398
rect 18379 21396 18403 21398
rect 18459 21396 18465 21398
rect 18157 21387 18465 21396
rect 17497 20908 17805 20917
rect 17497 20906 17503 20908
rect 17559 20906 17583 20908
rect 17639 20906 17663 20908
rect 17719 20906 17743 20908
rect 17799 20906 17805 20908
rect 17559 20854 17561 20906
rect 17741 20854 17743 20906
rect 17497 20852 17503 20854
rect 17559 20852 17583 20854
rect 17639 20852 17663 20854
rect 17719 20852 17743 20854
rect 17799 20852 17805 20854
rect 17497 20843 17805 20852
rect 14339 20364 14647 20373
rect 14339 20362 14345 20364
rect 14401 20362 14425 20364
rect 14481 20362 14505 20364
rect 14561 20362 14585 20364
rect 14641 20362 14647 20364
rect 14401 20310 14403 20362
rect 14583 20310 14585 20362
rect 14339 20308 14345 20310
rect 14401 20308 14425 20310
rect 14481 20308 14505 20310
rect 14561 20308 14585 20310
rect 14641 20308 14647 20310
rect 14339 20299 14647 20308
rect 18157 20364 18465 20373
rect 18157 20362 18163 20364
rect 18219 20362 18243 20364
rect 18299 20362 18323 20364
rect 18379 20362 18403 20364
rect 18459 20362 18465 20364
rect 18219 20310 18221 20362
rect 18401 20310 18403 20362
rect 18157 20308 18163 20310
rect 18219 20308 18243 20310
rect 18299 20308 18323 20310
rect 18379 20308 18403 20310
rect 18459 20308 18465 20310
rect 18157 20299 18465 20308
rect 17497 19820 17805 19829
rect 17497 19818 17503 19820
rect 17559 19818 17583 19820
rect 17639 19818 17663 19820
rect 17719 19818 17743 19820
rect 17799 19818 17805 19820
rect 17559 19766 17561 19818
rect 17741 19766 17743 19818
rect 17497 19764 17503 19766
rect 17559 19764 17583 19766
rect 17639 19764 17663 19766
rect 17719 19764 17743 19766
rect 17799 19764 17805 19766
rect 17497 19755 17805 19764
rect 14339 19276 14647 19285
rect 14339 19274 14345 19276
rect 14401 19274 14425 19276
rect 14481 19274 14505 19276
rect 14561 19274 14585 19276
rect 14641 19274 14647 19276
rect 14401 19222 14403 19274
rect 14583 19222 14585 19274
rect 14339 19220 14345 19222
rect 14401 19220 14425 19222
rect 14481 19220 14505 19222
rect 14561 19220 14585 19222
rect 14641 19220 14647 19222
rect 14339 19211 14647 19220
rect 18157 19276 18465 19285
rect 18157 19274 18163 19276
rect 18219 19274 18243 19276
rect 18299 19274 18323 19276
rect 18379 19274 18403 19276
rect 18459 19274 18465 19276
rect 18219 19222 18221 19274
rect 18401 19222 18403 19274
rect 18157 19220 18163 19222
rect 18219 19220 18243 19222
rect 18299 19220 18323 19222
rect 18379 19220 18403 19222
rect 18459 19220 18465 19222
rect 18157 19211 18465 19220
rect 17497 18732 17805 18741
rect 17497 18730 17503 18732
rect 17559 18730 17583 18732
rect 17639 18730 17663 18732
rect 17719 18730 17743 18732
rect 17799 18730 17805 18732
rect 17559 18678 17561 18730
rect 17741 18678 17743 18730
rect 17497 18676 17503 18678
rect 17559 18676 17583 18678
rect 17639 18676 17663 18678
rect 17719 18676 17743 18678
rect 17799 18676 17805 18678
rect 17497 18667 17805 18676
rect 14339 18188 14647 18197
rect 14339 18186 14345 18188
rect 14401 18186 14425 18188
rect 14481 18186 14505 18188
rect 14561 18186 14585 18188
rect 14641 18186 14647 18188
rect 14401 18134 14403 18186
rect 14583 18134 14585 18186
rect 14339 18132 14345 18134
rect 14401 18132 14425 18134
rect 14481 18132 14505 18134
rect 14561 18132 14585 18134
rect 14641 18132 14647 18134
rect 14339 18123 14647 18132
rect 18157 18188 18465 18197
rect 18157 18186 18163 18188
rect 18219 18186 18243 18188
rect 18299 18186 18323 18188
rect 18379 18186 18403 18188
rect 18459 18186 18465 18188
rect 18219 18134 18221 18186
rect 18401 18134 18403 18186
rect 18157 18132 18163 18134
rect 18219 18132 18243 18134
rect 18299 18132 18323 18134
rect 18379 18132 18403 18134
rect 18459 18132 18465 18134
rect 18157 18123 18465 18132
rect 17497 17644 17805 17653
rect 17497 17642 17503 17644
rect 17559 17642 17583 17644
rect 17639 17642 17663 17644
rect 17719 17642 17743 17644
rect 17799 17642 17805 17644
rect 17559 17590 17561 17642
rect 17741 17590 17743 17642
rect 17497 17588 17503 17590
rect 17559 17588 17583 17590
rect 17639 17588 17663 17590
rect 17719 17588 17743 17590
rect 17799 17588 17805 17590
rect 17497 17579 17805 17588
rect 14339 17100 14647 17109
rect 14339 17098 14345 17100
rect 14401 17098 14425 17100
rect 14481 17098 14505 17100
rect 14561 17098 14585 17100
rect 14641 17098 14647 17100
rect 14401 17046 14403 17098
rect 14583 17046 14585 17098
rect 14339 17044 14345 17046
rect 14401 17044 14425 17046
rect 14481 17044 14505 17046
rect 14561 17044 14585 17046
rect 14641 17044 14647 17046
rect 14339 17035 14647 17044
rect 18157 17100 18465 17109
rect 18157 17098 18163 17100
rect 18219 17098 18243 17100
rect 18299 17098 18323 17100
rect 18379 17098 18403 17100
rect 18459 17098 18465 17100
rect 18219 17046 18221 17098
rect 18401 17046 18403 17098
rect 18157 17044 18163 17046
rect 18219 17044 18243 17046
rect 18299 17044 18323 17046
rect 18379 17044 18403 17046
rect 18459 17044 18465 17046
rect 18157 17035 18465 17044
rect 17497 16556 17805 16565
rect 17497 16554 17503 16556
rect 17559 16554 17583 16556
rect 17639 16554 17663 16556
rect 17719 16554 17743 16556
rect 17799 16554 17805 16556
rect 17559 16502 17561 16554
rect 17741 16502 17743 16554
rect 17497 16500 17503 16502
rect 17559 16500 17583 16502
rect 17639 16500 17663 16502
rect 17719 16500 17743 16502
rect 17799 16500 17805 16502
rect 17497 16491 17805 16500
rect 14339 16012 14647 16021
rect 14339 16010 14345 16012
rect 14401 16010 14425 16012
rect 14481 16010 14505 16012
rect 14561 16010 14585 16012
rect 14641 16010 14647 16012
rect 14401 15958 14403 16010
rect 14583 15958 14585 16010
rect 14339 15956 14345 15958
rect 14401 15956 14425 15958
rect 14481 15956 14505 15958
rect 14561 15956 14585 15958
rect 14641 15956 14647 15958
rect 14339 15947 14647 15956
rect 18157 16012 18465 16021
rect 18157 16010 18163 16012
rect 18219 16010 18243 16012
rect 18299 16010 18323 16012
rect 18379 16010 18403 16012
rect 18459 16010 18465 16012
rect 18219 15958 18221 16010
rect 18401 15958 18403 16010
rect 18157 15956 18163 15958
rect 18219 15956 18243 15958
rect 18299 15956 18323 15958
rect 18379 15956 18403 15958
rect 18459 15956 18465 15958
rect 18157 15947 18465 15956
rect 17497 15468 17805 15477
rect 17497 15466 17503 15468
rect 17559 15466 17583 15468
rect 17639 15466 17663 15468
rect 17719 15466 17743 15468
rect 17799 15466 17805 15468
rect 17559 15414 17561 15466
rect 17741 15414 17743 15466
rect 17497 15412 17503 15414
rect 17559 15412 17583 15414
rect 17639 15412 17663 15414
rect 17719 15412 17743 15414
rect 17799 15412 17805 15414
rect 17497 15403 17805 15412
rect 15364 15160 15416 15166
rect 15364 15102 15416 15108
rect 14339 14924 14647 14933
rect 14339 14922 14345 14924
rect 14401 14922 14425 14924
rect 14481 14922 14505 14924
rect 14561 14922 14585 14924
rect 14641 14922 14647 14924
rect 14401 14870 14403 14922
rect 14583 14870 14585 14922
rect 14339 14868 14345 14870
rect 14401 14868 14425 14870
rect 14481 14868 14505 14870
rect 14561 14868 14585 14870
rect 14641 14868 14647 14870
rect 14339 14859 14647 14868
rect 14996 14752 15048 14758
rect 14996 14694 15048 14700
rect 14260 14616 14312 14622
rect 14260 14558 14312 14564
rect 14036 14156 14116 14162
rect 13984 14150 14116 14156
rect 13996 14134 14116 14150
rect 14168 14072 14220 14078
rect 14168 14014 14220 14020
rect 14076 13460 14128 13466
rect 14076 13402 14128 13408
rect 13679 13292 13987 13301
rect 13679 13290 13685 13292
rect 13741 13290 13765 13292
rect 13821 13290 13845 13292
rect 13901 13290 13925 13292
rect 13981 13290 13987 13292
rect 13741 13238 13743 13290
rect 13923 13238 13925 13290
rect 13679 13236 13685 13238
rect 13741 13236 13765 13238
rect 13821 13236 13845 13238
rect 13901 13236 13925 13238
rect 13981 13236 13987 13238
rect 13679 13227 13987 13236
rect 14088 12650 14116 13402
rect 14180 12854 14208 14014
rect 14272 12922 14300 14558
rect 14352 14480 14404 14486
rect 14352 14422 14404 14428
rect 14364 14078 14392 14422
rect 14352 14072 14404 14078
rect 14352 14014 14404 14020
rect 14812 14072 14864 14078
rect 14812 14014 14864 14020
rect 14720 13936 14772 13942
rect 14720 13878 14772 13884
rect 14339 13836 14647 13845
rect 14339 13834 14345 13836
rect 14401 13834 14425 13836
rect 14481 13834 14505 13836
rect 14561 13834 14585 13836
rect 14641 13834 14647 13836
rect 14401 13782 14403 13834
rect 14583 13782 14585 13834
rect 14339 13780 14345 13782
rect 14401 13780 14425 13782
rect 14481 13780 14505 13782
rect 14561 13780 14585 13782
rect 14641 13780 14647 13782
rect 14339 13771 14647 13780
rect 14732 13534 14760 13878
rect 14720 13528 14772 13534
rect 14720 13470 14772 13476
rect 14444 13392 14496 13398
rect 14444 13334 14496 13340
rect 14456 13194 14484 13334
rect 14444 13188 14496 13194
rect 14444 13130 14496 13136
rect 14824 13126 14852 14014
rect 15008 13126 15036 14694
rect 15376 14282 15404 15102
rect 16100 15024 16152 15030
rect 16100 14966 16152 14972
rect 15548 14548 15600 14554
rect 15548 14490 15600 14496
rect 16008 14548 16060 14554
rect 16008 14490 16060 14496
rect 15364 14276 15416 14282
rect 15364 14218 15416 14224
rect 15088 13596 15140 13602
rect 15088 13538 15140 13544
rect 14720 13120 14772 13126
rect 14720 13062 14772 13068
rect 14812 13120 14864 13126
rect 14812 13062 14864 13068
rect 14996 13120 15048 13126
rect 14996 13062 15048 13068
rect 14260 12916 14312 12922
rect 14260 12858 14312 12864
rect 14168 12848 14220 12854
rect 14168 12790 14220 12796
rect 14076 12644 14128 12650
rect 14076 12586 14128 12592
rect 14180 12514 14208 12790
rect 14339 12748 14647 12757
rect 14339 12746 14345 12748
rect 14401 12746 14425 12748
rect 14481 12746 14505 12748
rect 14561 12746 14585 12748
rect 14641 12746 14647 12748
rect 14401 12694 14403 12746
rect 14583 12694 14585 12746
rect 14339 12692 14345 12694
rect 14401 12692 14425 12694
rect 14481 12692 14505 12694
rect 14561 12692 14585 12694
rect 14641 12692 14647 12694
rect 14339 12683 14647 12692
rect 14732 12650 14760 13062
rect 14720 12644 14772 12650
rect 14720 12586 14772 12592
rect 15100 12514 15128 13538
rect 15560 13058 15588 14490
rect 15640 14480 15692 14486
rect 15640 14422 15692 14428
rect 15652 14282 15680 14422
rect 16020 14282 16048 14490
rect 16112 14282 16140 14966
rect 18157 14924 18465 14933
rect 18157 14922 18163 14924
rect 18219 14922 18243 14924
rect 18299 14922 18323 14924
rect 18379 14922 18403 14924
rect 18459 14922 18465 14924
rect 18219 14870 18221 14922
rect 18401 14870 18403 14922
rect 18157 14868 18163 14870
rect 18219 14868 18243 14870
rect 18299 14868 18323 14870
rect 18379 14868 18403 14870
rect 18459 14868 18465 14870
rect 18157 14859 18465 14868
rect 16284 14616 16336 14622
rect 16284 14558 16336 14564
rect 15640 14276 15692 14282
rect 15640 14218 15692 14224
rect 16008 14276 16060 14282
rect 16008 14218 16060 14224
rect 16100 14276 16152 14282
rect 16100 14218 16152 14224
rect 15652 13534 15680 14218
rect 15732 13936 15784 13942
rect 15732 13878 15784 13884
rect 15640 13528 15692 13534
rect 15640 13470 15692 13476
rect 15548 13052 15600 13058
rect 15548 12994 15600 13000
rect 14168 12508 14220 12514
rect 14168 12450 14220 12456
rect 15088 12508 15140 12514
rect 15088 12450 15140 12456
rect 13156 12440 13208 12446
rect 13156 12382 13208 12388
rect 13432 12440 13484 12446
rect 13432 12382 13484 12388
rect 15560 12310 15588 12994
rect 15744 12514 15772 13878
rect 16296 13738 16324 14558
rect 17497 14380 17805 14389
rect 17497 14378 17503 14380
rect 17559 14378 17583 14380
rect 17639 14378 17663 14380
rect 17719 14378 17743 14380
rect 17799 14378 17805 14380
rect 17559 14326 17561 14378
rect 17741 14326 17743 14378
rect 17497 14324 17503 14326
rect 17559 14324 17583 14326
rect 17639 14324 17663 14326
rect 17719 14324 17743 14326
rect 17799 14324 17805 14326
rect 17497 14315 17805 14324
rect 16468 14140 16520 14146
rect 16468 14082 16520 14088
rect 16480 13738 16508 14082
rect 17112 13936 17164 13942
rect 17112 13878 17164 13884
rect 16284 13732 16336 13738
rect 16284 13674 16336 13680
rect 16468 13732 16520 13738
rect 16468 13674 16520 13680
rect 16296 13194 16324 13674
rect 17124 13602 17152 13878
rect 18157 13836 18465 13845
rect 18157 13834 18163 13836
rect 18219 13834 18243 13836
rect 18299 13834 18323 13836
rect 18379 13834 18403 13836
rect 18459 13834 18465 13836
rect 18219 13782 18221 13834
rect 18401 13782 18403 13834
rect 18157 13780 18163 13782
rect 18219 13780 18243 13782
rect 18299 13780 18323 13782
rect 18379 13780 18403 13782
rect 18459 13780 18465 13782
rect 18157 13771 18465 13780
rect 18780 13602 18808 26934
rect 17112 13596 17164 13602
rect 17112 13538 17164 13544
rect 18768 13596 18820 13602
rect 18768 13538 18820 13544
rect 16928 13528 16980 13534
rect 16928 13470 16980 13476
rect 16284 13188 16336 13194
rect 16284 13130 16336 13136
rect 15732 12508 15784 12514
rect 15732 12450 15784 12456
rect 16940 12446 16968 13470
rect 17020 13392 17072 13398
rect 17020 13334 17072 13340
rect 17032 13194 17060 13334
rect 17497 13292 17805 13301
rect 17497 13290 17503 13292
rect 17559 13290 17583 13292
rect 17639 13290 17663 13292
rect 17719 13290 17743 13292
rect 17799 13290 17805 13292
rect 17559 13238 17561 13290
rect 17741 13238 17743 13290
rect 17497 13236 17503 13238
rect 17559 13236 17583 13238
rect 17639 13236 17663 13238
rect 17719 13236 17743 13238
rect 17799 13236 17805 13238
rect 17497 13227 17805 13236
rect 17020 13188 17072 13194
rect 17020 13130 17072 13136
rect 17572 12984 17624 12990
rect 17572 12926 17624 12932
rect 17584 12446 17612 12926
rect 18157 12748 18465 12757
rect 18157 12746 18163 12748
rect 18219 12746 18243 12748
rect 18299 12746 18323 12748
rect 18379 12746 18403 12748
rect 18459 12746 18465 12748
rect 18219 12694 18221 12746
rect 18401 12694 18403 12746
rect 18157 12692 18163 12694
rect 18219 12692 18243 12694
rect 18299 12692 18323 12694
rect 18379 12692 18403 12694
rect 18459 12692 18465 12694
rect 18157 12683 18465 12692
rect 16928 12440 16980 12446
rect 16928 12382 16980 12388
rect 17572 12440 17624 12446
rect 17572 12382 17624 12388
rect 15640 12372 15692 12378
rect 15640 12314 15692 12320
rect 17848 12372 17900 12378
rect 17848 12314 17900 12320
rect 19964 12372 20016 12378
rect 19964 12314 20016 12320
rect 12880 12304 12932 12310
rect 13616 12304 13668 12310
rect 12880 12246 12932 12252
rect 13536 12252 13616 12258
rect 13536 12246 13668 12252
rect 15548 12304 15600 12310
rect 15548 12246 15600 12252
rect 13536 12230 13656 12246
rect 13536 11170 13564 12230
rect 13679 12204 13987 12213
rect 13679 12202 13685 12204
rect 13741 12202 13765 12204
rect 13821 12202 13845 12204
rect 13901 12202 13925 12204
rect 13981 12202 13987 12204
rect 13741 12150 13743 12202
rect 13923 12150 13925 12202
rect 13679 12148 13685 12150
rect 13741 12148 13765 12150
rect 13821 12148 13845 12150
rect 13901 12148 13925 12150
rect 13981 12148 13987 12150
rect 13679 12139 13987 12148
rect 15652 11170 15680 12314
rect 17497 12204 17805 12213
rect 17497 12202 17503 12204
rect 17559 12202 17583 12204
rect 17639 12202 17663 12204
rect 17719 12202 17743 12204
rect 17799 12202 17805 12204
rect 17559 12150 17561 12202
rect 17741 12150 17743 12202
rect 17497 12148 17503 12150
rect 17559 12148 17583 12150
rect 17639 12148 17663 12150
rect 17719 12148 17743 12150
rect 17799 12148 17805 12150
rect 17497 12139 17805 12148
rect 13536 11142 13656 11170
rect 15652 11142 15772 11170
rect 13628 10800 13656 11142
rect 15744 10800 15772 11142
rect 17860 10800 17888 12314
rect 19976 10800 20004 12314
rect 5150 10180 5206 10800
rect 5140 10160 5260 10180
rect 7266 10160 7322 10800
rect 9382 10200 9438 10800
rect 11498 10200 11554 10800
rect 13614 10200 13670 10800
rect 15730 10200 15786 10800
rect 9340 10190 9470 10200
rect 5140 10020 5160 10160
rect 5140 10010 5260 10020
rect 7240 10150 7370 10160
rect 5150 10000 5206 10010
rect 9340 10010 9470 10020
rect 11430 10190 11560 10200
rect 11430 10010 11560 10020
rect 13600 10190 13730 10200
rect 13600 10010 13730 10020
rect 15720 10190 15850 10200
rect 17846 10190 17902 10800
rect 19962 10200 20018 10800
rect 19940 10190 20070 10200
rect 15720 10010 15850 10020
rect 17810 10180 17940 10190
rect 19940 10010 20070 10020
rect 9382 10000 9438 10010
rect 11498 10000 11554 10010
rect 13614 10000 13670 10010
rect 15730 10000 15786 10010
rect 17810 10000 17940 10010
rect 19962 10000 20018 10010
rect 7240 9970 7370 9980
rect 28530 7780 35010 8200
rect 28530 7570 28950 7780
rect 25190 7540 28950 7570
rect 25190 7410 25210 7540
rect 25340 7530 28950 7540
rect 25340 7410 25410 7530
rect 25190 7400 25410 7410
rect 25540 7520 28950 7530
rect 25540 7400 25600 7520
rect 25190 7390 25600 7400
rect 25730 7390 28950 7520
rect 25190 7360 28950 7390
rect 25190 7230 25220 7360
rect 25350 7340 28950 7360
rect 25350 7230 25400 7340
rect 25190 7210 25400 7230
rect 25530 7330 28950 7340
rect 25530 7210 25580 7330
rect 25190 7200 25580 7210
rect 25710 7200 28950 7330
rect 25190 7180 28950 7200
rect 32060 7330 32260 7340
rect 32060 7190 32070 7330
rect 32220 7320 32260 7330
rect 32060 7180 32080 7190
rect 32230 7180 32260 7320
rect 25190 7150 28900 7180
rect 32060 7150 32260 7180
rect 3400 6850 28610 6880
rect 3400 6810 28380 6850
rect 3400 6790 16930 6810
rect 3400 6730 13360 6790
rect 3400 6720 10040 6730
rect 3400 6480 3430 6720
rect 3650 6610 10040 6720
rect 3650 6490 6730 6610
rect 6940 6490 10040 6610
rect 3650 6480 10040 6490
rect 3400 6470 10040 6480
rect 10240 6480 13360 6730
rect 13560 6500 16930 6790
rect 17150 6780 28380 6810
rect 17150 6500 19490 6780
rect 13560 6490 19490 6500
rect 19820 6500 22560 6780
rect 22860 6710 28380 6780
rect 22860 6500 25170 6710
rect 19820 6490 25170 6500
rect 25500 6520 28380 6710
rect 28590 6520 28610 6850
rect 25500 6490 28610 6520
rect 13560 6480 28610 6490
rect 10240 6470 28610 6480
rect 3400 6460 28610 6470
rect 33830 6360 33960 6380
rect 31240 6290 31360 6310
rect 31240 6210 31260 6290
rect 31340 6210 31360 6290
rect 31240 6190 31360 6210
rect 33830 6200 33850 6360
rect 33950 6200 33960 6360
rect 33830 6190 33960 6200
rect 31260 5950 31340 6190
rect 30560 5930 31340 5950
rect 33840 5930 33950 6190
rect 34930 5930 35010 7780
rect 30560 5850 30580 5930
rect 30640 5870 31340 5930
rect 32935 5910 35015 5930
rect 30640 5850 30660 5870
rect 30560 5830 30660 5850
rect 32935 5830 34920 5910
rect 35010 5830 35015 5910
rect 32935 5820 35015 5830
rect 30670 5080 30750 5090
rect 30670 5020 30680 5080
rect 30740 5020 30750 5080
rect 30670 5010 30750 5020
rect 29480 4870 29560 4880
rect 30690 4870 30740 5010
rect 29480 4810 29490 4870
rect 29550 4820 30740 4870
rect 29550 4810 29560 4820
rect 29480 4800 29560 4810
rect 32935 4540 33045 5820
rect 32935 4460 32950 4540
rect 33030 4460 33045 4540
rect 32935 4415 33045 4460
rect 30900 4210 31050 4220
rect 29100 4090 29400 4100
rect 1870 4050 2050 4060
rect 1870 3950 1890 4050
rect 2030 3950 2050 4050
rect 1870 3940 2050 3950
rect 5170 4050 5350 4060
rect 5170 3950 5190 4050
rect 5330 3950 5350 4050
rect 5170 3940 5350 3950
rect 8470 4050 8650 4060
rect 8470 3950 8490 4050
rect 8630 3950 8650 4050
rect 8470 3940 8650 3950
rect 11770 4050 11950 4060
rect 11770 3950 11790 4050
rect 11930 3950 11950 4050
rect 11770 3940 11950 3950
rect 15370 4050 15550 4060
rect 15370 3950 15390 4050
rect 15530 3950 15550 4050
rect 15370 3940 15550 3950
rect 18870 4050 19050 4060
rect 18870 3950 18890 4050
rect 19030 3950 19050 4050
rect 18870 3940 19050 3950
rect 22570 4050 22750 4060
rect 22570 3950 22590 4050
rect 22730 3950 22750 4050
rect 22570 3940 22750 3950
rect 26370 4050 26550 4060
rect 26370 3950 26390 4050
rect 26530 3950 26550 4050
rect 26370 3940 26550 3950
rect 420 3630 620 3640
rect 420 3450 430 3630
rect 610 3450 620 3630
rect 420 3440 620 3450
rect 1040 3620 1240 3630
rect 1040 3440 1050 3620
rect 1230 3440 1240 3620
rect 1040 3430 1240 3440
rect 430 2690 650 2700
rect 430 2510 440 2690
rect 620 2510 650 2690
rect 430 2500 650 2510
rect 1050 2690 1250 2700
rect 1050 2510 1060 2690
rect 1240 2510 1250 2690
rect 1050 2500 1250 2510
rect 1920 2120 2000 3940
rect 4350 3630 4550 3640
rect 4350 3450 4360 3630
rect 4540 3450 4550 3630
rect 4350 3440 4550 3450
rect 4340 2690 4540 2700
rect 4340 2510 4350 2690
rect 4530 2510 4540 2690
rect 4340 2500 4540 2510
rect 5220 2120 5300 3940
rect 7650 3630 7850 3640
rect 7650 3450 7660 3630
rect 7840 3450 7850 3630
rect 7650 3440 7850 3450
rect 7650 2690 7850 2700
rect 7650 2510 7660 2690
rect 7840 2510 7850 2690
rect 7650 2500 7850 2510
rect 8520 2120 8600 3940
rect 10950 3630 11150 3640
rect 10950 3450 10960 3630
rect 11140 3450 11150 3630
rect 10950 3440 11150 3450
rect 10950 2690 11150 2700
rect 10950 2510 10960 2690
rect 11140 2510 11150 2690
rect 10950 2500 11150 2510
rect 11820 2120 11900 3940
rect 14550 3630 14750 3640
rect 14550 3450 14560 3630
rect 14740 3450 14750 3630
rect 14550 3440 14750 3450
rect 14540 2690 14740 2700
rect 14540 2510 14550 2690
rect 14730 2510 14740 2690
rect 14540 2500 14740 2510
rect 15420 2120 15500 3940
rect 18050 3630 18250 3640
rect 18050 3450 18060 3630
rect 18240 3450 18250 3630
rect 18050 3440 18250 3450
rect 18050 2680 18250 2690
rect 18050 2500 18060 2680
rect 18240 2500 18250 2680
rect 18050 2490 18250 2500
rect 18920 2120 19000 3940
rect 21750 3630 21950 3640
rect 21750 3450 21760 3630
rect 21940 3450 21950 3630
rect 21750 3440 21950 3450
rect 21750 2690 21950 2700
rect 21750 2510 21760 2690
rect 21940 2510 21950 2690
rect 21750 2500 21950 2510
rect 22620 2120 22700 3940
rect 25550 3630 25750 3640
rect 25550 3450 25560 3630
rect 25740 3450 25750 3630
rect 25550 3440 25750 3450
rect 25550 2690 25750 2700
rect 25550 2510 25560 2690
rect 25740 2510 25750 2690
rect 25550 2500 25750 2510
rect 26420 2120 26500 3940
rect 30900 4090 30920 4210
rect 31040 4090 31050 4210
rect 32940 4200 33040 4415
rect 32940 4100 32950 4200
rect 33030 4100 33040 4200
rect 32940 4090 33040 4100
rect 30900 4080 31050 4090
rect 29100 3880 29400 3890
rect 1920 2100 2050 2120
rect 1920 2000 1930 2100
rect 2040 2000 2050 2100
rect 1920 1980 2050 2000
rect 1920 1880 1930 1980
rect 2040 1880 2050 1980
rect 1920 1860 2050 1880
rect 1920 1760 1930 1860
rect 2040 1760 2050 1860
rect 1920 1730 2050 1760
rect 5220 2100 5350 2120
rect 5220 2000 5230 2100
rect 5340 2000 5350 2100
rect 5220 1980 5350 2000
rect 5220 1880 5230 1980
rect 5340 1880 5350 1980
rect 5220 1860 5350 1880
rect 5220 1760 5230 1860
rect 5340 1760 5350 1860
rect 5220 1730 5350 1760
rect 8520 2100 8650 2120
rect 8520 2000 8530 2100
rect 8640 2000 8650 2100
rect 8520 1980 8650 2000
rect 8520 1880 8530 1980
rect 8640 1880 8650 1980
rect 8520 1860 8650 1880
rect 8520 1760 8530 1860
rect 8640 1760 8650 1860
rect 8520 1730 8650 1760
rect 11820 2100 11950 2120
rect 11820 2000 11830 2100
rect 11940 2000 11950 2100
rect 11820 1980 11950 2000
rect 11820 1880 11830 1980
rect 11940 1880 11950 1980
rect 11820 1860 11950 1880
rect 11820 1760 11830 1860
rect 11940 1760 11950 1860
rect 11820 1730 11950 1760
rect 15420 2100 15550 2120
rect 15420 2000 15430 2100
rect 15540 2000 15550 2100
rect 15420 1980 15550 2000
rect 15420 1880 15430 1980
rect 15540 1880 15550 1980
rect 15420 1860 15550 1880
rect 15420 1760 15430 1860
rect 15540 1760 15550 1860
rect 15420 1730 15550 1760
rect 18920 2100 19050 2120
rect 18920 2000 18930 2100
rect 19040 2000 19050 2100
rect 18920 1980 19050 2000
rect 18920 1880 18930 1980
rect 19040 1880 19050 1980
rect 18920 1860 19050 1880
rect 18920 1760 18930 1860
rect 19040 1760 19050 1860
rect 18920 1730 19050 1760
rect 22620 2100 22750 2120
rect 22620 2000 22630 2100
rect 22740 2000 22750 2100
rect 22620 1980 22750 2000
rect 22620 1880 22630 1980
rect 22740 1880 22750 1980
rect 22620 1860 22750 1880
rect 22620 1760 22630 1860
rect 22740 1760 22750 1860
rect 22620 1730 22750 1760
rect 26420 2100 26550 2120
rect 26420 2000 26430 2100
rect 26540 2000 26550 2100
rect 26420 1980 26550 2000
rect 26420 1880 26430 1980
rect 26540 1880 26550 1980
rect 26420 1860 26550 1880
rect 26420 1760 26430 1860
rect 26540 1760 26550 1860
rect 26420 1730 26550 1760
<< via2 >>
rect 6049 27434 6105 27436
rect 6129 27434 6185 27436
rect 6209 27434 6265 27436
rect 6289 27434 6345 27436
rect 6049 27382 6095 27434
rect 6095 27382 6105 27434
rect 6129 27382 6159 27434
rect 6159 27382 6171 27434
rect 6171 27382 6185 27434
rect 6209 27382 6223 27434
rect 6223 27382 6235 27434
rect 6235 27382 6265 27434
rect 6289 27382 6299 27434
rect 6299 27382 6345 27434
rect 6049 27380 6105 27382
rect 6129 27380 6185 27382
rect 6209 27380 6265 27382
rect 6289 27380 6345 27382
rect 9867 27434 9923 27436
rect 9947 27434 10003 27436
rect 10027 27434 10083 27436
rect 10107 27434 10163 27436
rect 9867 27382 9913 27434
rect 9913 27382 9923 27434
rect 9947 27382 9977 27434
rect 9977 27382 9989 27434
rect 9989 27382 10003 27434
rect 10027 27382 10041 27434
rect 10041 27382 10053 27434
rect 10053 27382 10083 27434
rect 10107 27382 10117 27434
rect 10117 27382 10163 27434
rect 9867 27380 9923 27382
rect 9947 27380 10003 27382
rect 10027 27380 10083 27382
rect 10107 27380 10163 27382
rect 13685 27434 13741 27436
rect 13765 27434 13821 27436
rect 13845 27434 13901 27436
rect 13925 27434 13981 27436
rect 13685 27382 13731 27434
rect 13731 27382 13741 27434
rect 13765 27382 13795 27434
rect 13795 27382 13807 27434
rect 13807 27382 13821 27434
rect 13845 27382 13859 27434
rect 13859 27382 13871 27434
rect 13871 27382 13901 27434
rect 13925 27382 13935 27434
rect 13935 27382 13981 27434
rect 13685 27380 13741 27382
rect 13765 27380 13821 27382
rect 13845 27380 13901 27382
rect 13925 27380 13981 27382
rect 6709 26890 6765 26892
rect 6789 26890 6845 26892
rect 6869 26890 6925 26892
rect 6949 26890 7005 26892
rect 6709 26838 6755 26890
rect 6755 26838 6765 26890
rect 6789 26838 6819 26890
rect 6819 26838 6831 26890
rect 6831 26838 6845 26890
rect 6869 26838 6883 26890
rect 6883 26838 6895 26890
rect 6895 26838 6925 26890
rect 6949 26838 6959 26890
rect 6959 26838 7005 26890
rect 6709 26836 6765 26838
rect 6789 26836 6845 26838
rect 6869 26836 6925 26838
rect 6949 26836 7005 26838
rect 10527 26890 10583 26892
rect 10607 26890 10663 26892
rect 10687 26890 10743 26892
rect 10767 26890 10823 26892
rect 10527 26838 10573 26890
rect 10573 26838 10583 26890
rect 10607 26838 10637 26890
rect 10637 26838 10649 26890
rect 10649 26838 10663 26890
rect 10687 26838 10701 26890
rect 10701 26838 10713 26890
rect 10713 26838 10743 26890
rect 10767 26838 10777 26890
rect 10777 26838 10823 26890
rect 10527 26836 10583 26838
rect 10607 26836 10663 26838
rect 10687 26836 10743 26838
rect 10767 26836 10823 26838
rect 6049 26346 6105 26348
rect 6129 26346 6185 26348
rect 6209 26346 6265 26348
rect 6289 26346 6345 26348
rect 6049 26294 6095 26346
rect 6095 26294 6105 26346
rect 6129 26294 6159 26346
rect 6159 26294 6171 26346
rect 6171 26294 6185 26346
rect 6209 26294 6223 26346
rect 6223 26294 6235 26346
rect 6235 26294 6265 26346
rect 6289 26294 6299 26346
rect 6299 26294 6345 26346
rect 6049 26292 6105 26294
rect 6129 26292 6185 26294
rect 6209 26292 6265 26294
rect 6289 26292 6345 26294
rect 9867 26346 9923 26348
rect 9947 26346 10003 26348
rect 10027 26346 10083 26348
rect 10107 26346 10163 26348
rect 9867 26294 9913 26346
rect 9913 26294 9923 26346
rect 9947 26294 9977 26346
rect 9977 26294 9989 26346
rect 9989 26294 10003 26346
rect 10027 26294 10041 26346
rect 10041 26294 10053 26346
rect 10053 26294 10083 26346
rect 10107 26294 10117 26346
rect 10117 26294 10163 26346
rect 9867 26292 9923 26294
rect 9947 26292 10003 26294
rect 10027 26292 10083 26294
rect 10107 26292 10163 26294
rect 6709 25802 6765 25804
rect 6789 25802 6845 25804
rect 6869 25802 6925 25804
rect 6949 25802 7005 25804
rect 6709 25750 6755 25802
rect 6755 25750 6765 25802
rect 6789 25750 6819 25802
rect 6819 25750 6831 25802
rect 6831 25750 6845 25802
rect 6869 25750 6883 25802
rect 6883 25750 6895 25802
rect 6895 25750 6925 25802
rect 6949 25750 6959 25802
rect 6959 25750 7005 25802
rect 6709 25748 6765 25750
rect 6789 25748 6845 25750
rect 6869 25748 6925 25750
rect 6949 25748 7005 25750
rect 10527 25802 10583 25804
rect 10607 25802 10663 25804
rect 10687 25802 10743 25804
rect 10767 25802 10823 25804
rect 10527 25750 10573 25802
rect 10573 25750 10583 25802
rect 10607 25750 10637 25802
rect 10637 25750 10649 25802
rect 10649 25750 10663 25802
rect 10687 25750 10701 25802
rect 10701 25750 10713 25802
rect 10713 25750 10743 25802
rect 10767 25750 10777 25802
rect 10777 25750 10823 25802
rect 10527 25748 10583 25750
rect 10607 25748 10663 25750
rect 10687 25748 10743 25750
rect 10767 25748 10823 25750
rect 6049 25258 6105 25260
rect 6129 25258 6185 25260
rect 6209 25258 6265 25260
rect 6289 25258 6345 25260
rect 6049 25206 6095 25258
rect 6095 25206 6105 25258
rect 6129 25206 6159 25258
rect 6159 25206 6171 25258
rect 6171 25206 6185 25258
rect 6209 25206 6223 25258
rect 6223 25206 6235 25258
rect 6235 25206 6265 25258
rect 6289 25206 6299 25258
rect 6299 25206 6345 25258
rect 6049 25204 6105 25206
rect 6129 25204 6185 25206
rect 6209 25204 6265 25206
rect 6289 25204 6345 25206
rect 9867 25258 9923 25260
rect 9947 25258 10003 25260
rect 10027 25258 10083 25260
rect 10107 25258 10163 25260
rect 9867 25206 9913 25258
rect 9913 25206 9923 25258
rect 9947 25206 9977 25258
rect 9977 25206 9989 25258
rect 9989 25206 10003 25258
rect 10027 25206 10041 25258
rect 10041 25206 10053 25258
rect 10053 25206 10083 25258
rect 10107 25206 10117 25258
rect 10117 25206 10163 25258
rect 9867 25204 9923 25206
rect 9947 25204 10003 25206
rect 10027 25204 10083 25206
rect 10107 25204 10163 25206
rect 6709 24714 6765 24716
rect 6789 24714 6845 24716
rect 6869 24714 6925 24716
rect 6949 24714 7005 24716
rect 6709 24662 6755 24714
rect 6755 24662 6765 24714
rect 6789 24662 6819 24714
rect 6819 24662 6831 24714
rect 6831 24662 6845 24714
rect 6869 24662 6883 24714
rect 6883 24662 6895 24714
rect 6895 24662 6925 24714
rect 6949 24662 6959 24714
rect 6959 24662 7005 24714
rect 6709 24660 6765 24662
rect 6789 24660 6845 24662
rect 6869 24660 6925 24662
rect 6949 24660 7005 24662
rect 10527 24714 10583 24716
rect 10607 24714 10663 24716
rect 10687 24714 10743 24716
rect 10767 24714 10823 24716
rect 10527 24662 10573 24714
rect 10573 24662 10583 24714
rect 10607 24662 10637 24714
rect 10637 24662 10649 24714
rect 10649 24662 10663 24714
rect 10687 24662 10701 24714
rect 10701 24662 10713 24714
rect 10713 24662 10743 24714
rect 10767 24662 10777 24714
rect 10777 24662 10823 24714
rect 10527 24660 10583 24662
rect 10607 24660 10663 24662
rect 10687 24660 10743 24662
rect 10767 24660 10823 24662
rect 6049 24170 6105 24172
rect 6129 24170 6185 24172
rect 6209 24170 6265 24172
rect 6289 24170 6345 24172
rect 6049 24118 6095 24170
rect 6095 24118 6105 24170
rect 6129 24118 6159 24170
rect 6159 24118 6171 24170
rect 6171 24118 6185 24170
rect 6209 24118 6223 24170
rect 6223 24118 6235 24170
rect 6235 24118 6265 24170
rect 6289 24118 6299 24170
rect 6299 24118 6345 24170
rect 6049 24116 6105 24118
rect 6129 24116 6185 24118
rect 6209 24116 6265 24118
rect 6289 24116 6345 24118
rect 9867 24170 9923 24172
rect 9947 24170 10003 24172
rect 10027 24170 10083 24172
rect 10107 24170 10163 24172
rect 9867 24118 9913 24170
rect 9913 24118 9923 24170
rect 9947 24118 9977 24170
rect 9977 24118 9989 24170
rect 9989 24118 10003 24170
rect 10027 24118 10041 24170
rect 10041 24118 10053 24170
rect 10053 24118 10083 24170
rect 10107 24118 10117 24170
rect 10117 24118 10163 24170
rect 9867 24116 9923 24118
rect 9947 24116 10003 24118
rect 10027 24116 10083 24118
rect 10107 24116 10163 24118
rect 6709 23626 6765 23628
rect 6789 23626 6845 23628
rect 6869 23626 6925 23628
rect 6949 23626 7005 23628
rect 6709 23574 6755 23626
rect 6755 23574 6765 23626
rect 6789 23574 6819 23626
rect 6819 23574 6831 23626
rect 6831 23574 6845 23626
rect 6869 23574 6883 23626
rect 6883 23574 6895 23626
rect 6895 23574 6925 23626
rect 6949 23574 6959 23626
rect 6959 23574 7005 23626
rect 6709 23572 6765 23574
rect 6789 23572 6845 23574
rect 6869 23572 6925 23574
rect 6949 23572 7005 23574
rect 10527 23626 10583 23628
rect 10607 23626 10663 23628
rect 10687 23626 10743 23628
rect 10767 23626 10823 23628
rect 10527 23574 10573 23626
rect 10573 23574 10583 23626
rect 10607 23574 10637 23626
rect 10637 23574 10649 23626
rect 10649 23574 10663 23626
rect 10687 23574 10701 23626
rect 10701 23574 10713 23626
rect 10713 23574 10743 23626
rect 10767 23574 10777 23626
rect 10777 23574 10823 23626
rect 10527 23572 10583 23574
rect 10607 23572 10663 23574
rect 10687 23572 10743 23574
rect 10767 23572 10823 23574
rect 6049 23082 6105 23084
rect 6129 23082 6185 23084
rect 6209 23082 6265 23084
rect 6289 23082 6345 23084
rect 6049 23030 6095 23082
rect 6095 23030 6105 23082
rect 6129 23030 6159 23082
rect 6159 23030 6171 23082
rect 6171 23030 6185 23082
rect 6209 23030 6223 23082
rect 6223 23030 6235 23082
rect 6235 23030 6265 23082
rect 6289 23030 6299 23082
rect 6299 23030 6345 23082
rect 6049 23028 6105 23030
rect 6129 23028 6185 23030
rect 6209 23028 6265 23030
rect 6289 23028 6345 23030
rect 9867 23082 9923 23084
rect 9947 23082 10003 23084
rect 10027 23082 10083 23084
rect 10107 23082 10163 23084
rect 9867 23030 9913 23082
rect 9913 23030 9923 23082
rect 9947 23030 9977 23082
rect 9977 23030 9989 23082
rect 9989 23030 10003 23082
rect 10027 23030 10041 23082
rect 10041 23030 10053 23082
rect 10053 23030 10083 23082
rect 10107 23030 10117 23082
rect 10117 23030 10163 23082
rect 9867 23028 9923 23030
rect 9947 23028 10003 23030
rect 10027 23028 10083 23030
rect 10107 23028 10163 23030
rect 6709 22538 6765 22540
rect 6789 22538 6845 22540
rect 6869 22538 6925 22540
rect 6949 22538 7005 22540
rect 6709 22486 6755 22538
rect 6755 22486 6765 22538
rect 6789 22486 6819 22538
rect 6819 22486 6831 22538
rect 6831 22486 6845 22538
rect 6869 22486 6883 22538
rect 6883 22486 6895 22538
rect 6895 22486 6925 22538
rect 6949 22486 6959 22538
rect 6959 22486 7005 22538
rect 6709 22484 6765 22486
rect 6789 22484 6845 22486
rect 6869 22484 6925 22486
rect 6949 22484 7005 22486
rect 10527 22538 10583 22540
rect 10607 22538 10663 22540
rect 10687 22538 10743 22540
rect 10767 22538 10823 22540
rect 10527 22486 10573 22538
rect 10573 22486 10583 22538
rect 10607 22486 10637 22538
rect 10637 22486 10649 22538
rect 10649 22486 10663 22538
rect 10687 22486 10701 22538
rect 10701 22486 10713 22538
rect 10713 22486 10743 22538
rect 10767 22486 10777 22538
rect 10777 22486 10823 22538
rect 10527 22484 10583 22486
rect 10607 22484 10663 22486
rect 10687 22484 10743 22486
rect 10767 22484 10823 22486
rect 6049 21994 6105 21996
rect 6129 21994 6185 21996
rect 6209 21994 6265 21996
rect 6289 21994 6345 21996
rect 6049 21942 6095 21994
rect 6095 21942 6105 21994
rect 6129 21942 6159 21994
rect 6159 21942 6171 21994
rect 6171 21942 6185 21994
rect 6209 21942 6223 21994
rect 6223 21942 6235 21994
rect 6235 21942 6265 21994
rect 6289 21942 6299 21994
rect 6299 21942 6345 21994
rect 6049 21940 6105 21942
rect 6129 21940 6185 21942
rect 6209 21940 6265 21942
rect 6289 21940 6345 21942
rect 9867 21994 9923 21996
rect 9947 21994 10003 21996
rect 10027 21994 10083 21996
rect 10107 21994 10163 21996
rect 9867 21942 9913 21994
rect 9913 21942 9923 21994
rect 9947 21942 9977 21994
rect 9977 21942 9989 21994
rect 9989 21942 10003 21994
rect 10027 21942 10041 21994
rect 10041 21942 10053 21994
rect 10053 21942 10083 21994
rect 10107 21942 10117 21994
rect 10117 21942 10163 21994
rect 9867 21940 9923 21942
rect 9947 21940 10003 21942
rect 10027 21940 10083 21942
rect 10107 21940 10163 21942
rect 6709 21450 6765 21452
rect 6789 21450 6845 21452
rect 6869 21450 6925 21452
rect 6949 21450 7005 21452
rect 6709 21398 6755 21450
rect 6755 21398 6765 21450
rect 6789 21398 6819 21450
rect 6819 21398 6831 21450
rect 6831 21398 6845 21450
rect 6869 21398 6883 21450
rect 6883 21398 6895 21450
rect 6895 21398 6925 21450
rect 6949 21398 6959 21450
rect 6959 21398 7005 21450
rect 6709 21396 6765 21398
rect 6789 21396 6845 21398
rect 6869 21396 6925 21398
rect 6949 21396 7005 21398
rect 10527 21450 10583 21452
rect 10607 21450 10663 21452
rect 10687 21450 10743 21452
rect 10767 21450 10823 21452
rect 10527 21398 10573 21450
rect 10573 21398 10583 21450
rect 10607 21398 10637 21450
rect 10637 21398 10649 21450
rect 10649 21398 10663 21450
rect 10687 21398 10701 21450
rect 10701 21398 10713 21450
rect 10713 21398 10743 21450
rect 10767 21398 10777 21450
rect 10777 21398 10823 21450
rect 10527 21396 10583 21398
rect 10607 21396 10663 21398
rect 10687 21396 10743 21398
rect 10767 21396 10823 21398
rect 6049 20906 6105 20908
rect 6129 20906 6185 20908
rect 6209 20906 6265 20908
rect 6289 20906 6345 20908
rect 6049 20854 6095 20906
rect 6095 20854 6105 20906
rect 6129 20854 6159 20906
rect 6159 20854 6171 20906
rect 6171 20854 6185 20906
rect 6209 20854 6223 20906
rect 6223 20854 6235 20906
rect 6235 20854 6265 20906
rect 6289 20854 6299 20906
rect 6299 20854 6345 20906
rect 6049 20852 6105 20854
rect 6129 20852 6185 20854
rect 6209 20852 6265 20854
rect 6289 20852 6345 20854
rect 9867 20906 9923 20908
rect 9947 20906 10003 20908
rect 10027 20906 10083 20908
rect 10107 20906 10163 20908
rect 9867 20854 9913 20906
rect 9913 20854 9923 20906
rect 9947 20854 9977 20906
rect 9977 20854 9989 20906
rect 9989 20854 10003 20906
rect 10027 20854 10041 20906
rect 10041 20854 10053 20906
rect 10053 20854 10083 20906
rect 10107 20854 10117 20906
rect 10117 20854 10163 20906
rect 9867 20852 9923 20854
rect 9947 20852 10003 20854
rect 10027 20852 10083 20854
rect 10107 20852 10163 20854
rect 6709 20362 6765 20364
rect 6789 20362 6845 20364
rect 6869 20362 6925 20364
rect 6949 20362 7005 20364
rect 6709 20310 6755 20362
rect 6755 20310 6765 20362
rect 6789 20310 6819 20362
rect 6819 20310 6831 20362
rect 6831 20310 6845 20362
rect 6869 20310 6883 20362
rect 6883 20310 6895 20362
rect 6895 20310 6925 20362
rect 6949 20310 6959 20362
rect 6959 20310 7005 20362
rect 6709 20308 6765 20310
rect 6789 20308 6845 20310
rect 6869 20308 6925 20310
rect 6949 20308 7005 20310
rect 10527 20362 10583 20364
rect 10607 20362 10663 20364
rect 10687 20362 10743 20364
rect 10767 20362 10823 20364
rect 10527 20310 10573 20362
rect 10573 20310 10583 20362
rect 10607 20310 10637 20362
rect 10637 20310 10649 20362
rect 10649 20310 10663 20362
rect 10687 20310 10701 20362
rect 10701 20310 10713 20362
rect 10713 20310 10743 20362
rect 10767 20310 10777 20362
rect 10777 20310 10823 20362
rect 10527 20308 10583 20310
rect 10607 20308 10663 20310
rect 10687 20308 10743 20310
rect 10767 20308 10823 20310
rect 6049 19818 6105 19820
rect 6129 19818 6185 19820
rect 6209 19818 6265 19820
rect 6289 19818 6345 19820
rect 6049 19766 6095 19818
rect 6095 19766 6105 19818
rect 6129 19766 6159 19818
rect 6159 19766 6171 19818
rect 6171 19766 6185 19818
rect 6209 19766 6223 19818
rect 6223 19766 6235 19818
rect 6235 19766 6265 19818
rect 6289 19766 6299 19818
rect 6299 19766 6345 19818
rect 6049 19764 6105 19766
rect 6129 19764 6185 19766
rect 6209 19764 6265 19766
rect 6289 19764 6345 19766
rect 9867 19818 9923 19820
rect 9947 19818 10003 19820
rect 10027 19818 10083 19820
rect 10107 19818 10163 19820
rect 9867 19766 9913 19818
rect 9913 19766 9923 19818
rect 9947 19766 9977 19818
rect 9977 19766 9989 19818
rect 9989 19766 10003 19818
rect 10027 19766 10041 19818
rect 10041 19766 10053 19818
rect 10053 19766 10083 19818
rect 10107 19766 10117 19818
rect 10117 19766 10163 19818
rect 9867 19764 9923 19766
rect 9947 19764 10003 19766
rect 10027 19764 10083 19766
rect 10107 19764 10163 19766
rect 6709 19274 6765 19276
rect 6789 19274 6845 19276
rect 6869 19274 6925 19276
rect 6949 19274 7005 19276
rect 6709 19222 6755 19274
rect 6755 19222 6765 19274
rect 6789 19222 6819 19274
rect 6819 19222 6831 19274
rect 6831 19222 6845 19274
rect 6869 19222 6883 19274
rect 6883 19222 6895 19274
rect 6895 19222 6925 19274
rect 6949 19222 6959 19274
rect 6959 19222 7005 19274
rect 6709 19220 6765 19222
rect 6789 19220 6845 19222
rect 6869 19220 6925 19222
rect 6949 19220 7005 19222
rect 10527 19274 10583 19276
rect 10607 19274 10663 19276
rect 10687 19274 10743 19276
rect 10767 19274 10823 19276
rect 10527 19222 10573 19274
rect 10573 19222 10583 19274
rect 10607 19222 10637 19274
rect 10637 19222 10649 19274
rect 10649 19222 10663 19274
rect 10687 19222 10701 19274
rect 10701 19222 10713 19274
rect 10713 19222 10743 19274
rect 10767 19222 10777 19274
rect 10777 19222 10823 19274
rect 10527 19220 10583 19222
rect 10607 19220 10663 19222
rect 10687 19220 10743 19222
rect 10767 19220 10823 19222
rect 6049 18730 6105 18732
rect 6129 18730 6185 18732
rect 6209 18730 6265 18732
rect 6289 18730 6345 18732
rect 6049 18678 6095 18730
rect 6095 18678 6105 18730
rect 6129 18678 6159 18730
rect 6159 18678 6171 18730
rect 6171 18678 6185 18730
rect 6209 18678 6223 18730
rect 6223 18678 6235 18730
rect 6235 18678 6265 18730
rect 6289 18678 6299 18730
rect 6299 18678 6345 18730
rect 6049 18676 6105 18678
rect 6129 18676 6185 18678
rect 6209 18676 6265 18678
rect 6289 18676 6345 18678
rect 9867 18730 9923 18732
rect 9947 18730 10003 18732
rect 10027 18730 10083 18732
rect 10107 18730 10163 18732
rect 9867 18678 9913 18730
rect 9913 18678 9923 18730
rect 9947 18678 9977 18730
rect 9977 18678 9989 18730
rect 9989 18678 10003 18730
rect 10027 18678 10041 18730
rect 10041 18678 10053 18730
rect 10053 18678 10083 18730
rect 10107 18678 10117 18730
rect 10117 18678 10163 18730
rect 9867 18676 9923 18678
rect 9947 18676 10003 18678
rect 10027 18676 10083 18678
rect 10107 18676 10163 18678
rect 6709 18186 6765 18188
rect 6789 18186 6845 18188
rect 6869 18186 6925 18188
rect 6949 18186 7005 18188
rect 6709 18134 6755 18186
rect 6755 18134 6765 18186
rect 6789 18134 6819 18186
rect 6819 18134 6831 18186
rect 6831 18134 6845 18186
rect 6869 18134 6883 18186
rect 6883 18134 6895 18186
rect 6895 18134 6925 18186
rect 6949 18134 6959 18186
rect 6959 18134 7005 18186
rect 6709 18132 6765 18134
rect 6789 18132 6845 18134
rect 6869 18132 6925 18134
rect 6949 18132 7005 18134
rect 10527 18186 10583 18188
rect 10607 18186 10663 18188
rect 10687 18186 10743 18188
rect 10767 18186 10823 18188
rect 10527 18134 10573 18186
rect 10573 18134 10583 18186
rect 10607 18134 10637 18186
rect 10637 18134 10649 18186
rect 10649 18134 10663 18186
rect 10687 18134 10701 18186
rect 10701 18134 10713 18186
rect 10713 18134 10743 18186
rect 10767 18134 10777 18186
rect 10777 18134 10823 18186
rect 10527 18132 10583 18134
rect 10607 18132 10663 18134
rect 10687 18132 10743 18134
rect 10767 18132 10823 18134
rect 6049 17642 6105 17644
rect 6129 17642 6185 17644
rect 6209 17642 6265 17644
rect 6289 17642 6345 17644
rect 6049 17590 6095 17642
rect 6095 17590 6105 17642
rect 6129 17590 6159 17642
rect 6159 17590 6171 17642
rect 6171 17590 6185 17642
rect 6209 17590 6223 17642
rect 6223 17590 6235 17642
rect 6235 17590 6265 17642
rect 6289 17590 6299 17642
rect 6299 17590 6345 17642
rect 6049 17588 6105 17590
rect 6129 17588 6185 17590
rect 6209 17588 6265 17590
rect 6289 17588 6345 17590
rect 9867 17642 9923 17644
rect 9947 17642 10003 17644
rect 10027 17642 10083 17644
rect 10107 17642 10163 17644
rect 9867 17590 9913 17642
rect 9913 17590 9923 17642
rect 9947 17590 9977 17642
rect 9977 17590 9989 17642
rect 9989 17590 10003 17642
rect 10027 17590 10041 17642
rect 10041 17590 10053 17642
rect 10053 17590 10083 17642
rect 10107 17590 10117 17642
rect 10117 17590 10163 17642
rect 9867 17588 9923 17590
rect 9947 17588 10003 17590
rect 10027 17588 10083 17590
rect 10107 17588 10163 17590
rect 6709 17098 6765 17100
rect 6789 17098 6845 17100
rect 6869 17098 6925 17100
rect 6949 17098 7005 17100
rect 6709 17046 6755 17098
rect 6755 17046 6765 17098
rect 6789 17046 6819 17098
rect 6819 17046 6831 17098
rect 6831 17046 6845 17098
rect 6869 17046 6883 17098
rect 6883 17046 6895 17098
rect 6895 17046 6925 17098
rect 6949 17046 6959 17098
rect 6959 17046 7005 17098
rect 6709 17044 6765 17046
rect 6789 17044 6845 17046
rect 6869 17044 6925 17046
rect 6949 17044 7005 17046
rect 10527 17098 10583 17100
rect 10607 17098 10663 17100
rect 10687 17098 10743 17100
rect 10767 17098 10823 17100
rect 10527 17046 10573 17098
rect 10573 17046 10583 17098
rect 10607 17046 10637 17098
rect 10637 17046 10649 17098
rect 10649 17046 10663 17098
rect 10687 17046 10701 17098
rect 10701 17046 10713 17098
rect 10713 17046 10743 17098
rect 10767 17046 10777 17098
rect 10777 17046 10823 17098
rect 10527 17044 10583 17046
rect 10607 17044 10663 17046
rect 10687 17044 10743 17046
rect 10767 17044 10823 17046
rect 6049 16554 6105 16556
rect 6129 16554 6185 16556
rect 6209 16554 6265 16556
rect 6289 16554 6345 16556
rect 6049 16502 6095 16554
rect 6095 16502 6105 16554
rect 6129 16502 6159 16554
rect 6159 16502 6171 16554
rect 6171 16502 6185 16554
rect 6209 16502 6223 16554
rect 6223 16502 6235 16554
rect 6235 16502 6265 16554
rect 6289 16502 6299 16554
rect 6299 16502 6345 16554
rect 6049 16500 6105 16502
rect 6129 16500 6185 16502
rect 6209 16500 6265 16502
rect 6289 16500 6345 16502
rect 9867 16554 9923 16556
rect 9947 16554 10003 16556
rect 10027 16554 10083 16556
rect 10107 16554 10163 16556
rect 9867 16502 9913 16554
rect 9913 16502 9923 16554
rect 9947 16502 9977 16554
rect 9977 16502 9989 16554
rect 9989 16502 10003 16554
rect 10027 16502 10041 16554
rect 10041 16502 10053 16554
rect 10053 16502 10083 16554
rect 10107 16502 10117 16554
rect 10117 16502 10163 16554
rect 9867 16500 9923 16502
rect 9947 16500 10003 16502
rect 10027 16500 10083 16502
rect 10107 16500 10163 16502
rect 6709 16010 6765 16012
rect 6789 16010 6845 16012
rect 6869 16010 6925 16012
rect 6949 16010 7005 16012
rect 6709 15958 6755 16010
rect 6755 15958 6765 16010
rect 6789 15958 6819 16010
rect 6819 15958 6831 16010
rect 6831 15958 6845 16010
rect 6869 15958 6883 16010
rect 6883 15958 6895 16010
rect 6895 15958 6925 16010
rect 6949 15958 6959 16010
rect 6959 15958 7005 16010
rect 6709 15956 6765 15958
rect 6789 15956 6845 15958
rect 6869 15956 6925 15958
rect 6949 15956 7005 15958
rect 10527 16010 10583 16012
rect 10607 16010 10663 16012
rect 10687 16010 10743 16012
rect 10767 16010 10823 16012
rect 10527 15958 10573 16010
rect 10573 15958 10583 16010
rect 10607 15958 10637 16010
rect 10637 15958 10649 16010
rect 10649 15958 10663 16010
rect 10687 15958 10701 16010
rect 10701 15958 10713 16010
rect 10713 15958 10743 16010
rect 10767 15958 10777 16010
rect 10777 15958 10823 16010
rect 10527 15956 10583 15958
rect 10607 15956 10663 15958
rect 10687 15956 10743 15958
rect 10767 15956 10823 15958
rect 6049 15466 6105 15468
rect 6129 15466 6185 15468
rect 6209 15466 6265 15468
rect 6289 15466 6345 15468
rect 6049 15414 6095 15466
rect 6095 15414 6105 15466
rect 6129 15414 6159 15466
rect 6159 15414 6171 15466
rect 6171 15414 6185 15466
rect 6209 15414 6223 15466
rect 6223 15414 6235 15466
rect 6235 15414 6265 15466
rect 6289 15414 6299 15466
rect 6299 15414 6345 15466
rect 6049 15412 6105 15414
rect 6129 15412 6185 15414
rect 6209 15412 6265 15414
rect 6289 15412 6345 15414
rect 9867 15466 9923 15468
rect 9947 15466 10003 15468
rect 10027 15466 10083 15468
rect 10107 15466 10163 15468
rect 9867 15414 9913 15466
rect 9913 15414 9923 15466
rect 9947 15414 9977 15466
rect 9977 15414 9989 15466
rect 9989 15414 10003 15466
rect 10027 15414 10041 15466
rect 10041 15414 10053 15466
rect 10053 15414 10083 15466
rect 10107 15414 10117 15466
rect 10117 15414 10163 15466
rect 9867 15412 9923 15414
rect 9947 15412 10003 15414
rect 10027 15412 10083 15414
rect 10107 15412 10163 15414
rect 6709 14922 6765 14924
rect 6789 14922 6845 14924
rect 6869 14922 6925 14924
rect 6949 14922 7005 14924
rect 6709 14870 6755 14922
rect 6755 14870 6765 14922
rect 6789 14870 6819 14922
rect 6819 14870 6831 14922
rect 6831 14870 6845 14922
rect 6869 14870 6883 14922
rect 6883 14870 6895 14922
rect 6895 14870 6925 14922
rect 6949 14870 6959 14922
rect 6959 14870 7005 14922
rect 6709 14868 6765 14870
rect 6789 14868 6845 14870
rect 6869 14868 6925 14870
rect 6949 14868 7005 14870
rect 10527 14922 10583 14924
rect 10607 14922 10663 14924
rect 10687 14922 10743 14924
rect 10767 14922 10823 14924
rect 10527 14870 10573 14922
rect 10573 14870 10583 14922
rect 10607 14870 10637 14922
rect 10637 14870 10649 14922
rect 10649 14870 10663 14922
rect 10687 14870 10701 14922
rect 10701 14870 10713 14922
rect 10713 14870 10743 14922
rect 10767 14870 10777 14922
rect 10777 14870 10823 14922
rect 10527 14868 10583 14870
rect 10607 14868 10663 14870
rect 10687 14868 10743 14870
rect 10767 14868 10823 14870
rect 14345 26890 14401 26892
rect 14425 26890 14481 26892
rect 14505 26890 14561 26892
rect 14585 26890 14641 26892
rect 14345 26838 14391 26890
rect 14391 26838 14401 26890
rect 14425 26838 14455 26890
rect 14455 26838 14467 26890
rect 14467 26838 14481 26890
rect 14505 26838 14519 26890
rect 14519 26838 14531 26890
rect 14531 26838 14561 26890
rect 14585 26838 14595 26890
rect 14595 26838 14641 26890
rect 14345 26836 14401 26838
rect 14425 26836 14481 26838
rect 14505 26836 14561 26838
rect 14585 26836 14641 26838
rect 13685 26346 13741 26348
rect 13765 26346 13821 26348
rect 13845 26346 13901 26348
rect 13925 26346 13981 26348
rect 13685 26294 13731 26346
rect 13731 26294 13741 26346
rect 13765 26294 13795 26346
rect 13795 26294 13807 26346
rect 13807 26294 13821 26346
rect 13845 26294 13859 26346
rect 13859 26294 13871 26346
rect 13871 26294 13901 26346
rect 13925 26294 13935 26346
rect 13935 26294 13981 26346
rect 13685 26292 13741 26294
rect 13765 26292 13821 26294
rect 13845 26292 13901 26294
rect 13925 26292 13981 26294
rect 14345 25802 14401 25804
rect 14425 25802 14481 25804
rect 14505 25802 14561 25804
rect 14585 25802 14641 25804
rect 14345 25750 14391 25802
rect 14391 25750 14401 25802
rect 14425 25750 14455 25802
rect 14455 25750 14467 25802
rect 14467 25750 14481 25802
rect 14505 25750 14519 25802
rect 14519 25750 14531 25802
rect 14531 25750 14561 25802
rect 14585 25750 14595 25802
rect 14595 25750 14641 25802
rect 14345 25748 14401 25750
rect 14425 25748 14481 25750
rect 14505 25748 14561 25750
rect 14585 25748 14641 25750
rect 17503 27434 17559 27436
rect 17583 27434 17639 27436
rect 17663 27434 17719 27436
rect 17743 27434 17799 27436
rect 17503 27382 17549 27434
rect 17549 27382 17559 27434
rect 17583 27382 17613 27434
rect 17613 27382 17625 27434
rect 17625 27382 17639 27434
rect 17663 27382 17677 27434
rect 17677 27382 17689 27434
rect 17689 27382 17719 27434
rect 17743 27382 17753 27434
rect 17753 27382 17799 27434
rect 17503 27380 17559 27382
rect 17583 27380 17639 27382
rect 17663 27380 17719 27382
rect 17743 27380 17799 27382
rect 18163 26890 18219 26892
rect 18243 26890 18299 26892
rect 18323 26890 18379 26892
rect 18403 26890 18459 26892
rect 18163 26838 18209 26890
rect 18209 26838 18219 26890
rect 18243 26838 18273 26890
rect 18273 26838 18285 26890
rect 18285 26838 18299 26890
rect 18323 26838 18337 26890
rect 18337 26838 18349 26890
rect 18349 26838 18379 26890
rect 18403 26838 18413 26890
rect 18413 26838 18459 26890
rect 18163 26836 18219 26838
rect 18243 26836 18299 26838
rect 18323 26836 18379 26838
rect 18403 26836 18459 26838
rect 17503 26346 17559 26348
rect 17583 26346 17639 26348
rect 17663 26346 17719 26348
rect 17743 26346 17799 26348
rect 17503 26294 17549 26346
rect 17549 26294 17559 26346
rect 17583 26294 17613 26346
rect 17613 26294 17625 26346
rect 17625 26294 17639 26346
rect 17663 26294 17677 26346
rect 17677 26294 17689 26346
rect 17689 26294 17719 26346
rect 17743 26294 17753 26346
rect 17753 26294 17799 26346
rect 17503 26292 17559 26294
rect 17583 26292 17639 26294
rect 17663 26292 17719 26294
rect 17743 26292 17799 26294
rect 18163 25802 18219 25804
rect 18243 25802 18299 25804
rect 18323 25802 18379 25804
rect 18403 25802 18459 25804
rect 18163 25750 18209 25802
rect 18209 25750 18219 25802
rect 18243 25750 18273 25802
rect 18273 25750 18285 25802
rect 18285 25750 18299 25802
rect 18323 25750 18337 25802
rect 18337 25750 18349 25802
rect 18349 25750 18379 25802
rect 18403 25750 18413 25802
rect 18413 25750 18459 25802
rect 18163 25748 18219 25750
rect 18243 25748 18299 25750
rect 18323 25748 18379 25750
rect 18403 25748 18459 25750
rect 13685 25258 13741 25260
rect 13765 25258 13821 25260
rect 13845 25258 13901 25260
rect 13925 25258 13981 25260
rect 13685 25206 13731 25258
rect 13731 25206 13741 25258
rect 13765 25206 13795 25258
rect 13795 25206 13807 25258
rect 13807 25206 13821 25258
rect 13845 25206 13859 25258
rect 13859 25206 13871 25258
rect 13871 25206 13901 25258
rect 13925 25206 13935 25258
rect 13935 25206 13981 25258
rect 13685 25204 13741 25206
rect 13765 25204 13821 25206
rect 13845 25204 13901 25206
rect 13925 25204 13981 25206
rect 13685 24170 13741 24172
rect 13765 24170 13821 24172
rect 13845 24170 13901 24172
rect 13925 24170 13981 24172
rect 13685 24118 13731 24170
rect 13731 24118 13741 24170
rect 13765 24118 13795 24170
rect 13795 24118 13807 24170
rect 13807 24118 13821 24170
rect 13845 24118 13859 24170
rect 13859 24118 13871 24170
rect 13871 24118 13901 24170
rect 13925 24118 13935 24170
rect 13935 24118 13981 24170
rect 13685 24116 13741 24118
rect 13765 24116 13821 24118
rect 13845 24116 13901 24118
rect 13925 24116 13981 24118
rect 13685 23082 13741 23084
rect 13765 23082 13821 23084
rect 13845 23082 13901 23084
rect 13925 23082 13981 23084
rect 13685 23030 13731 23082
rect 13731 23030 13741 23082
rect 13765 23030 13795 23082
rect 13795 23030 13807 23082
rect 13807 23030 13821 23082
rect 13845 23030 13859 23082
rect 13859 23030 13871 23082
rect 13871 23030 13901 23082
rect 13925 23030 13935 23082
rect 13935 23030 13981 23082
rect 13685 23028 13741 23030
rect 13765 23028 13821 23030
rect 13845 23028 13901 23030
rect 13925 23028 13981 23030
rect 13685 21994 13741 21996
rect 13765 21994 13821 21996
rect 13845 21994 13901 21996
rect 13925 21994 13981 21996
rect 13685 21942 13731 21994
rect 13731 21942 13741 21994
rect 13765 21942 13795 21994
rect 13795 21942 13807 21994
rect 13807 21942 13821 21994
rect 13845 21942 13859 21994
rect 13859 21942 13871 21994
rect 13871 21942 13901 21994
rect 13925 21942 13935 21994
rect 13935 21942 13981 21994
rect 13685 21940 13741 21942
rect 13765 21940 13821 21942
rect 13845 21940 13901 21942
rect 13925 21940 13981 21942
rect 13685 20906 13741 20908
rect 13765 20906 13821 20908
rect 13845 20906 13901 20908
rect 13925 20906 13981 20908
rect 13685 20854 13731 20906
rect 13731 20854 13741 20906
rect 13765 20854 13795 20906
rect 13795 20854 13807 20906
rect 13807 20854 13821 20906
rect 13845 20854 13859 20906
rect 13859 20854 13871 20906
rect 13871 20854 13901 20906
rect 13925 20854 13935 20906
rect 13935 20854 13981 20906
rect 13685 20852 13741 20854
rect 13765 20852 13821 20854
rect 13845 20852 13901 20854
rect 13925 20852 13981 20854
rect 13685 19818 13741 19820
rect 13765 19818 13821 19820
rect 13845 19818 13901 19820
rect 13925 19818 13981 19820
rect 13685 19766 13731 19818
rect 13731 19766 13741 19818
rect 13765 19766 13795 19818
rect 13795 19766 13807 19818
rect 13807 19766 13821 19818
rect 13845 19766 13859 19818
rect 13859 19766 13871 19818
rect 13871 19766 13901 19818
rect 13925 19766 13935 19818
rect 13935 19766 13981 19818
rect 13685 19764 13741 19766
rect 13765 19764 13821 19766
rect 13845 19764 13901 19766
rect 13925 19764 13981 19766
rect 13685 18730 13741 18732
rect 13765 18730 13821 18732
rect 13845 18730 13901 18732
rect 13925 18730 13981 18732
rect 13685 18678 13731 18730
rect 13731 18678 13741 18730
rect 13765 18678 13795 18730
rect 13795 18678 13807 18730
rect 13807 18678 13821 18730
rect 13845 18678 13859 18730
rect 13859 18678 13871 18730
rect 13871 18678 13901 18730
rect 13925 18678 13935 18730
rect 13935 18678 13981 18730
rect 13685 18676 13741 18678
rect 13765 18676 13821 18678
rect 13845 18676 13901 18678
rect 13925 18676 13981 18678
rect 13685 17642 13741 17644
rect 13765 17642 13821 17644
rect 13845 17642 13901 17644
rect 13925 17642 13981 17644
rect 13685 17590 13731 17642
rect 13731 17590 13741 17642
rect 13765 17590 13795 17642
rect 13795 17590 13807 17642
rect 13807 17590 13821 17642
rect 13845 17590 13859 17642
rect 13859 17590 13871 17642
rect 13871 17590 13901 17642
rect 13925 17590 13935 17642
rect 13935 17590 13981 17642
rect 13685 17588 13741 17590
rect 13765 17588 13821 17590
rect 13845 17588 13901 17590
rect 13925 17588 13981 17590
rect 13685 16554 13741 16556
rect 13765 16554 13821 16556
rect 13845 16554 13901 16556
rect 13925 16554 13981 16556
rect 13685 16502 13731 16554
rect 13731 16502 13741 16554
rect 13765 16502 13795 16554
rect 13795 16502 13807 16554
rect 13807 16502 13821 16554
rect 13845 16502 13859 16554
rect 13859 16502 13871 16554
rect 13871 16502 13901 16554
rect 13925 16502 13935 16554
rect 13935 16502 13981 16554
rect 13685 16500 13741 16502
rect 13765 16500 13821 16502
rect 13845 16500 13901 16502
rect 13925 16500 13981 16502
rect 13685 15466 13741 15468
rect 13765 15466 13821 15468
rect 13845 15466 13901 15468
rect 13925 15466 13981 15468
rect 13685 15414 13731 15466
rect 13731 15414 13741 15466
rect 13765 15414 13795 15466
rect 13795 15414 13807 15466
rect 13807 15414 13821 15466
rect 13845 15414 13859 15466
rect 13859 15414 13871 15466
rect 13871 15414 13901 15466
rect 13925 15414 13935 15466
rect 13935 15414 13981 15466
rect 13685 15412 13741 15414
rect 13765 15412 13821 15414
rect 13845 15412 13901 15414
rect 13925 15412 13981 15414
rect 6049 14378 6105 14380
rect 6129 14378 6185 14380
rect 6209 14378 6265 14380
rect 6289 14378 6345 14380
rect 6049 14326 6095 14378
rect 6095 14326 6105 14378
rect 6129 14326 6159 14378
rect 6159 14326 6171 14378
rect 6171 14326 6185 14378
rect 6209 14326 6223 14378
rect 6223 14326 6235 14378
rect 6235 14326 6265 14378
rect 6289 14326 6299 14378
rect 6299 14326 6345 14378
rect 6049 14324 6105 14326
rect 6129 14324 6185 14326
rect 6209 14324 6265 14326
rect 6289 14324 6345 14326
rect 9867 14378 9923 14380
rect 9947 14378 10003 14380
rect 10027 14378 10083 14380
rect 10107 14378 10163 14380
rect 9867 14326 9913 14378
rect 9913 14326 9923 14378
rect 9947 14326 9977 14378
rect 9977 14326 9989 14378
rect 9989 14326 10003 14378
rect 10027 14326 10041 14378
rect 10041 14326 10053 14378
rect 10053 14326 10083 14378
rect 10107 14326 10117 14378
rect 10117 14326 10163 14378
rect 9867 14324 9923 14326
rect 9947 14324 10003 14326
rect 10027 14324 10083 14326
rect 10107 14324 10163 14326
rect 6709 13834 6765 13836
rect 6789 13834 6845 13836
rect 6869 13834 6925 13836
rect 6949 13834 7005 13836
rect 6709 13782 6755 13834
rect 6755 13782 6765 13834
rect 6789 13782 6819 13834
rect 6819 13782 6831 13834
rect 6831 13782 6845 13834
rect 6869 13782 6883 13834
rect 6883 13782 6895 13834
rect 6895 13782 6925 13834
rect 6949 13782 6959 13834
rect 6959 13782 7005 13834
rect 6709 13780 6765 13782
rect 6789 13780 6845 13782
rect 6869 13780 6925 13782
rect 6949 13780 7005 13782
rect 6049 13290 6105 13292
rect 6129 13290 6185 13292
rect 6209 13290 6265 13292
rect 6289 13290 6345 13292
rect 6049 13238 6095 13290
rect 6095 13238 6105 13290
rect 6129 13238 6159 13290
rect 6159 13238 6171 13290
rect 6171 13238 6185 13290
rect 6209 13238 6223 13290
rect 6223 13238 6235 13290
rect 6235 13238 6265 13290
rect 6289 13238 6299 13290
rect 6299 13238 6345 13290
rect 6049 13236 6105 13238
rect 6129 13236 6185 13238
rect 6209 13236 6265 13238
rect 6289 13236 6345 13238
rect 6709 12746 6765 12748
rect 6789 12746 6845 12748
rect 6869 12746 6925 12748
rect 6949 12746 7005 12748
rect 6709 12694 6755 12746
rect 6755 12694 6765 12746
rect 6789 12694 6819 12746
rect 6819 12694 6831 12746
rect 6831 12694 6845 12746
rect 6869 12694 6883 12746
rect 6883 12694 6895 12746
rect 6895 12694 6925 12746
rect 6949 12694 6959 12746
rect 6959 12694 7005 12746
rect 6709 12692 6765 12694
rect 6789 12692 6845 12694
rect 6869 12692 6925 12694
rect 6949 12692 7005 12694
rect 9867 13290 9923 13292
rect 9947 13290 10003 13292
rect 10027 13290 10083 13292
rect 10107 13290 10163 13292
rect 9867 13238 9913 13290
rect 9913 13238 9923 13290
rect 9947 13238 9977 13290
rect 9977 13238 9989 13290
rect 9989 13238 10003 13290
rect 10027 13238 10041 13290
rect 10041 13238 10053 13290
rect 10053 13238 10083 13290
rect 10107 13238 10117 13290
rect 10117 13238 10163 13290
rect 9867 13236 9923 13238
rect 9947 13236 10003 13238
rect 10027 13236 10083 13238
rect 10107 13236 10163 13238
rect 10527 13834 10583 13836
rect 10607 13834 10663 13836
rect 10687 13834 10743 13836
rect 10767 13834 10823 13836
rect 10527 13782 10573 13834
rect 10573 13782 10583 13834
rect 10607 13782 10637 13834
rect 10637 13782 10649 13834
rect 10649 13782 10663 13834
rect 10687 13782 10701 13834
rect 10701 13782 10713 13834
rect 10713 13782 10743 13834
rect 10767 13782 10777 13834
rect 10777 13782 10823 13834
rect 10527 13780 10583 13782
rect 10607 13780 10663 13782
rect 10687 13780 10743 13782
rect 10767 13780 10823 13782
rect 10527 12746 10583 12748
rect 10607 12746 10663 12748
rect 10687 12746 10743 12748
rect 10767 12746 10823 12748
rect 10527 12694 10573 12746
rect 10573 12694 10583 12746
rect 10607 12694 10637 12746
rect 10637 12694 10649 12746
rect 10649 12694 10663 12746
rect 10687 12694 10701 12746
rect 10701 12694 10713 12746
rect 10713 12694 10743 12746
rect 10767 12694 10777 12746
rect 10777 12694 10823 12746
rect 10527 12692 10583 12694
rect 10607 12692 10663 12694
rect 10687 12692 10743 12694
rect 10767 12692 10823 12694
rect 6049 12202 6105 12204
rect 6129 12202 6185 12204
rect 6209 12202 6265 12204
rect 6289 12202 6345 12204
rect 6049 12150 6095 12202
rect 6095 12150 6105 12202
rect 6129 12150 6159 12202
rect 6159 12150 6171 12202
rect 6171 12150 6185 12202
rect 6209 12150 6223 12202
rect 6223 12150 6235 12202
rect 6235 12150 6265 12202
rect 6289 12150 6299 12202
rect 6299 12150 6345 12202
rect 6049 12148 6105 12150
rect 6129 12148 6185 12150
rect 6209 12148 6265 12150
rect 6289 12148 6345 12150
rect 9867 12202 9923 12204
rect 9947 12202 10003 12204
rect 10027 12202 10083 12204
rect 10107 12202 10163 12204
rect 9867 12150 9913 12202
rect 9913 12150 9923 12202
rect 9947 12150 9977 12202
rect 9977 12150 9989 12202
rect 9989 12150 10003 12202
rect 10027 12150 10041 12202
rect 10041 12150 10053 12202
rect 10053 12150 10083 12202
rect 10107 12150 10117 12202
rect 10117 12150 10163 12202
rect 9867 12148 9923 12150
rect 9947 12148 10003 12150
rect 10027 12148 10083 12150
rect 10107 12148 10163 12150
rect 13685 14378 13741 14380
rect 13765 14378 13821 14380
rect 13845 14378 13901 14380
rect 13925 14378 13981 14380
rect 13685 14326 13731 14378
rect 13731 14326 13741 14378
rect 13765 14326 13795 14378
rect 13795 14326 13807 14378
rect 13807 14326 13821 14378
rect 13845 14326 13859 14378
rect 13859 14326 13871 14378
rect 13871 14326 13901 14378
rect 13925 14326 13935 14378
rect 13935 14326 13981 14378
rect 13685 14324 13741 14326
rect 13765 14324 13821 14326
rect 13845 14324 13901 14326
rect 13925 14324 13981 14326
rect 17503 25258 17559 25260
rect 17583 25258 17639 25260
rect 17663 25258 17719 25260
rect 17743 25258 17799 25260
rect 17503 25206 17549 25258
rect 17549 25206 17559 25258
rect 17583 25206 17613 25258
rect 17613 25206 17625 25258
rect 17625 25206 17639 25258
rect 17663 25206 17677 25258
rect 17677 25206 17689 25258
rect 17689 25206 17719 25258
rect 17743 25206 17753 25258
rect 17753 25206 17799 25258
rect 17503 25204 17559 25206
rect 17583 25204 17639 25206
rect 17663 25204 17719 25206
rect 17743 25204 17799 25206
rect 14345 24714 14401 24716
rect 14425 24714 14481 24716
rect 14505 24714 14561 24716
rect 14585 24714 14641 24716
rect 14345 24662 14391 24714
rect 14391 24662 14401 24714
rect 14425 24662 14455 24714
rect 14455 24662 14467 24714
rect 14467 24662 14481 24714
rect 14505 24662 14519 24714
rect 14519 24662 14531 24714
rect 14531 24662 14561 24714
rect 14585 24662 14595 24714
rect 14595 24662 14641 24714
rect 14345 24660 14401 24662
rect 14425 24660 14481 24662
rect 14505 24660 14561 24662
rect 14585 24660 14641 24662
rect 18163 24714 18219 24716
rect 18243 24714 18299 24716
rect 18323 24714 18379 24716
rect 18403 24714 18459 24716
rect 18163 24662 18209 24714
rect 18209 24662 18219 24714
rect 18243 24662 18273 24714
rect 18273 24662 18285 24714
rect 18285 24662 18299 24714
rect 18323 24662 18337 24714
rect 18337 24662 18349 24714
rect 18349 24662 18379 24714
rect 18403 24662 18413 24714
rect 18413 24662 18459 24714
rect 18163 24660 18219 24662
rect 18243 24660 18299 24662
rect 18323 24660 18379 24662
rect 18403 24660 18459 24662
rect 17503 24170 17559 24172
rect 17583 24170 17639 24172
rect 17663 24170 17719 24172
rect 17743 24170 17799 24172
rect 17503 24118 17549 24170
rect 17549 24118 17559 24170
rect 17583 24118 17613 24170
rect 17613 24118 17625 24170
rect 17625 24118 17639 24170
rect 17663 24118 17677 24170
rect 17677 24118 17689 24170
rect 17689 24118 17719 24170
rect 17743 24118 17753 24170
rect 17753 24118 17799 24170
rect 17503 24116 17559 24118
rect 17583 24116 17639 24118
rect 17663 24116 17719 24118
rect 17743 24116 17799 24118
rect 14345 23626 14401 23628
rect 14425 23626 14481 23628
rect 14505 23626 14561 23628
rect 14585 23626 14641 23628
rect 14345 23574 14391 23626
rect 14391 23574 14401 23626
rect 14425 23574 14455 23626
rect 14455 23574 14467 23626
rect 14467 23574 14481 23626
rect 14505 23574 14519 23626
rect 14519 23574 14531 23626
rect 14531 23574 14561 23626
rect 14585 23574 14595 23626
rect 14595 23574 14641 23626
rect 14345 23572 14401 23574
rect 14425 23572 14481 23574
rect 14505 23572 14561 23574
rect 14585 23572 14641 23574
rect 18163 23626 18219 23628
rect 18243 23626 18299 23628
rect 18323 23626 18379 23628
rect 18403 23626 18459 23628
rect 18163 23574 18209 23626
rect 18209 23574 18219 23626
rect 18243 23574 18273 23626
rect 18273 23574 18285 23626
rect 18285 23574 18299 23626
rect 18323 23574 18337 23626
rect 18337 23574 18349 23626
rect 18349 23574 18379 23626
rect 18403 23574 18413 23626
rect 18413 23574 18459 23626
rect 18163 23572 18219 23574
rect 18243 23572 18299 23574
rect 18323 23572 18379 23574
rect 18403 23572 18459 23574
rect 17503 23082 17559 23084
rect 17583 23082 17639 23084
rect 17663 23082 17719 23084
rect 17743 23082 17799 23084
rect 17503 23030 17549 23082
rect 17549 23030 17559 23082
rect 17583 23030 17613 23082
rect 17613 23030 17625 23082
rect 17625 23030 17639 23082
rect 17663 23030 17677 23082
rect 17677 23030 17689 23082
rect 17689 23030 17719 23082
rect 17743 23030 17753 23082
rect 17753 23030 17799 23082
rect 17503 23028 17559 23030
rect 17583 23028 17639 23030
rect 17663 23028 17719 23030
rect 17743 23028 17799 23030
rect 14345 22538 14401 22540
rect 14425 22538 14481 22540
rect 14505 22538 14561 22540
rect 14585 22538 14641 22540
rect 14345 22486 14391 22538
rect 14391 22486 14401 22538
rect 14425 22486 14455 22538
rect 14455 22486 14467 22538
rect 14467 22486 14481 22538
rect 14505 22486 14519 22538
rect 14519 22486 14531 22538
rect 14531 22486 14561 22538
rect 14585 22486 14595 22538
rect 14595 22486 14641 22538
rect 14345 22484 14401 22486
rect 14425 22484 14481 22486
rect 14505 22484 14561 22486
rect 14585 22484 14641 22486
rect 18163 22538 18219 22540
rect 18243 22538 18299 22540
rect 18323 22538 18379 22540
rect 18403 22538 18459 22540
rect 18163 22486 18209 22538
rect 18209 22486 18219 22538
rect 18243 22486 18273 22538
rect 18273 22486 18285 22538
rect 18285 22486 18299 22538
rect 18323 22486 18337 22538
rect 18337 22486 18349 22538
rect 18349 22486 18379 22538
rect 18403 22486 18413 22538
rect 18413 22486 18459 22538
rect 18163 22484 18219 22486
rect 18243 22484 18299 22486
rect 18323 22484 18379 22486
rect 18403 22484 18459 22486
rect 17503 21994 17559 21996
rect 17583 21994 17639 21996
rect 17663 21994 17719 21996
rect 17743 21994 17799 21996
rect 17503 21942 17549 21994
rect 17549 21942 17559 21994
rect 17583 21942 17613 21994
rect 17613 21942 17625 21994
rect 17625 21942 17639 21994
rect 17663 21942 17677 21994
rect 17677 21942 17689 21994
rect 17689 21942 17719 21994
rect 17743 21942 17753 21994
rect 17753 21942 17799 21994
rect 17503 21940 17559 21942
rect 17583 21940 17639 21942
rect 17663 21940 17719 21942
rect 17743 21940 17799 21942
rect 14345 21450 14401 21452
rect 14425 21450 14481 21452
rect 14505 21450 14561 21452
rect 14585 21450 14641 21452
rect 14345 21398 14391 21450
rect 14391 21398 14401 21450
rect 14425 21398 14455 21450
rect 14455 21398 14467 21450
rect 14467 21398 14481 21450
rect 14505 21398 14519 21450
rect 14519 21398 14531 21450
rect 14531 21398 14561 21450
rect 14585 21398 14595 21450
rect 14595 21398 14641 21450
rect 14345 21396 14401 21398
rect 14425 21396 14481 21398
rect 14505 21396 14561 21398
rect 14585 21396 14641 21398
rect 18163 21450 18219 21452
rect 18243 21450 18299 21452
rect 18323 21450 18379 21452
rect 18403 21450 18459 21452
rect 18163 21398 18209 21450
rect 18209 21398 18219 21450
rect 18243 21398 18273 21450
rect 18273 21398 18285 21450
rect 18285 21398 18299 21450
rect 18323 21398 18337 21450
rect 18337 21398 18349 21450
rect 18349 21398 18379 21450
rect 18403 21398 18413 21450
rect 18413 21398 18459 21450
rect 18163 21396 18219 21398
rect 18243 21396 18299 21398
rect 18323 21396 18379 21398
rect 18403 21396 18459 21398
rect 17503 20906 17559 20908
rect 17583 20906 17639 20908
rect 17663 20906 17719 20908
rect 17743 20906 17799 20908
rect 17503 20854 17549 20906
rect 17549 20854 17559 20906
rect 17583 20854 17613 20906
rect 17613 20854 17625 20906
rect 17625 20854 17639 20906
rect 17663 20854 17677 20906
rect 17677 20854 17689 20906
rect 17689 20854 17719 20906
rect 17743 20854 17753 20906
rect 17753 20854 17799 20906
rect 17503 20852 17559 20854
rect 17583 20852 17639 20854
rect 17663 20852 17719 20854
rect 17743 20852 17799 20854
rect 14345 20362 14401 20364
rect 14425 20362 14481 20364
rect 14505 20362 14561 20364
rect 14585 20362 14641 20364
rect 14345 20310 14391 20362
rect 14391 20310 14401 20362
rect 14425 20310 14455 20362
rect 14455 20310 14467 20362
rect 14467 20310 14481 20362
rect 14505 20310 14519 20362
rect 14519 20310 14531 20362
rect 14531 20310 14561 20362
rect 14585 20310 14595 20362
rect 14595 20310 14641 20362
rect 14345 20308 14401 20310
rect 14425 20308 14481 20310
rect 14505 20308 14561 20310
rect 14585 20308 14641 20310
rect 18163 20362 18219 20364
rect 18243 20362 18299 20364
rect 18323 20362 18379 20364
rect 18403 20362 18459 20364
rect 18163 20310 18209 20362
rect 18209 20310 18219 20362
rect 18243 20310 18273 20362
rect 18273 20310 18285 20362
rect 18285 20310 18299 20362
rect 18323 20310 18337 20362
rect 18337 20310 18349 20362
rect 18349 20310 18379 20362
rect 18403 20310 18413 20362
rect 18413 20310 18459 20362
rect 18163 20308 18219 20310
rect 18243 20308 18299 20310
rect 18323 20308 18379 20310
rect 18403 20308 18459 20310
rect 17503 19818 17559 19820
rect 17583 19818 17639 19820
rect 17663 19818 17719 19820
rect 17743 19818 17799 19820
rect 17503 19766 17549 19818
rect 17549 19766 17559 19818
rect 17583 19766 17613 19818
rect 17613 19766 17625 19818
rect 17625 19766 17639 19818
rect 17663 19766 17677 19818
rect 17677 19766 17689 19818
rect 17689 19766 17719 19818
rect 17743 19766 17753 19818
rect 17753 19766 17799 19818
rect 17503 19764 17559 19766
rect 17583 19764 17639 19766
rect 17663 19764 17719 19766
rect 17743 19764 17799 19766
rect 14345 19274 14401 19276
rect 14425 19274 14481 19276
rect 14505 19274 14561 19276
rect 14585 19274 14641 19276
rect 14345 19222 14391 19274
rect 14391 19222 14401 19274
rect 14425 19222 14455 19274
rect 14455 19222 14467 19274
rect 14467 19222 14481 19274
rect 14505 19222 14519 19274
rect 14519 19222 14531 19274
rect 14531 19222 14561 19274
rect 14585 19222 14595 19274
rect 14595 19222 14641 19274
rect 14345 19220 14401 19222
rect 14425 19220 14481 19222
rect 14505 19220 14561 19222
rect 14585 19220 14641 19222
rect 18163 19274 18219 19276
rect 18243 19274 18299 19276
rect 18323 19274 18379 19276
rect 18403 19274 18459 19276
rect 18163 19222 18209 19274
rect 18209 19222 18219 19274
rect 18243 19222 18273 19274
rect 18273 19222 18285 19274
rect 18285 19222 18299 19274
rect 18323 19222 18337 19274
rect 18337 19222 18349 19274
rect 18349 19222 18379 19274
rect 18403 19222 18413 19274
rect 18413 19222 18459 19274
rect 18163 19220 18219 19222
rect 18243 19220 18299 19222
rect 18323 19220 18379 19222
rect 18403 19220 18459 19222
rect 17503 18730 17559 18732
rect 17583 18730 17639 18732
rect 17663 18730 17719 18732
rect 17743 18730 17799 18732
rect 17503 18678 17549 18730
rect 17549 18678 17559 18730
rect 17583 18678 17613 18730
rect 17613 18678 17625 18730
rect 17625 18678 17639 18730
rect 17663 18678 17677 18730
rect 17677 18678 17689 18730
rect 17689 18678 17719 18730
rect 17743 18678 17753 18730
rect 17753 18678 17799 18730
rect 17503 18676 17559 18678
rect 17583 18676 17639 18678
rect 17663 18676 17719 18678
rect 17743 18676 17799 18678
rect 14345 18186 14401 18188
rect 14425 18186 14481 18188
rect 14505 18186 14561 18188
rect 14585 18186 14641 18188
rect 14345 18134 14391 18186
rect 14391 18134 14401 18186
rect 14425 18134 14455 18186
rect 14455 18134 14467 18186
rect 14467 18134 14481 18186
rect 14505 18134 14519 18186
rect 14519 18134 14531 18186
rect 14531 18134 14561 18186
rect 14585 18134 14595 18186
rect 14595 18134 14641 18186
rect 14345 18132 14401 18134
rect 14425 18132 14481 18134
rect 14505 18132 14561 18134
rect 14585 18132 14641 18134
rect 18163 18186 18219 18188
rect 18243 18186 18299 18188
rect 18323 18186 18379 18188
rect 18403 18186 18459 18188
rect 18163 18134 18209 18186
rect 18209 18134 18219 18186
rect 18243 18134 18273 18186
rect 18273 18134 18285 18186
rect 18285 18134 18299 18186
rect 18323 18134 18337 18186
rect 18337 18134 18349 18186
rect 18349 18134 18379 18186
rect 18403 18134 18413 18186
rect 18413 18134 18459 18186
rect 18163 18132 18219 18134
rect 18243 18132 18299 18134
rect 18323 18132 18379 18134
rect 18403 18132 18459 18134
rect 17503 17642 17559 17644
rect 17583 17642 17639 17644
rect 17663 17642 17719 17644
rect 17743 17642 17799 17644
rect 17503 17590 17549 17642
rect 17549 17590 17559 17642
rect 17583 17590 17613 17642
rect 17613 17590 17625 17642
rect 17625 17590 17639 17642
rect 17663 17590 17677 17642
rect 17677 17590 17689 17642
rect 17689 17590 17719 17642
rect 17743 17590 17753 17642
rect 17753 17590 17799 17642
rect 17503 17588 17559 17590
rect 17583 17588 17639 17590
rect 17663 17588 17719 17590
rect 17743 17588 17799 17590
rect 14345 17098 14401 17100
rect 14425 17098 14481 17100
rect 14505 17098 14561 17100
rect 14585 17098 14641 17100
rect 14345 17046 14391 17098
rect 14391 17046 14401 17098
rect 14425 17046 14455 17098
rect 14455 17046 14467 17098
rect 14467 17046 14481 17098
rect 14505 17046 14519 17098
rect 14519 17046 14531 17098
rect 14531 17046 14561 17098
rect 14585 17046 14595 17098
rect 14595 17046 14641 17098
rect 14345 17044 14401 17046
rect 14425 17044 14481 17046
rect 14505 17044 14561 17046
rect 14585 17044 14641 17046
rect 18163 17098 18219 17100
rect 18243 17098 18299 17100
rect 18323 17098 18379 17100
rect 18403 17098 18459 17100
rect 18163 17046 18209 17098
rect 18209 17046 18219 17098
rect 18243 17046 18273 17098
rect 18273 17046 18285 17098
rect 18285 17046 18299 17098
rect 18323 17046 18337 17098
rect 18337 17046 18349 17098
rect 18349 17046 18379 17098
rect 18403 17046 18413 17098
rect 18413 17046 18459 17098
rect 18163 17044 18219 17046
rect 18243 17044 18299 17046
rect 18323 17044 18379 17046
rect 18403 17044 18459 17046
rect 17503 16554 17559 16556
rect 17583 16554 17639 16556
rect 17663 16554 17719 16556
rect 17743 16554 17799 16556
rect 17503 16502 17549 16554
rect 17549 16502 17559 16554
rect 17583 16502 17613 16554
rect 17613 16502 17625 16554
rect 17625 16502 17639 16554
rect 17663 16502 17677 16554
rect 17677 16502 17689 16554
rect 17689 16502 17719 16554
rect 17743 16502 17753 16554
rect 17753 16502 17799 16554
rect 17503 16500 17559 16502
rect 17583 16500 17639 16502
rect 17663 16500 17719 16502
rect 17743 16500 17799 16502
rect 14345 16010 14401 16012
rect 14425 16010 14481 16012
rect 14505 16010 14561 16012
rect 14585 16010 14641 16012
rect 14345 15958 14391 16010
rect 14391 15958 14401 16010
rect 14425 15958 14455 16010
rect 14455 15958 14467 16010
rect 14467 15958 14481 16010
rect 14505 15958 14519 16010
rect 14519 15958 14531 16010
rect 14531 15958 14561 16010
rect 14585 15958 14595 16010
rect 14595 15958 14641 16010
rect 14345 15956 14401 15958
rect 14425 15956 14481 15958
rect 14505 15956 14561 15958
rect 14585 15956 14641 15958
rect 18163 16010 18219 16012
rect 18243 16010 18299 16012
rect 18323 16010 18379 16012
rect 18403 16010 18459 16012
rect 18163 15958 18209 16010
rect 18209 15958 18219 16010
rect 18243 15958 18273 16010
rect 18273 15958 18285 16010
rect 18285 15958 18299 16010
rect 18323 15958 18337 16010
rect 18337 15958 18349 16010
rect 18349 15958 18379 16010
rect 18403 15958 18413 16010
rect 18413 15958 18459 16010
rect 18163 15956 18219 15958
rect 18243 15956 18299 15958
rect 18323 15956 18379 15958
rect 18403 15956 18459 15958
rect 17503 15466 17559 15468
rect 17583 15466 17639 15468
rect 17663 15466 17719 15468
rect 17743 15466 17799 15468
rect 17503 15414 17549 15466
rect 17549 15414 17559 15466
rect 17583 15414 17613 15466
rect 17613 15414 17625 15466
rect 17625 15414 17639 15466
rect 17663 15414 17677 15466
rect 17677 15414 17689 15466
rect 17689 15414 17719 15466
rect 17743 15414 17753 15466
rect 17753 15414 17799 15466
rect 17503 15412 17559 15414
rect 17583 15412 17639 15414
rect 17663 15412 17719 15414
rect 17743 15412 17799 15414
rect 14345 14922 14401 14924
rect 14425 14922 14481 14924
rect 14505 14922 14561 14924
rect 14585 14922 14641 14924
rect 14345 14870 14391 14922
rect 14391 14870 14401 14922
rect 14425 14870 14455 14922
rect 14455 14870 14467 14922
rect 14467 14870 14481 14922
rect 14505 14870 14519 14922
rect 14519 14870 14531 14922
rect 14531 14870 14561 14922
rect 14585 14870 14595 14922
rect 14595 14870 14641 14922
rect 14345 14868 14401 14870
rect 14425 14868 14481 14870
rect 14505 14868 14561 14870
rect 14585 14868 14641 14870
rect 13685 13290 13741 13292
rect 13765 13290 13821 13292
rect 13845 13290 13901 13292
rect 13925 13290 13981 13292
rect 13685 13238 13731 13290
rect 13731 13238 13741 13290
rect 13765 13238 13795 13290
rect 13795 13238 13807 13290
rect 13807 13238 13821 13290
rect 13845 13238 13859 13290
rect 13859 13238 13871 13290
rect 13871 13238 13901 13290
rect 13925 13238 13935 13290
rect 13935 13238 13981 13290
rect 13685 13236 13741 13238
rect 13765 13236 13821 13238
rect 13845 13236 13901 13238
rect 13925 13236 13981 13238
rect 14345 13834 14401 13836
rect 14425 13834 14481 13836
rect 14505 13834 14561 13836
rect 14585 13834 14641 13836
rect 14345 13782 14391 13834
rect 14391 13782 14401 13834
rect 14425 13782 14455 13834
rect 14455 13782 14467 13834
rect 14467 13782 14481 13834
rect 14505 13782 14519 13834
rect 14519 13782 14531 13834
rect 14531 13782 14561 13834
rect 14585 13782 14595 13834
rect 14595 13782 14641 13834
rect 14345 13780 14401 13782
rect 14425 13780 14481 13782
rect 14505 13780 14561 13782
rect 14585 13780 14641 13782
rect 14345 12746 14401 12748
rect 14425 12746 14481 12748
rect 14505 12746 14561 12748
rect 14585 12746 14641 12748
rect 14345 12694 14391 12746
rect 14391 12694 14401 12746
rect 14425 12694 14455 12746
rect 14455 12694 14467 12746
rect 14467 12694 14481 12746
rect 14505 12694 14519 12746
rect 14519 12694 14531 12746
rect 14531 12694 14561 12746
rect 14585 12694 14595 12746
rect 14595 12694 14641 12746
rect 14345 12692 14401 12694
rect 14425 12692 14481 12694
rect 14505 12692 14561 12694
rect 14585 12692 14641 12694
rect 18163 14922 18219 14924
rect 18243 14922 18299 14924
rect 18323 14922 18379 14924
rect 18403 14922 18459 14924
rect 18163 14870 18209 14922
rect 18209 14870 18219 14922
rect 18243 14870 18273 14922
rect 18273 14870 18285 14922
rect 18285 14870 18299 14922
rect 18323 14870 18337 14922
rect 18337 14870 18349 14922
rect 18349 14870 18379 14922
rect 18403 14870 18413 14922
rect 18413 14870 18459 14922
rect 18163 14868 18219 14870
rect 18243 14868 18299 14870
rect 18323 14868 18379 14870
rect 18403 14868 18459 14870
rect 17503 14378 17559 14380
rect 17583 14378 17639 14380
rect 17663 14378 17719 14380
rect 17743 14378 17799 14380
rect 17503 14326 17549 14378
rect 17549 14326 17559 14378
rect 17583 14326 17613 14378
rect 17613 14326 17625 14378
rect 17625 14326 17639 14378
rect 17663 14326 17677 14378
rect 17677 14326 17689 14378
rect 17689 14326 17719 14378
rect 17743 14326 17753 14378
rect 17753 14326 17799 14378
rect 17503 14324 17559 14326
rect 17583 14324 17639 14326
rect 17663 14324 17719 14326
rect 17743 14324 17799 14326
rect 18163 13834 18219 13836
rect 18243 13834 18299 13836
rect 18323 13834 18379 13836
rect 18403 13834 18459 13836
rect 18163 13782 18209 13834
rect 18209 13782 18219 13834
rect 18243 13782 18273 13834
rect 18273 13782 18285 13834
rect 18285 13782 18299 13834
rect 18323 13782 18337 13834
rect 18337 13782 18349 13834
rect 18349 13782 18379 13834
rect 18403 13782 18413 13834
rect 18413 13782 18459 13834
rect 18163 13780 18219 13782
rect 18243 13780 18299 13782
rect 18323 13780 18379 13782
rect 18403 13780 18459 13782
rect 17503 13290 17559 13292
rect 17583 13290 17639 13292
rect 17663 13290 17719 13292
rect 17743 13290 17799 13292
rect 17503 13238 17549 13290
rect 17549 13238 17559 13290
rect 17583 13238 17613 13290
rect 17613 13238 17625 13290
rect 17625 13238 17639 13290
rect 17663 13238 17677 13290
rect 17677 13238 17689 13290
rect 17689 13238 17719 13290
rect 17743 13238 17753 13290
rect 17753 13238 17799 13290
rect 17503 13236 17559 13238
rect 17583 13236 17639 13238
rect 17663 13236 17719 13238
rect 17743 13236 17799 13238
rect 18163 12746 18219 12748
rect 18243 12746 18299 12748
rect 18323 12746 18379 12748
rect 18403 12746 18459 12748
rect 18163 12694 18209 12746
rect 18209 12694 18219 12746
rect 18243 12694 18273 12746
rect 18273 12694 18285 12746
rect 18285 12694 18299 12746
rect 18323 12694 18337 12746
rect 18337 12694 18349 12746
rect 18349 12694 18379 12746
rect 18403 12694 18413 12746
rect 18413 12694 18459 12746
rect 18163 12692 18219 12694
rect 18243 12692 18299 12694
rect 18323 12692 18379 12694
rect 18403 12692 18459 12694
rect 13685 12202 13741 12204
rect 13765 12202 13821 12204
rect 13845 12202 13901 12204
rect 13925 12202 13981 12204
rect 13685 12150 13731 12202
rect 13731 12150 13741 12202
rect 13765 12150 13795 12202
rect 13795 12150 13807 12202
rect 13807 12150 13821 12202
rect 13845 12150 13859 12202
rect 13859 12150 13871 12202
rect 13871 12150 13901 12202
rect 13925 12150 13935 12202
rect 13935 12150 13981 12202
rect 13685 12148 13741 12150
rect 13765 12148 13821 12150
rect 13845 12148 13901 12150
rect 13925 12148 13981 12150
rect 17503 12202 17559 12204
rect 17583 12202 17639 12204
rect 17663 12202 17719 12204
rect 17743 12202 17799 12204
rect 17503 12150 17549 12202
rect 17549 12150 17559 12202
rect 17583 12150 17613 12202
rect 17613 12150 17625 12202
rect 17625 12150 17639 12202
rect 17663 12150 17677 12202
rect 17677 12150 17689 12202
rect 17689 12150 17719 12202
rect 17743 12150 17753 12202
rect 17753 12150 17799 12202
rect 17503 12148 17559 12150
rect 17583 12148 17639 12150
rect 17663 12148 17719 12150
rect 17743 12148 17799 12150
rect 32070 7320 32220 7330
rect 32070 7190 32080 7320
rect 32080 7190 32220 7320
rect 430 3450 610 3630
rect 1050 3440 1230 3620
rect 440 2510 620 2690
rect 1060 2510 1240 2690
rect 4360 3450 4540 3630
rect 4350 2510 4530 2690
rect 7660 3450 7840 3630
rect 7660 2510 7840 2690
rect 10960 3450 11140 3630
rect 10960 2510 11140 2690
rect 14560 3450 14740 3630
rect 14550 2510 14730 2690
rect 18060 3450 18240 3630
rect 18060 2500 18240 2680
rect 21760 3450 21940 3630
rect 21760 2510 21940 2690
rect 25560 3450 25740 3630
rect 25560 2510 25740 2690
rect 29100 3890 29400 4090
rect 30920 4090 31040 4210
rect 32950 4100 33030 4200
<< metal3 >>
rect 6039 27440 6355 27441
rect 6039 27376 6045 27440
rect 6109 27376 6125 27440
rect 6189 27376 6205 27440
rect 6269 27376 6285 27440
rect 6349 27376 6355 27440
rect 6039 27375 6355 27376
rect 9857 27440 10173 27441
rect 9857 27376 9863 27440
rect 9927 27376 9943 27440
rect 10007 27376 10023 27440
rect 10087 27376 10103 27440
rect 10167 27376 10173 27440
rect 9857 27375 10173 27376
rect 13675 27440 13991 27441
rect 13675 27376 13681 27440
rect 13745 27376 13761 27440
rect 13825 27376 13841 27440
rect 13905 27376 13921 27440
rect 13985 27376 13991 27440
rect 13675 27375 13991 27376
rect 17493 27440 17809 27441
rect 17493 27376 17499 27440
rect 17563 27376 17579 27440
rect 17643 27376 17659 27440
rect 17723 27376 17739 27440
rect 17803 27376 17809 27440
rect 17493 27375 17809 27376
rect 6699 26896 7015 26897
rect 6699 26832 6705 26896
rect 6769 26832 6785 26896
rect 6849 26832 6865 26896
rect 6929 26832 6945 26896
rect 7009 26832 7015 26896
rect 6699 26831 7015 26832
rect 10517 26896 10833 26897
rect 10517 26832 10523 26896
rect 10587 26832 10603 26896
rect 10667 26832 10683 26896
rect 10747 26832 10763 26896
rect 10827 26832 10833 26896
rect 10517 26831 10833 26832
rect 14335 26896 14651 26897
rect 14335 26832 14341 26896
rect 14405 26832 14421 26896
rect 14485 26832 14501 26896
rect 14565 26832 14581 26896
rect 14645 26832 14651 26896
rect 14335 26831 14651 26832
rect 18153 26896 18469 26897
rect 18153 26832 18159 26896
rect 18223 26832 18239 26896
rect 18303 26832 18319 26896
rect 18383 26832 18399 26896
rect 18463 26832 18469 26896
rect 18153 26831 18469 26832
rect 6039 26352 6355 26353
rect 6039 26288 6045 26352
rect 6109 26288 6125 26352
rect 6189 26288 6205 26352
rect 6269 26288 6285 26352
rect 6349 26288 6355 26352
rect 6039 26287 6355 26288
rect 9857 26352 10173 26353
rect 9857 26288 9863 26352
rect 9927 26288 9943 26352
rect 10007 26288 10023 26352
rect 10087 26288 10103 26352
rect 10167 26288 10173 26352
rect 9857 26287 10173 26288
rect 13675 26352 13991 26353
rect 13675 26288 13681 26352
rect 13745 26288 13761 26352
rect 13825 26288 13841 26352
rect 13905 26288 13921 26352
rect 13985 26288 13991 26352
rect 13675 26287 13991 26288
rect 17493 26352 17809 26353
rect 17493 26288 17499 26352
rect 17563 26288 17579 26352
rect 17643 26288 17659 26352
rect 17723 26288 17739 26352
rect 17803 26288 17809 26352
rect 17493 26287 17809 26288
rect 6699 25808 7015 25809
rect 6699 25744 6705 25808
rect 6769 25744 6785 25808
rect 6849 25744 6865 25808
rect 6929 25744 6945 25808
rect 7009 25744 7015 25808
rect 6699 25743 7015 25744
rect 10517 25808 10833 25809
rect 10517 25744 10523 25808
rect 10587 25744 10603 25808
rect 10667 25744 10683 25808
rect 10747 25744 10763 25808
rect 10827 25744 10833 25808
rect 10517 25743 10833 25744
rect 14335 25808 14651 25809
rect 14335 25744 14341 25808
rect 14405 25744 14421 25808
rect 14485 25744 14501 25808
rect 14565 25744 14581 25808
rect 14645 25744 14651 25808
rect 14335 25743 14651 25744
rect 18153 25808 18469 25809
rect 18153 25744 18159 25808
rect 18223 25744 18239 25808
rect 18303 25744 18319 25808
rect 18383 25744 18399 25808
rect 18463 25744 18469 25808
rect 18153 25743 18469 25744
rect 6039 25264 6355 25265
rect 6039 25200 6045 25264
rect 6109 25200 6125 25264
rect 6189 25200 6205 25264
rect 6269 25200 6285 25264
rect 6349 25200 6355 25264
rect 6039 25199 6355 25200
rect 9857 25264 10173 25265
rect 9857 25200 9863 25264
rect 9927 25200 9943 25264
rect 10007 25200 10023 25264
rect 10087 25200 10103 25264
rect 10167 25200 10173 25264
rect 9857 25199 10173 25200
rect 13675 25264 13991 25265
rect 13675 25200 13681 25264
rect 13745 25200 13761 25264
rect 13825 25200 13841 25264
rect 13905 25200 13921 25264
rect 13985 25200 13991 25264
rect 13675 25199 13991 25200
rect 17493 25264 17809 25265
rect 17493 25200 17499 25264
rect 17563 25200 17579 25264
rect 17643 25200 17659 25264
rect 17723 25200 17739 25264
rect 17803 25200 17809 25264
rect 17493 25199 17809 25200
rect 6699 24720 7015 24721
rect 6699 24656 6705 24720
rect 6769 24656 6785 24720
rect 6849 24656 6865 24720
rect 6929 24656 6945 24720
rect 7009 24656 7015 24720
rect 6699 24655 7015 24656
rect 10517 24720 10833 24721
rect 10517 24656 10523 24720
rect 10587 24656 10603 24720
rect 10667 24656 10683 24720
rect 10747 24656 10763 24720
rect 10827 24656 10833 24720
rect 10517 24655 10833 24656
rect 14335 24720 14651 24721
rect 14335 24656 14341 24720
rect 14405 24656 14421 24720
rect 14485 24656 14501 24720
rect 14565 24656 14581 24720
rect 14645 24656 14651 24720
rect 14335 24655 14651 24656
rect 18153 24720 18469 24721
rect 18153 24656 18159 24720
rect 18223 24656 18239 24720
rect 18303 24656 18319 24720
rect 18383 24656 18399 24720
rect 18463 24656 18469 24720
rect 18153 24655 18469 24656
rect 6039 24176 6355 24177
rect 6039 24112 6045 24176
rect 6109 24112 6125 24176
rect 6189 24112 6205 24176
rect 6269 24112 6285 24176
rect 6349 24112 6355 24176
rect 6039 24111 6355 24112
rect 9857 24176 10173 24177
rect 9857 24112 9863 24176
rect 9927 24112 9943 24176
rect 10007 24112 10023 24176
rect 10087 24112 10103 24176
rect 10167 24112 10173 24176
rect 9857 24111 10173 24112
rect 13675 24176 13991 24177
rect 13675 24112 13681 24176
rect 13745 24112 13761 24176
rect 13825 24112 13841 24176
rect 13905 24112 13921 24176
rect 13985 24112 13991 24176
rect 13675 24111 13991 24112
rect 17493 24176 17809 24177
rect 17493 24112 17499 24176
rect 17563 24112 17579 24176
rect 17643 24112 17659 24176
rect 17723 24112 17739 24176
rect 17803 24112 17809 24176
rect 17493 24111 17809 24112
rect 6699 23632 7015 23633
rect 6699 23568 6705 23632
rect 6769 23568 6785 23632
rect 6849 23568 6865 23632
rect 6929 23568 6945 23632
rect 7009 23568 7015 23632
rect 6699 23567 7015 23568
rect 10517 23632 10833 23633
rect 10517 23568 10523 23632
rect 10587 23568 10603 23632
rect 10667 23568 10683 23632
rect 10747 23568 10763 23632
rect 10827 23568 10833 23632
rect 10517 23567 10833 23568
rect 14335 23632 14651 23633
rect 14335 23568 14341 23632
rect 14405 23568 14421 23632
rect 14485 23568 14501 23632
rect 14565 23568 14581 23632
rect 14645 23568 14651 23632
rect 14335 23567 14651 23568
rect 18153 23632 18469 23633
rect 18153 23568 18159 23632
rect 18223 23568 18239 23632
rect 18303 23568 18319 23632
rect 18383 23568 18399 23632
rect 18463 23568 18469 23632
rect 18153 23567 18469 23568
rect 6039 23088 6355 23089
rect 6039 23024 6045 23088
rect 6109 23024 6125 23088
rect 6189 23024 6205 23088
rect 6269 23024 6285 23088
rect 6349 23024 6355 23088
rect 6039 23023 6355 23024
rect 9857 23088 10173 23089
rect 9857 23024 9863 23088
rect 9927 23024 9943 23088
rect 10007 23024 10023 23088
rect 10087 23024 10103 23088
rect 10167 23024 10173 23088
rect 9857 23023 10173 23024
rect 13675 23088 13991 23089
rect 13675 23024 13681 23088
rect 13745 23024 13761 23088
rect 13825 23024 13841 23088
rect 13905 23024 13921 23088
rect 13985 23024 13991 23088
rect 13675 23023 13991 23024
rect 17493 23088 17809 23089
rect 17493 23024 17499 23088
rect 17563 23024 17579 23088
rect 17643 23024 17659 23088
rect 17723 23024 17739 23088
rect 17803 23024 17809 23088
rect 17493 23023 17809 23024
rect 6699 22544 7015 22545
rect 6699 22480 6705 22544
rect 6769 22480 6785 22544
rect 6849 22480 6865 22544
rect 6929 22480 6945 22544
rect 7009 22480 7015 22544
rect 6699 22479 7015 22480
rect 10517 22544 10833 22545
rect 10517 22480 10523 22544
rect 10587 22480 10603 22544
rect 10667 22480 10683 22544
rect 10747 22480 10763 22544
rect 10827 22480 10833 22544
rect 10517 22479 10833 22480
rect 14335 22544 14651 22545
rect 14335 22480 14341 22544
rect 14405 22480 14421 22544
rect 14485 22480 14501 22544
rect 14565 22480 14581 22544
rect 14645 22480 14651 22544
rect 14335 22479 14651 22480
rect 18153 22544 18469 22545
rect 18153 22480 18159 22544
rect 18223 22480 18239 22544
rect 18303 22480 18319 22544
rect 18383 22480 18399 22544
rect 18463 22480 18469 22544
rect 18153 22479 18469 22480
rect 6039 22000 6355 22001
rect 6039 21936 6045 22000
rect 6109 21936 6125 22000
rect 6189 21936 6205 22000
rect 6269 21936 6285 22000
rect 6349 21936 6355 22000
rect 6039 21935 6355 21936
rect 9857 22000 10173 22001
rect 9857 21936 9863 22000
rect 9927 21936 9943 22000
rect 10007 21936 10023 22000
rect 10087 21936 10103 22000
rect 10167 21936 10173 22000
rect 9857 21935 10173 21936
rect 13675 22000 13991 22001
rect 13675 21936 13681 22000
rect 13745 21936 13761 22000
rect 13825 21936 13841 22000
rect 13905 21936 13921 22000
rect 13985 21936 13991 22000
rect 13675 21935 13991 21936
rect 17493 22000 17809 22001
rect 17493 21936 17499 22000
rect 17563 21936 17579 22000
rect 17643 21936 17659 22000
rect 17723 21936 17739 22000
rect 17803 21936 17809 22000
rect 17493 21935 17809 21936
rect 6699 21456 7015 21457
rect 6699 21392 6705 21456
rect 6769 21392 6785 21456
rect 6849 21392 6865 21456
rect 6929 21392 6945 21456
rect 7009 21392 7015 21456
rect 6699 21391 7015 21392
rect 10517 21456 10833 21457
rect 10517 21392 10523 21456
rect 10587 21392 10603 21456
rect 10667 21392 10683 21456
rect 10747 21392 10763 21456
rect 10827 21392 10833 21456
rect 10517 21391 10833 21392
rect 14335 21456 14651 21457
rect 14335 21392 14341 21456
rect 14405 21392 14421 21456
rect 14485 21392 14501 21456
rect 14565 21392 14581 21456
rect 14645 21392 14651 21456
rect 14335 21391 14651 21392
rect 18153 21456 18469 21457
rect 18153 21392 18159 21456
rect 18223 21392 18239 21456
rect 18303 21392 18319 21456
rect 18383 21392 18399 21456
rect 18463 21392 18469 21456
rect 18153 21391 18469 21392
rect 6039 20912 6355 20913
rect 6039 20848 6045 20912
rect 6109 20848 6125 20912
rect 6189 20848 6205 20912
rect 6269 20848 6285 20912
rect 6349 20848 6355 20912
rect 6039 20847 6355 20848
rect 9857 20912 10173 20913
rect 9857 20848 9863 20912
rect 9927 20848 9943 20912
rect 10007 20848 10023 20912
rect 10087 20848 10103 20912
rect 10167 20848 10173 20912
rect 9857 20847 10173 20848
rect 13675 20912 13991 20913
rect 13675 20848 13681 20912
rect 13745 20848 13761 20912
rect 13825 20848 13841 20912
rect 13905 20848 13921 20912
rect 13985 20848 13991 20912
rect 13675 20847 13991 20848
rect 17493 20912 17809 20913
rect 17493 20848 17499 20912
rect 17563 20848 17579 20912
rect 17643 20848 17659 20912
rect 17723 20848 17739 20912
rect 17803 20848 17809 20912
rect 17493 20847 17809 20848
rect 6699 20368 7015 20369
rect 6699 20304 6705 20368
rect 6769 20304 6785 20368
rect 6849 20304 6865 20368
rect 6929 20304 6945 20368
rect 7009 20304 7015 20368
rect 6699 20303 7015 20304
rect 10517 20368 10833 20369
rect 10517 20304 10523 20368
rect 10587 20304 10603 20368
rect 10667 20304 10683 20368
rect 10747 20304 10763 20368
rect 10827 20304 10833 20368
rect 10517 20303 10833 20304
rect 14335 20368 14651 20369
rect 14335 20304 14341 20368
rect 14405 20304 14421 20368
rect 14485 20304 14501 20368
rect 14565 20304 14581 20368
rect 14645 20304 14651 20368
rect 14335 20303 14651 20304
rect 18153 20368 18469 20369
rect 18153 20304 18159 20368
rect 18223 20304 18239 20368
rect 18303 20304 18319 20368
rect 18383 20304 18399 20368
rect 18463 20304 18469 20368
rect 18153 20303 18469 20304
rect 6039 19824 6355 19825
rect 6039 19760 6045 19824
rect 6109 19760 6125 19824
rect 6189 19760 6205 19824
rect 6269 19760 6285 19824
rect 6349 19760 6355 19824
rect 6039 19759 6355 19760
rect 9857 19824 10173 19825
rect 9857 19760 9863 19824
rect 9927 19760 9943 19824
rect 10007 19760 10023 19824
rect 10087 19760 10103 19824
rect 10167 19760 10173 19824
rect 9857 19759 10173 19760
rect 13675 19824 13991 19825
rect 13675 19760 13681 19824
rect 13745 19760 13761 19824
rect 13825 19760 13841 19824
rect 13905 19760 13921 19824
rect 13985 19760 13991 19824
rect 13675 19759 13991 19760
rect 17493 19824 17809 19825
rect 17493 19760 17499 19824
rect 17563 19760 17579 19824
rect 17643 19760 17659 19824
rect 17723 19760 17739 19824
rect 17803 19760 17809 19824
rect 17493 19759 17809 19760
rect 6699 19280 7015 19281
rect 6699 19216 6705 19280
rect 6769 19216 6785 19280
rect 6849 19216 6865 19280
rect 6929 19216 6945 19280
rect 7009 19216 7015 19280
rect 6699 19215 7015 19216
rect 10517 19280 10833 19281
rect 10517 19216 10523 19280
rect 10587 19216 10603 19280
rect 10667 19216 10683 19280
rect 10747 19216 10763 19280
rect 10827 19216 10833 19280
rect 10517 19215 10833 19216
rect 14335 19280 14651 19281
rect 14335 19216 14341 19280
rect 14405 19216 14421 19280
rect 14485 19216 14501 19280
rect 14565 19216 14581 19280
rect 14645 19216 14651 19280
rect 14335 19215 14651 19216
rect 18153 19280 18469 19281
rect 18153 19216 18159 19280
rect 18223 19216 18239 19280
rect 18303 19216 18319 19280
rect 18383 19216 18399 19280
rect 18463 19216 18469 19280
rect 18153 19215 18469 19216
rect 6039 18736 6355 18737
rect 6039 18672 6045 18736
rect 6109 18672 6125 18736
rect 6189 18672 6205 18736
rect 6269 18672 6285 18736
rect 6349 18672 6355 18736
rect 6039 18671 6355 18672
rect 9857 18736 10173 18737
rect 9857 18672 9863 18736
rect 9927 18672 9943 18736
rect 10007 18672 10023 18736
rect 10087 18672 10103 18736
rect 10167 18672 10173 18736
rect 9857 18671 10173 18672
rect 13675 18736 13991 18737
rect 13675 18672 13681 18736
rect 13745 18672 13761 18736
rect 13825 18672 13841 18736
rect 13905 18672 13921 18736
rect 13985 18672 13991 18736
rect 13675 18671 13991 18672
rect 17493 18736 17809 18737
rect 17493 18672 17499 18736
rect 17563 18672 17579 18736
rect 17643 18672 17659 18736
rect 17723 18672 17739 18736
rect 17803 18672 17809 18736
rect 17493 18671 17809 18672
rect 6699 18192 7015 18193
rect 6699 18128 6705 18192
rect 6769 18128 6785 18192
rect 6849 18128 6865 18192
rect 6929 18128 6945 18192
rect 7009 18128 7015 18192
rect 6699 18127 7015 18128
rect 10517 18192 10833 18193
rect 10517 18128 10523 18192
rect 10587 18128 10603 18192
rect 10667 18128 10683 18192
rect 10747 18128 10763 18192
rect 10827 18128 10833 18192
rect 10517 18127 10833 18128
rect 14335 18192 14651 18193
rect 14335 18128 14341 18192
rect 14405 18128 14421 18192
rect 14485 18128 14501 18192
rect 14565 18128 14581 18192
rect 14645 18128 14651 18192
rect 14335 18127 14651 18128
rect 18153 18192 18469 18193
rect 18153 18128 18159 18192
rect 18223 18128 18239 18192
rect 18303 18128 18319 18192
rect 18383 18128 18399 18192
rect 18463 18128 18469 18192
rect 18153 18127 18469 18128
rect 6039 17648 6355 17649
rect 6039 17584 6045 17648
rect 6109 17584 6125 17648
rect 6189 17584 6205 17648
rect 6269 17584 6285 17648
rect 6349 17584 6355 17648
rect 6039 17583 6355 17584
rect 9857 17648 10173 17649
rect 9857 17584 9863 17648
rect 9927 17584 9943 17648
rect 10007 17584 10023 17648
rect 10087 17584 10103 17648
rect 10167 17584 10173 17648
rect 9857 17583 10173 17584
rect 13675 17648 13991 17649
rect 13675 17584 13681 17648
rect 13745 17584 13761 17648
rect 13825 17584 13841 17648
rect 13905 17584 13921 17648
rect 13985 17584 13991 17648
rect 13675 17583 13991 17584
rect 17493 17648 17809 17649
rect 17493 17584 17499 17648
rect 17563 17584 17579 17648
rect 17643 17584 17659 17648
rect 17723 17584 17739 17648
rect 17803 17584 17809 17648
rect 17493 17583 17809 17584
rect 6699 17104 7015 17105
rect 6699 17040 6705 17104
rect 6769 17040 6785 17104
rect 6849 17040 6865 17104
rect 6929 17040 6945 17104
rect 7009 17040 7015 17104
rect 6699 17039 7015 17040
rect 10517 17104 10833 17105
rect 10517 17040 10523 17104
rect 10587 17040 10603 17104
rect 10667 17040 10683 17104
rect 10747 17040 10763 17104
rect 10827 17040 10833 17104
rect 10517 17039 10833 17040
rect 14335 17104 14651 17105
rect 14335 17040 14341 17104
rect 14405 17040 14421 17104
rect 14485 17040 14501 17104
rect 14565 17040 14581 17104
rect 14645 17040 14651 17104
rect 14335 17039 14651 17040
rect 18153 17104 18469 17105
rect 18153 17040 18159 17104
rect 18223 17040 18239 17104
rect 18303 17040 18319 17104
rect 18383 17040 18399 17104
rect 18463 17040 18469 17104
rect 18153 17039 18469 17040
rect 6039 16560 6355 16561
rect 6039 16496 6045 16560
rect 6109 16496 6125 16560
rect 6189 16496 6205 16560
rect 6269 16496 6285 16560
rect 6349 16496 6355 16560
rect 6039 16495 6355 16496
rect 9857 16560 10173 16561
rect 9857 16496 9863 16560
rect 9927 16496 9943 16560
rect 10007 16496 10023 16560
rect 10087 16496 10103 16560
rect 10167 16496 10173 16560
rect 9857 16495 10173 16496
rect 13675 16560 13991 16561
rect 13675 16496 13681 16560
rect 13745 16496 13761 16560
rect 13825 16496 13841 16560
rect 13905 16496 13921 16560
rect 13985 16496 13991 16560
rect 13675 16495 13991 16496
rect 17493 16560 17809 16561
rect 17493 16496 17499 16560
rect 17563 16496 17579 16560
rect 17643 16496 17659 16560
rect 17723 16496 17739 16560
rect 17803 16496 17809 16560
rect 17493 16495 17809 16496
rect 6699 16016 7015 16017
rect 6699 15952 6705 16016
rect 6769 15952 6785 16016
rect 6849 15952 6865 16016
rect 6929 15952 6945 16016
rect 7009 15952 7015 16016
rect 6699 15951 7015 15952
rect 10517 16016 10833 16017
rect 10517 15952 10523 16016
rect 10587 15952 10603 16016
rect 10667 15952 10683 16016
rect 10747 15952 10763 16016
rect 10827 15952 10833 16016
rect 10517 15951 10833 15952
rect 14335 16016 14651 16017
rect 14335 15952 14341 16016
rect 14405 15952 14421 16016
rect 14485 15952 14501 16016
rect 14565 15952 14581 16016
rect 14645 15952 14651 16016
rect 14335 15951 14651 15952
rect 18153 16016 18469 16017
rect 18153 15952 18159 16016
rect 18223 15952 18239 16016
rect 18303 15952 18319 16016
rect 18383 15952 18399 16016
rect 18463 15952 18469 16016
rect 18153 15951 18469 15952
rect 6039 15472 6355 15473
rect 6039 15408 6045 15472
rect 6109 15408 6125 15472
rect 6189 15408 6205 15472
rect 6269 15408 6285 15472
rect 6349 15408 6355 15472
rect 6039 15407 6355 15408
rect 9857 15472 10173 15473
rect 9857 15408 9863 15472
rect 9927 15408 9943 15472
rect 10007 15408 10023 15472
rect 10087 15408 10103 15472
rect 10167 15408 10173 15472
rect 9857 15407 10173 15408
rect 13675 15472 13991 15473
rect 13675 15408 13681 15472
rect 13745 15408 13761 15472
rect 13825 15408 13841 15472
rect 13905 15408 13921 15472
rect 13985 15408 13991 15472
rect 13675 15407 13991 15408
rect 17493 15472 17809 15473
rect 17493 15408 17499 15472
rect 17563 15408 17579 15472
rect 17643 15408 17659 15472
rect 17723 15408 17739 15472
rect 17803 15408 17809 15472
rect 17493 15407 17809 15408
rect 6699 14928 7015 14929
rect 6699 14864 6705 14928
rect 6769 14864 6785 14928
rect 6849 14864 6865 14928
rect 6929 14864 6945 14928
rect 7009 14864 7015 14928
rect 6699 14863 7015 14864
rect 10517 14928 10833 14929
rect 10517 14864 10523 14928
rect 10587 14864 10603 14928
rect 10667 14864 10683 14928
rect 10747 14864 10763 14928
rect 10827 14864 10833 14928
rect 10517 14863 10833 14864
rect 14335 14928 14651 14929
rect 14335 14864 14341 14928
rect 14405 14864 14421 14928
rect 14485 14864 14501 14928
rect 14565 14864 14581 14928
rect 14645 14864 14651 14928
rect 14335 14863 14651 14864
rect 18153 14928 18469 14929
rect 18153 14864 18159 14928
rect 18223 14864 18239 14928
rect 18303 14864 18319 14928
rect 18383 14864 18399 14928
rect 18463 14864 18469 14928
rect 18153 14863 18469 14864
rect 6039 14384 6355 14385
rect 6039 14320 6045 14384
rect 6109 14320 6125 14384
rect 6189 14320 6205 14384
rect 6269 14320 6285 14384
rect 6349 14320 6355 14384
rect 6039 14319 6355 14320
rect 9857 14384 10173 14385
rect 9857 14320 9863 14384
rect 9927 14320 9943 14384
rect 10007 14320 10023 14384
rect 10087 14320 10103 14384
rect 10167 14320 10173 14384
rect 9857 14319 10173 14320
rect 13675 14384 13991 14385
rect 13675 14320 13681 14384
rect 13745 14320 13761 14384
rect 13825 14320 13841 14384
rect 13905 14320 13921 14384
rect 13985 14320 13991 14384
rect 13675 14319 13991 14320
rect 17493 14384 17809 14385
rect 17493 14320 17499 14384
rect 17563 14320 17579 14384
rect 17643 14320 17659 14384
rect 17723 14320 17739 14384
rect 17803 14320 17809 14384
rect 17493 14319 17809 14320
rect 6699 13840 7015 13841
rect 6699 13776 6705 13840
rect 6769 13776 6785 13840
rect 6849 13776 6865 13840
rect 6929 13776 6945 13840
rect 7009 13776 7015 13840
rect 6699 13775 7015 13776
rect 10517 13840 10833 13841
rect 10517 13776 10523 13840
rect 10587 13776 10603 13840
rect 10667 13776 10683 13840
rect 10747 13776 10763 13840
rect 10827 13776 10833 13840
rect 10517 13775 10833 13776
rect 14335 13840 14651 13841
rect 14335 13776 14341 13840
rect 14405 13776 14421 13840
rect 14485 13776 14501 13840
rect 14565 13776 14581 13840
rect 14645 13776 14651 13840
rect 14335 13775 14651 13776
rect 18153 13840 18469 13841
rect 18153 13776 18159 13840
rect 18223 13776 18239 13840
rect 18303 13776 18319 13840
rect 18383 13776 18399 13840
rect 18463 13776 18469 13840
rect 18153 13775 18469 13776
rect 6039 13296 6355 13297
rect 6039 13232 6045 13296
rect 6109 13232 6125 13296
rect 6189 13232 6205 13296
rect 6269 13232 6285 13296
rect 6349 13232 6355 13296
rect 6039 13231 6355 13232
rect 9857 13296 10173 13297
rect 9857 13232 9863 13296
rect 9927 13232 9943 13296
rect 10007 13232 10023 13296
rect 10087 13232 10103 13296
rect 10167 13232 10173 13296
rect 9857 13231 10173 13232
rect 13675 13296 13991 13297
rect 13675 13232 13681 13296
rect 13745 13232 13761 13296
rect 13825 13232 13841 13296
rect 13905 13232 13921 13296
rect 13985 13232 13991 13296
rect 13675 13231 13991 13232
rect 17493 13296 17809 13297
rect 17493 13232 17499 13296
rect 17563 13232 17579 13296
rect 17643 13232 17659 13296
rect 17723 13232 17739 13296
rect 17803 13232 17809 13296
rect 17493 13231 17809 13232
rect 6699 12752 7015 12753
rect 6699 12688 6705 12752
rect 6769 12688 6785 12752
rect 6849 12688 6865 12752
rect 6929 12688 6945 12752
rect 7009 12688 7015 12752
rect 6699 12687 7015 12688
rect 10517 12752 10833 12753
rect 10517 12688 10523 12752
rect 10587 12688 10603 12752
rect 10667 12688 10683 12752
rect 10747 12688 10763 12752
rect 10827 12688 10833 12752
rect 10517 12687 10833 12688
rect 14335 12752 14651 12753
rect 14335 12688 14341 12752
rect 14405 12688 14421 12752
rect 14485 12688 14501 12752
rect 14565 12688 14581 12752
rect 14645 12688 14651 12752
rect 14335 12687 14651 12688
rect 18153 12752 18469 12753
rect 18153 12688 18159 12752
rect 18223 12688 18239 12752
rect 18303 12688 18319 12752
rect 18383 12688 18399 12752
rect 18463 12688 18469 12752
rect 18153 12687 18469 12688
rect 6039 12208 6355 12209
rect 6039 12144 6045 12208
rect 6109 12144 6125 12208
rect 6189 12144 6205 12208
rect 6269 12144 6285 12208
rect 6349 12144 6355 12208
rect 6039 12143 6355 12144
rect 9857 12208 10173 12209
rect 9857 12144 9863 12208
rect 9927 12144 9943 12208
rect 10007 12144 10023 12208
rect 10087 12144 10103 12208
rect 10167 12144 10173 12208
rect 9857 12143 10173 12144
rect 13675 12208 13991 12209
rect 13675 12144 13681 12208
rect 13745 12144 13761 12208
rect 13825 12144 13841 12208
rect 13905 12144 13921 12208
rect 13985 12144 13991 12208
rect 13675 12143 13991 12144
rect 17493 12208 17809 12209
rect 17493 12144 17499 12208
rect 17563 12144 17579 12208
rect 17643 12144 17659 12208
rect 17723 12144 17739 12208
rect 17803 12144 17809 12208
rect 17493 12143 17809 12144
rect 28310 7330 32230 7350
rect 28310 7190 32070 7330
rect 32220 7190 32230 7330
rect 28310 7130 32230 7190
rect 28310 3650 28530 7130
rect 30900 4210 31050 4220
rect 420 3630 28530 3650
rect 420 3450 430 3630
rect 610 3620 4360 3630
rect 610 3450 1050 3620
rect 420 3440 1050 3450
rect 1230 3450 4360 3620
rect 4540 3450 7660 3630
rect 7840 3450 10960 3630
rect 11140 3450 14560 3630
rect 14740 3450 18060 3630
rect 18240 3450 21760 3630
rect 21940 3450 25560 3630
rect 25740 3450 28530 3630
rect 1230 3440 28530 3450
rect 420 3430 28530 3440
rect 29090 4095 29310 4200
rect 29090 4090 29410 4095
rect 29090 3890 29100 4090
rect 29400 3890 29410 4090
rect 30900 4090 30920 4210
rect 31040 4090 31050 4210
rect 32940 4200 33040 4210
rect 32940 4100 32950 4200
rect 33030 4100 33040 4200
rect 32940 4090 33040 4100
rect 30900 4080 31050 4090
rect 29090 3885 29410 3890
rect 29090 2710 29310 3885
rect 430 2690 29310 2710
rect 430 2510 440 2690
rect 620 2510 1060 2690
rect 1240 2510 4350 2690
rect 4530 2510 7660 2690
rect 7840 2510 10960 2690
rect 11140 2510 14550 2690
rect 14730 2680 21760 2690
rect 14730 2510 18060 2680
rect 430 2500 18060 2510
rect 18240 2510 21760 2680
rect 21940 2510 25560 2690
rect 25740 2510 29310 2690
rect 18240 2500 29310 2510
rect 430 2490 29310 2500
rect 29720 3862 34819 3890
rect 29720 918 29740 3862
rect 29804 918 34819 3862
rect 29720 890 34819 918
<< via3 >>
rect 6045 27436 6109 27440
rect 6045 27380 6049 27436
rect 6049 27380 6105 27436
rect 6105 27380 6109 27436
rect 6045 27376 6109 27380
rect 6125 27436 6189 27440
rect 6125 27380 6129 27436
rect 6129 27380 6185 27436
rect 6185 27380 6189 27436
rect 6125 27376 6189 27380
rect 6205 27436 6269 27440
rect 6205 27380 6209 27436
rect 6209 27380 6265 27436
rect 6265 27380 6269 27436
rect 6205 27376 6269 27380
rect 6285 27436 6349 27440
rect 6285 27380 6289 27436
rect 6289 27380 6345 27436
rect 6345 27380 6349 27436
rect 6285 27376 6349 27380
rect 9863 27436 9927 27440
rect 9863 27380 9867 27436
rect 9867 27380 9923 27436
rect 9923 27380 9927 27436
rect 9863 27376 9927 27380
rect 9943 27436 10007 27440
rect 9943 27380 9947 27436
rect 9947 27380 10003 27436
rect 10003 27380 10007 27436
rect 9943 27376 10007 27380
rect 10023 27436 10087 27440
rect 10023 27380 10027 27436
rect 10027 27380 10083 27436
rect 10083 27380 10087 27436
rect 10023 27376 10087 27380
rect 10103 27436 10167 27440
rect 10103 27380 10107 27436
rect 10107 27380 10163 27436
rect 10163 27380 10167 27436
rect 10103 27376 10167 27380
rect 13681 27436 13745 27440
rect 13681 27380 13685 27436
rect 13685 27380 13741 27436
rect 13741 27380 13745 27436
rect 13681 27376 13745 27380
rect 13761 27436 13825 27440
rect 13761 27380 13765 27436
rect 13765 27380 13821 27436
rect 13821 27380 13825 27436
rect 13761 27376 13825 27380
rect 13841 27436 13905 27440
rect 13841 27380 13845 27436
rect 13845 27380 13901 27436
rect 13901 27380 13905 27436
rect 13841 27376 13905 27380
rect 13921 27436 13985 27440
rect 13921 27380 13925 27436
rect 13925 27380 13981 27436
rect 13981 27380 13985 27436
rect 13921 27376 13985 27380
rect 17499 27436 17563 27440
rect 17499 27380 17503 27436
rect 17503 27380 17559 27436
rect 17559 27380 17563 27436
rect 17499 27376 17563 27380
rect 17579 27436 17643 27440
rect 17579 27380 17583 27436
rect 17583 27380 17639 27436
rect 17639 27380 17643 27436
rect 17579 27376 17643 27380
rect 17659 27436 17723 27440
rect 17659 27380 17663 27436
rect 17663 27380 17719 27436
rect 17719 27380 17723 27436
rect 17659 27376 17723 27380
rect 17739 27436 17803 27440
rect 17739 27380 17743 27436
rect 17743 27380 17799 27436
rect 17799 27380 17803 27436
rect 17739 27376 17803 27380
rect 6705 26892 6769 26896
rect 6705 26836 6709 26892
rect 6709 26836 6765 26892
rect 6765 26836 6769 26892
rect 6705 26832 6769 26836
rect 6785 26892 6849 26896
rect 6785 26836 6789 26892
rect 6789 26836 6845 26892
rect 6845 26836 6849 26892
rect 6785 26832 6849 26836
rect 6865 26892 6929 26896
rect 6865 26836 6869 26892
rect 6869 26836 6925 26892
rect 6925 26836 6929 26892
rect 6865 26832 6929 26836
rect 6945 26892 7009 26896
rect 6945 26836 6949 26892
rect 6949 26836 7005 26892
rect 7005 26836 7009 26892
rect 6945 26832 7009 26836
rect 10523 26892 10587 26896
rect 10523 26836 10527 26892
rect 10527 26836 10583 26892
rect 10583 26836 10587 26892
rect 10523 26832 10587 26836
rect 10603 26892 10667 26896
rect 10603 26836 10607 26892
rect 10607 26836 10663 26892
rect 10663 26836 10667 26892
rect 10603 26832 10667 26836
rect 10683 26892 10747 26896
rect 10683 26836 10687 26892
rect 10687 26836 10743 26892
rect 10743 26836 10747 26892
rect 10683 26832 10747 26836
rect 10763 26892 10827 26896
rect 10763 26836 10767 26892
rect 10767 26836 10823 26892
rect 10823 26836 10827 26892
rect 10763 26832 10827 26836
rect 14341 26892 14405 26896
rect 14341 26836 14345 26892
rect 14345 26836 14401 26892
rect 14401 26836 14405 26892
rect 14341 26832 14405 26836
rect 14421 26892 14485 26896
rect 14421 26836 14425 26892
rect 14425 26836 14481 26892
rect 14481 26836 14485 26892
rect 14421 26832 14485 26836
rect 14501 26892 14565 26896
rect 14501 26836 14505 26892
rect 14505 26836 14561 26892
rect 14561 26836 14565 26892
rect 14501 26832 14565 26836
rect 14581 26892 14645 26896
rect 14581 26836 14585 26892
rect 14585 26836 14641 26892
rect 14641 26836 14645 26892
rect 14581 26832 14645 26836
rect 18159 26892 18223 26896
rect 18159 26836 18163 26892
rect 18163 26836 18219 26892
rect 18219 26836 18223 26892
rect 18159 26832 18223 26836
rect 18239 26892 18303 26896
rect 18239 26836 18243 26892
rect 18243 26836 18299 26892
rect 18299 26836 18303 26892
rect 18239 26832 18303 26836
rect 18319 26892 18383 26896
rect 18319 26836 18323 26892
rect 18323 26836 18379 26892
rect 18379 26836 18383 26892
rect 18319 26832 18383 26836
rect 18399 26892 18463 26896
rect 18399 26836 18403 26892
rect 18403 26836 18459 26892
rect 18459 26836 18463 26892
rect 18399 26832 18463 26836
rect 6045 26348 6109 26352
rect 6045 26292 6049 26348
rect 6049 26292 6105 26348
rect 6105 26292 6109 26348
rect 6045 26288 6109 26292
rect 6125 26348 6189 26352
rect 6125 26292 6129 26348
rect 6129 26292 6185 26348
rect 6185 26292 6189 26348
rect 6125 26288 6189 26292
rect 6205 26348 6269 26352
rect 6205 26292 6209 26348
rect 6209 26292 6265 26348
rect 6265 26292 6269 26348
rect 6205 26288 6269 26292
rect 6285 26348 6349 26352
rect 6285 26292 6289 26348
rect 6289 26292 6345 26348
rect 6345 26292 6349 26348
rect 6285 26288 6349 26292
rect 9863 26348 9927 26352
rect 9863 26292 9867 26348
rect 9867 26292 9923 26348
rect 9923 26292 9927 26348
rect 9863 26288 9927 26292
rect 9943 26348 10007 26352
rect 9943 26292 9947 26348
rect 9947 26292 10003 26348
rect 10003 26292 10007 26348
rect 9943 26288 10007 26292
rect 10023 26348 10087 26352
rect 10023 26292 10027 26348
rect 10027 26292 10083 26348
rect 10083 26292 10087 26348
rect 10023 26288 10087 26292
rect 10103 26348 10167 26352
rect 10103 26292 10107 26348
rect 10107 26292 10163 26348
rect 10163 26292 10167 26348
rect 10103 26288 10167 26292
rect 13681 26348 13745 26352
rect 13681 26292 13685 26348
rect 13685 26292 13741 26348
rect 13741 26292 13745 26348
rect 13681 26288 13745 26292
rect 13761 26348 13825 26352
rect 13761 26292 13765 26348
rect 13765 26292 13821 26348
rect 13821 26292 13825 26348
rect 13761 26288 13825 26292
rect 13841 26348 13905 26352
rect 13841 26292 13845 26348
rect 13845 26292 13901 26348
rect 13901 26292 13905 26348
rect 13841 26288 13905 26292
rect 13921 26348 13985 26352
rect 13921 26292 13925 26348
rect 13925 26292 13981 26348
rect 13981 26292 13985 26348
rect 13921 26288 13985 26292
rect 17499 26348 17563 26352
rect 17499 26292 17503 26348
rect 17503 26292 17559 26348
rect 17559 26292 17563 26348
rect 17499 26288 17563 26292
rect 17579 26348 17643 26352
rect 17579 26292 17583 26348
rect 17583 26292 17639 26348
rect 17639 26292 17643 26348
rect 17579 26288 17643 26292
rect 17659 26348 17723 26352
rect 17659 26292 17663 26348
rect 17663 26292 17719 26348
rect 17719 26292 17723 26348
rect 17659 26288 17723 26292
rect 17739 26348 17803 26352
rect 17739 26292 17743 26348
rect 17743 26292 17799 26348
rect 17799 26292 17803 26348
rect 17739 26288 17803 26292
rect 6705 25804 6769 25808
rect 6705 25748 6709 25804
rect 6709 25748 6765 25804
rect 6765 25748 6769 25804
rect 6705 25744 6769 25748
rect 6785 25804 6849 25808
rect 6785 25748 6789 25804
rect 6789 25748 6845 25804
rect 6845 25748 6849 25804
rect 6785 25744 6849 25748
rect 6865 25804 6929 25808
rect 6865 25748 6869 25804
rect 6869 25748 6925 25804
rect 6925 25748 6929 25804
rect 6865 25744 6929 25748
rect 6945 25804 7009 25808
rect 6945 25748 6949 25804
rect 6949 25748 7005 25804
rect 7005 25748 7009 25804
rect 6945 25744 7009 25748
rect 10523 25804 10587 25808
rect 10523 25748 10527 25804
rect 10527 25748 10583 25804
rect 10583 25748 10587 25804
rect 10523 25744 10587 25748
rect 10603 25804 10667 25808
rect 10603 25748 10607 25804
rect 10607 25748 10663 25804
rect 10663 25748 10667 25804
rect 10603 25744 10667 25748
rect 10683 25804 10747 25808
rect 10683 25748 10687 25804
rect 10687 25748 10743 25804
rect 10743 25748 10747 25804
rect 10683 25744 10747 25748
rect 10763 25804 10827 25808
rect 10763 25748 10767 25804
rect 10767 25748 10823 25804
rect 10823 25748 10827 25804
rect 10763 25744 10827 25748
rect 14341 25804 14405 25808
rect 14341 25748 14345 25804
rect 14345 25748 14401 25804
rect 14401 25748 14405 25804
rect 14341 25744 14405 25748
rect 14421 25804 14485 25808
rect 14421 25748 14425 25804
rect 14425 25748 14481 25804
rect 14481 25748 14485 25804
rect 14421 25744 14485 25748
rect 14501 25804 14565 25808
rect 14501 25748 14505 25804
rect 14505 25748 14561 25804
rect 14561 25748 14565 25804
rect 14501 25744 14565 25748
rect 14581 25804 14645 25808
rect 14581 25748 14585 25804
rect 14585 25748 14641 25804
rect 14641 25748 14645 25804
rect 14581 25744 14645 25748
rect 18159 25804 18223 25808
rect 18159 25748 18163 25804
rect 18163 25748 18219 25804
rect 18219 25748 18223 25804
rect 18159 25744 18223 25748
rect 18239 25804 18303 25808
rect 18239 25748 18243 25804
rect 18243 25748 18299 25804
rect 18299 25748 18303 25804
rect 18239 25744 18303 25748
rect 18319 25804 18383 25808
rect 18319 25748 18323 25804
rect 18323 25748 18379 25804
rect 18379 25748 18383 25804
rect 18319 25744 18383 25748
rect 18399 25804 18463 25808
rect 18399 25748 18403 25804
rect 18403 25748 18459 25804
rect 18459 25748 18463 25804
rect 18399 25744 18463 25748
rect 6045 25260 6109 25264
rect 6045 25204 6049 25260
rect 6049 25204 6105 25260
rect 6105 25204 6109 25260
rect 6045 25200 6109 25204
rect 6125 25260 6189 25264
rect 6125 25204 6129 25260
rect 6129 25204 6185 25260
rect 6185 25204 6189 25260
rect 6125 25200 6189 25204
rect 6205 25260 6269 25264
rect 6205 25204 6209 25260
rect 6209 25204 6265 25260
rect 6265 25204 6269 25260
rect 6205 25200 6269 25204
rect 6285 25260 6349 25264
rect 6285 25204 6289 25260
rect 6289 25204 6345 25260
rect 6345 25204 6349 25260
rect 6285 25200 6349 25204
rect 9863 25260 9927 25264
rect 9863 25204 9867 25260
rect 9867 25204 9923 25260
rect 9923 25204 9927 25260
rect 9863 25200 9927 25204
rect 9943 25260 10007 25264
rect 9943 25204 9947 25260
rect 9947 25204 10003 25260
rect 10003 25204 10007 25260
rect 9943 25200 10007 25204
rect 10023 25260 10087 25264
rect 10023 25204 10027 25260
rect 10027 25204 10083 25260
rect 10083 25204 10087 25260
rect 10023 25200 10087 25204
rect 10103 25260 10167 25264
rect 10103 25204 10107 25260
rect 10107 25204 10163 25260
rect 10163 25204 10167 25260
rect 10103 25200 10167 25204
rect 13681 25260 13745 25264
rect 13681 25204 13685 25260
rect 13685 25204 13741 25260
rect 13741 25204 13745 25260
rect 13681 25200 13745 25204
rect 13761 25260 13825 25264
rect 13761 25204 13765 25260
rect 13765 25204 13821 25260
rect 13821 25204 13825 25260
rect 13761 25200 13825 25204
rect 13841 25260 13905 25264
rect 13841 25204 13845 25260
rect 13845 25204 13901 25260
rect 13901 25204 13905 25260
rect 13841 25200 13905 25204
rect 13921 25260 13985 25264
rect 13921 25204 13925 25260
rect 13925 25204 13981 25260
rect 13981 25204 13985 25260
rect 13921 25200 13985 25204
rect 17499 25260 17563 25264
rect 17499 25204 17503 25260
rect 17503 25204 17559 25260
rect 17559 25204 17563 25260
rect 17499 25200 17563 25204
rect 17579 25260 17643 25264
rect 17579 25204 17583 25260
rect 17583 25204 17639 25260
rect 17639 25204 17643 25260
rect 17579 25200 17643 25204
rect 17659 25260 17723 25264
rect 17659 25204 17663 25260
rect 17663 25204 17719 25260
rect 17719 25204 17723 25260
rect 17659 25200 17723 25204
rect 17739 25260 17803 25264
rect 17739 25204 17743 25260
rect 17743 25204 17799 25260
rect 17799 25204 17803 25260
rect 17739 25200 17803 25204
rect 6705 24716 6769 24720
rect 6705 24660 6709 24716
rect 6709 24660 6765 24716
rect 6765 24660 6769 24716
rect 6705 24656 6769 24660
rect 6785 24716 6849 24720
rect 6785 24660 6789 24716
rect 6789 24660 6845 24716
rect 6845 24660 6849 24716
rect 6785 24656 6849 24660
rect 6865 24716 6929 24720
rect 6865 24660 6869 24716
rect 6869 24660 6925 24716
rect 6925 24660 6929 24716
rect 6865 24656 6929 24660
rect 6945 24716 7009 24720
rect 6945 24660 6949 24716
rect 6949 24660 7005 24716
rect 7005 24660 7009 24716
rect 6945 24656 7009 24660
rect 10523 24716 10587 24720
rect 10523 24660 10527 24716
rect 10527 24660 10583 24716
rect 10583 24660 10587 24716
rect 10523 24656 10587 24660
rect 10603 24716 10667 24720
rect 10603 24660 10607 24716
rect 10607 24660 10663 24716
rect 10663 24660 10667 24716
rect 10603 24656 10667 24660
rect 10683 24716 10747 24720
rect 10683 24660 10687 24716
rect 10687 24660 10743 24716
rect 10743 24660 10747 24716
rect 10683 24656 10747 24660
rect 10763 24716 10827 24720
rect 10763 24660 10767 24716
rect 10767 24660 10823 24716
rect 10823 24660 10827 24716
rect 10763 24656 10827 24660
rect 14341 24716 14405 24720
rect 14341 24660 14345 24716
rect 14345 24660 14401 24716
rect 14401 24660 14405 24716
rect 14341 24656 14405 24660
rect 14421 24716 14485 24720
rect 14421 24660 14425 24716
rect 14425 24660 14481 24716
rect 14481 24660 14485 24716
rect 14421 24656 14485 24660
rect 14501 24716 14565 24720
rect 14501 24660 14505 24716
rect 14505 24660 14561 24716
rect 14561 24660 14565 24716
rect 14501 24656 14565 24660
rect 14581 24716 14645 24720
rect 14581 24660 14585 24716
rect 14585 24660 14641 24716
rect 14641 24660 14645 24716
rect 14581 24656 14645 24660
rect 18159 24716 18223 24720
rect 18159 24660 18163 24716
rect 18163 24660 18219 24716
rect 18219 24660 18223 24716
rect 18159 24656 18223 24660
rect 18239 24716 18303 24720
rect 18239 24660 18243 24716
rect 18243 24660 18299 24716
rect 18299 24660 18303 24716
rect 18239 24656 18303 24660
rect 18319 24716 18383 24720
rect 18319 24660 18323 24716
rect 18323 24660 18379 24716
rect 18379 24660 18383 24716
rect 18319 24656 18383 24660
rect 18399 24716 18463 24720
rect 18399 24660 18403 24716
rect 18403 24660 18459 24716
rect 18459 24660 18463 24716
rect 18399 24656 18463 24660
rect 6045 24172 6109 24176
rect 6045 24116 6049 24172
rect 6049 24116 6105 24172
rect 6105 24116 6109 24172
rect 6045 24112 6109 24116
rect 6125 24172 6189 24176
rect 6125 24116 6129 24172
rect 6129 24116 6185 24172
rect 6185 24116 6189 24172
rect 6125 24112 6189 24116
rect 6205 24172 6269 24176
rect 6205 24116 6209 24172
rect 6209 24116 6265 24172
rect 6265 24116 6269 24172
rect 6205 24112 6269 24116
rect 6285 24172 6349 24176
rect 6285 24116 6289 24172
rect 6289 24116 6345 24172
rect 6345 24116 6349 24172
rect 6285 24112 6349 24116
rect 9863 24172 9927 24176
rect 9863 24116 9867 24172
rect 9867 24116 9923 24172
rect 9923 24116 9927 24172
rect 9863 24112 9927 24116
rect 9943 24172 10007 24176
rect 9943 24116 9947 24172
rect 9947 24116 10003 24172
rect 10003 24116 10007 24172
rect 9943 24112 10007 24116
rect 10023 24172 10087 24176
rect 10023 24116 10027 24172
rect 10027 24116 10083 24172
rect 10083 24116 10087 24172
rect 10023 24112 10087 24116
rect 10103 24172 10167 24176
rect 10103 24116 10107 24172
rect 10107 24116 10163 24172
rect 10163 24116 10167 24172
rect 10103 24112 10167 24116
rect 13681 24172 13745 24176
rect 13681 24116 13685 24172
rect 13685 24116 13741 24172
rect 13741 24116 13745 24172
rect 13681 24112 13745 24116
rect 13761 24172 13825 24176
rect 13761 24116 13765 24172
rect 13765 24116 13821 24172
rect 13821 24116 13825 24172
rect 13761 24112 13825 24116
rect 13841 24172 13905 24176
rect 13841 24116 13845 24172
rect 13845 24116 13901 24172
rect 13901 24116 13905 24172
rect 13841 24112 13905 24116
rect 13921 24172 13985 24176
rect 13921 24116 13925 24172
rect 13925 24116 13981 24172
rect 13981 24116 13985 24172
rect 13921 24112 13985 24116
rect 17499 24172 17563 24176
rect 17499 24116 17503 24172
rect 17503 24116 17559 24172
rect 17559 24116 17563 24172
rect 17499 24112 17563 24116
rect 17579 24172 17643 24176
rect 17579 24116 17583 24172
rect 17583 24116 17639 24172
rect 17639 24116 17643 24172
rect 17579 24112 17643 24116
rect 17659 24172 17723 24176
rect 17659 24116 17663 24172
rect 17663 24116 17719 24172
rect 17719 24116 17723 24172
rect 17659 24112 17723 24116
rect 17739 24172 17803 24176
rect 17739 24116 17743 24172
rect 17743 24116 17799 24172
rect 17799 24116 17803 24172
rect 17739 24112 17803 24116
rect 6705 23628 6769 23632
rect 6705 23572 6709 23628
rect 6709 23572 6765 23628
rect 6765 23572 6769 23628
rect 6705 23568 6769 23572
rect 6785 23628 6849 23632
rect 6785 23572 6789 23628
rect 6789 23572 6845 23628
rect 6845 23572 6849 23628
rect 6785 23568 6849 23572
rect 6865 23628 6929 23632
rect 6865 23572 6869 23628
rect 6869 23572 6925 23628
rect 6925 23572 6929 23628
rect 6865 23568 6929 23572
rect 6945 23628 7009 23632
rect 6945 23572 6949 23628
rect 6949 23572 7005 23628
rect 7005 23572 7009 23628
rect 6945 23568 7009 23572
rect 10523 23628 10587 23632
rect 10523 23572 10527 23628
rect 10527 23572 10583 23628
rect 10583 23572 10587 23628
rect 10523 23568 10587 23572
rect 10603 23628 10667 23632
rect 10603 23572 10607 23628
rect 10607 23572 10663 23628
rect 10663 23572 10667 23628
rect 10603 23568 10667 23572
rect 10683 23628 10747 23632
rect 10683 23572 10687 23628
rect 10687 23572 10743 23628
rect 10743 23572 10747 23628
rect 10683 23568 10747 23572
rect 10763 23628 10827 23632
rect 10763 23572 10767 23628
rect 10767 23572 10823 23628
rect 10823 23572 10827 23628
rect 10763 23568 10827 23572
rect 14341 23628 14405 23632
rect 14341 23572 14345 23628
rect 14345 23572 14401 23628
rect 14401 23572 14405 23628
rect 14341 23568 14405 23572
rect 14421 23628 14485 23632
rect 14421 23572 14425 23628
rect 14425 23572 14481 23628
rect 14481 23572 14485 23628
rect 14421 23568 14485 23572
rect 14501 23628 14565 23632
rect 14501 23572 14505 23628
rect 14505 23572 14561 23628
rect 14561 23572 14565 23628
rect 14501 23568 14565 23572
rect 14581 23628 14645 23632
rect 14581 23572 14585 23628
rect 14585 23572 14641 23628
rect 14641 23572 14645 23628
rect 14581 23568 14645 23572
rect 18159 23628 18223 23632
rect 18159 23572 18163 23628
rect 18163 23572 18219 23628
rect 18219 23572 18223 23628
rect 18159 23568 18223 23572
rect 18239 23628 18303 23632
rect 18239 23572 18243 23628
rect 18243 23572 18299 23628
rect 18299 23572 18303 23628
rect 18239 23568 18303 23572
rect 18319 23628 18383 23632
rect 18319 23572 18323 23628
rect 18323 23572 18379 23628
rect 18379 23572 18383 23628
rect 18319 23568 18383 23572
rect 18399 23628 18463 23632
rect 18399 23572 18403 23628
rect 18403 23572 18459 23628
rect 18459 23572 18463 23628
rect 18399 23568 18463 23572
rect 6045 23084 6109 23088
rect 6045 23028 6049 23084
rect 6049 23028 6105 23084
rect 6105 23028 6109 23084
rect 6045 23024 6109 23028
rect 6125 23084 6189 23088
rect 6125 23028 6129 23084
rect 6129 23028 6185 23084
rect 6185 23028 6189 23084
rect 6125 23024 6189 23028
rect 6205 23084 6269 23088
rect 6205 23028 6209 23084
rect 6209 23028 6265 23084
rect 6265 23028 6269 23084
rect 6205 23024 6269 23028
rect 6285 23084 6349 23088
rect 6285 23028 6289 23084
rect 6289 23028 6345 23084
rect 6345 23028 6349 23084
rect 6285 23024 6349 23028
rect 9863 23084 9927 23088
rect 9863 23028 9867 23084
rect 9867 23028 9923 23084
rect 9923 23028 9927 23084
rect 9863 23024 9927 23028
rect 9943 23084 10007 23088
rect 9943 23028 9947 23084
rect 9947 23028 10003 23084
rect 10003 23028 10007 23084
rect 9943 23024 10007 23028
rect 10023 23084 10087 23088
rect 10023 23028 10027 23084
rect 10027 23028 10083 23084
rect 10083 23028 10087 23084
rect 10023 23024 10087 23028
rect 10103 23084 10167 23088
rect 10103 23028 10107 23084
rect 10107 23028 10163 23084
rect 10163 23028 10167 23084
rect 10103 23024 10167 23028
rect 13681 23084 13745 23088
rect 13681 23028 13685 23084
rect 13685 23028 13741 23084
rect 13741 23028 13745 23084
rect 13681 23024 13745 23028
rect 13761 23084 13825 23088
rect 13761 23028 13765 23084
rect 13765 23028 13821 23084
rect 13821 23028 13825 23084
rect 13761 23024 13825 23028
rect 13841 23084 13905 23088
rect 13841 23028 13845 23084
rect 13845 23028 13901 23084
rect 13901 23028 13905 23084
rect 13841 23024 13905 23028
rect 13921 23084 13985 23088
rect 13921 23028 13925 23084
rect 13925 23028 13981 23084
rect 13981 23028 13985 23084
rect 13921 23024 13985 23028
rect 17499 23084 17563 23088
rect 17499 23028 17503 23084
rect 17503 23028 17559 23084
rect 17559 23028 17563 23084
rect 17499 23024 17563 23028
rect 17579 23084 17643 23088
rect 17579 23028 17583 23084
rect 17583 23028 17639 23084
rect 17639 23028 17643 23084
rect 17579 23024 17643 23028
rect 17659 23084 17723 23088
rect 17659 23028 17663 23084
rect 17663 23028 17719 23084
rect 17719 23028 17723 23084
rect 17659 23024 17723 23028
rect 17739 23084 17803 23088
rect 17739 23028 17743 23084
rect 17743 23028 17799 23084
rect 17799 23028 17803 23084
rect 17739 23024 17803 23028
rect 6705 22540 6769 22544
rect 6705 22484 6709 22540
rect 6709 22484 6765 22540
rect 6765 22484 6769 22540
rect 6705 22480 6769 22484
rect 6785 22540 6849 22544
rect 6785 22484 6789 22540
rect 6789 22484 6845 22540
rect 6845 22484 6849 22540
rect 6785 22480 6849 22484
rect 6865 22540 6929 22544
rect 6865 22484 6869 22540
rect 6869 22484 6925 22540
rect 6925 22484 6929 22540
rect 6865 22480 6929 22484
rect 6945 22540 7009 22544
rect 6945 22484 6949 22540
rect 6949 22484 7005 22540
rect 7005 22484 7009 22540
rect 6945 22480 7009 22484
rect 10523 22540 10587 22544
rect 10523 22484 10527 22540
rect 10527 22484 10583 22540
rect 10583 22484 10587 22540
rect 10523 22480 10587 22484
rect 10603 22540 10667 22544
rect 10603 22484 10607 22540
rect 10607 22484 10663 22540
rect 10663 22484 10667 22540
rect 10603 22480 10667 22484
rect 10683 22540 10747 22544
rect 10683 22484 10687 22540
rect 10687 22484 10743 22540
rect 10743 22484 10747 22540
rect 10683 22480 10747 22484
rect 10763 22540 10827 22544
rect 10763 22484 10767 22540
rect 10767 22484 10823 22540
rect 10823 22484 10827 22540
rect 10763 22480 10827 22484
rect 14341 22540 14405 22544
rect 14341 22484 14345 22540
rect 14345 22484 14401 22540
rect 14401 22484 14405 22540
rect 14341 22480 14405 22484
rect 14421 22540 14485 22544
rect 14421 22484 14425 22540
rect 14425 22484 14481 22540
rect 14481 22484 14485 22540
rect 14421 22480 14485 22484
rect 14501 22540 14565 22544
rect 14501 22484 14505 22540
rect 14505 22484 14561 22540
rect 14561 22484 14565 22540
rect 14501 22480 14565 22484
rect 14581 22540 14645 22544
rect 14581 22484 14585 22540
rect 14585 22484 14641 22540
rect 14641 22484 14645 22540
rect 14581 22480 14645 22484
rect 18159 22540 18223 22544
rect 18159 22484 18163 22540
rect 18163 22484 18219 22540
rect 18219 22484 18223 22540
rect 18159 22480 18223 22484
rect 18239 22540 18303 22544
rect 18239 22484 18243 22540
rect 18243 22484 18299 22540
rect 18299 22484 18303 22540
rect 18239 22480 18303 22484
rect 18319 22540 18383 22544
rect 18319 22484 18323 22540
rect 18323 22484 18379 22540
rect 18379 22484 18383 22540
rect 18319 22480 18383 22484
rect 18399 22540 18463 22544
rect 18399 22484 18403 22540
rect 18403 22484 18459 22540
rect 18459 22484 18463 22540
rect 18399 22480 18463 22484
rect 6045 21996 6109 22000
rect 6045 21940 6049 21996
rect 6049 21940 6105 21996
rect 6105 21940 6109 21996
rect 6045 21936 6109 21940
rect 6125 21996 6189 22000
rect 6125 21940 6129 21996
rect 6129 21940 6185 21996
rect 6185 21940 6189 21996
rect 6125 21936 6189 21940
rect 6205 21996 6269 22000
rect 6205 21940 6209 21996
rect 6209 21940 6265 21996
rect 6265 21940 6269 21996
rect 6205 21936 6269 21940
rect 6285 21996 6349 22000
rect 6285 21940 6289 21996
rect 6289 21940 6345 21996
rect 6345 21940 6349 21996
rect 6285 21936 6349 21940
rect 9863 21996 9927 22000
rect 9863 21940 9867 21996
rect 9867 21940 9923 21996
rect 9923 21940 9927 21996
rect 9863 21936 9927 21940
rect 9943 21996 10007 22000
rect 9943 21940 9947 21996
rect 9947 21940 10003 21996
rect 10003 21940 10007 21996
rect 9943 21936 10007 21940
rect 10023 21996 10087 22000
rect 10023 21940 10027 21996
rect 10027 21940 10083 21996
rect 10083 21940 10087 21996
rect 10023 21936 10087 21940
rect 10103 21996 10167 22000
rect 10103 21940 10107 21996
rect 10107 21940 10163 21996
rect 10163 21940 10167 21996
rect 10103 21936 10167 21940
rect 13681 21996 13745 22000
rect 13681 21940 13685 21996
rect 13685 21940 13741 21996
rect 13741 21940 13745 21996
rect 13681 21936 13745 21940
rect 13761 21996 13825 22000
rect 13761 21940 13765 21996
rect 13765 21940 13821 21996
rect 13821 21940 13825 21996
rect 13761 21936 13825 21940
rect 13841 21996 13905 22000
rect 13841 21940 13845 21996
rect 13845 21940 13901 21996
rect 13901 21940 13905 21996
rect 13841 21936 13905 21940
rect 13921 21996 13985 22000
rect 13921 21940 13925 21996
rect 13925 21940 13981 21996
rect 13981 21940 13985 21996
rect 13921 21936 13985 21940
rect 17499 21996 17563 22000
rect 17499 21940 17503 21996
rect 17503 21940 17559 21996
rect 17559 21940 17563 21996
rect 17499 21936 17563 21940
rect 17579 21996 17643 22000
rect 17579 21940 17583 21996
rect 17583 21940 17639 21996
rect 17639 21940 17643 21996
rect 17579 21936 17643 21940
rect 17659 21996 17723 22000
rect 17659 21940 17663 21996
rect 17663 21940 17719 21996
rect 17719 21940 17723 21996
rect 17659 21936 17723 21940
rect 17739 21996 17803 22000
rect 17739 21940 17743 21996
rect 17743 21940 17799 21996
rect 17799 21940 17803 21996
rect 17739 21936 17803 21940
rect 6705 21452 6769 21456
rect 6705 21396 6709 21452
rect 6709 21396 6765 21452
rect 6765 21396 6769 21452
rect 6705 21392 6769 21396
rect 6785 21452 6849 21456
rect 6785 21396 6789 21452
rect 6789 21396 6845 21452
rect 6845 21396 6849 21452
rect 6785 21392 6849 21396
rect 6865 21452 6929 21456
rect 6865 21396 6869 21452
rect 6869 21396 6925 21452
rect 6925 21396 6929 21452
rect 6865 21392 6929 21396
rect 6945 21452 7009 21456
rect 6945 21396 6949 21452
rect 6949 21396 7005 21452
rect 7005 21396 7009 21452
rect 6945 21392 7009 21396
rect 10523 21452 10587 21456
rect 10523 21396 10527 21452
rect 10527 21396 10583 21452
rect 10583 21396 10587 21452
rect 10523 21392 10587 21396
rect 10603 21452 10667 21456
rect 10603 21396 10607 21452
rect 10607 21396 10663 21452
rect 10663 21396 10667 21452
rect 10603 21392 10667 21396
rect 10683 21452 10747 21456
rect 10683 21396 10687 21452
rect 10687 21396 10743 21452
rect 10743 21396 10747 21452
rect 10683 21392 10747 21396
rect 10763 21452 10827 21456
rect 10763 21396 10767 21452
rect 10767 21396 10823 21452
rect 10823 21396 10827 21452
rect 10763 21392 10827 21396
rect 14341 21452 14405 21456
rect 14341 21396 14345 21452
rect 14345 21396 14401 21452
rect 14401 21396 14405 21452
rect 14341 21392 14405 21396
rect 14421 21452 14485 21456
rect 14421 21396 14425 21452
rect 14425 21396 14481 21452
rect 14481 21396 14485 21452
rect 14421 21392 14485 21396
rect 14501 21452 14565 21456
rect 14501 21396 14505 21452
rect 14505 21396 14561 21452
rect 14561 21396 14565 21452
rect 14501 21392 14565 21396
rect 14581 21452 14645 21456
rect 14581 21396 14585 21452
rect 14585 21396 14641 21452
rect 14641 21396 14645 21452
rect 14581 21392 14645 21396
rect 18159 21452 18223 21456
rect 18159 21396 18163 21452
rect 18163 21396 18219 21452
rect 18219 21396 18223 21452
rect 18159 21392 18223 21396
rect 18239 21452 18303 21456
rect 18239 21396 18243 21452
rect 18243 21396 18299 21452
rect 18299 21396 18303 21452
rect 18239 21392 18303 21396
rect 18319 21452 18383 21456
rect 18319 21396 18323 21452
rect 18323 21396 18379 21452
rect 18379 21396 18383 21452
rect 18319 21392 18383 21396
rect 18399 21452 18463 21456
rect 18399 21396 18403 21452
rect 18403 21396 18459 21452
rect 18459 21396 18463 21452
rect 18399 21392 18463 21396
rect 6045 20908 6109 20912
rect 6045 20852 6049 20908
rect 6049 20852 6105 20908
rect 6105 20852 6109 20908
rect 6045 20848 6109 20852
rect 6125 20908 6189 20912
rect 6125 20852 6129 20908
rect 6129 20852 6185 20908
rect 6185 20852 6189 20908
rect 6125 20848 6189 20852
rect 6205 20908 6269 20912
rect 6205 20852 6209 20908
rect 6209 20852 6265 20908
rect 6265 20852 6269 20908
rect 6205 20848 6269 20852
rect 6285 20908 6349 20912
rect 6285 20852 6289 20908
rect 6289 20852 6345 20908
rect 6345 20852 6349 20908
rect 6285 20848 6349 20852
rect 9863 20908 9927 20912
rect 9863 20852 9867 20908
rect 9867 20852 9923 20908
rect 9923 20852 9927 20908
rect 9863 20848 9927 20852
rect 9943 20908 10007 20912
rect 9943 20852 9947 20908
rect 9947 20852 10003 20908
rect 10003 20852 10007 20908
rect 9943 20848 10007 20852
rect 10023 20908 10087 20912
rect 10023 20852 10027 20908
rect 10027 20852 10083 20908
rect 10083 20852 10087 20908
rect 10023 20848 10087 20852
rect 10103 20908 10167 20912
rect 10103 20852 10107 20908
rect 10107 20852 10163 20908
rect 10163 20852 10167 20908
rect 10103 20848 10167 20852
rect 13681 20908 13745 20912
rect 13681 20852 13685 20908
rect 13685 20852 13741 20908
rect 13741 20852 13745 20908
rect 13681 20848 13745 20852
rect 13761 20908 13825 20912
rect 13761 20852 13765 20908
rect 13765 20852 13821 20908
rect 13821 20852 13825 20908
rect 13761 20848 13825 20852
rect 13841 20908 13905 20912
rect 13841 20852 13845 20908
rect 13845 20852 13901 20908
rect 13901 20852 13905 20908
rect 13841 20848 13905 20852
rect 13921 20908 13985 20912
rect 13921 20852 13925 20908
rect 13925 20852 13981 20908
rect 13981 20852 13985 20908
rect 13921 20848 13985 20852
rect 17499 20908 17563 20912
rect 17499 20852 17503 20908
rect 17503 20852 17559 20908
rect 17559 20852 17563 20908
rect 17499 20848 17563 20852
rect 17579 20908 17643 20912
rect 17579 20852 17583 20908
rect 17583 20852 17639 20908
rect 17639 20852 17643 20908
rect 17579 20848 17643 20852
rect 17659 20908 17723 20912
rect 17659 20852 17663 20908
rect 17663 20852 17719 20908
rect 17719 20852 17723 20908
rect 17659 20848 17723 20852
rect 17739 20908 17803 20912
rect 17739 20852 17743 20908
rect 17743 20852 17799 20908
rect 17799 20852 17803 20908
rect 17739 20848 17803 20852
rect 6705 20364 6769 20368
rect 6705 20308 6709 20364
rect 6709 20308 6765 20364
rect 6765 20308 6769 20364
rect 6705 20304 6769 20308
rect 6785 20364 6849 20368
rect 6785 20308 6789 20364
rect 6789 20308 6845 20364
rect 6845 20308 6849 20364
rect 6785 20304 6849 20308
rect 6865 20364 6929 20368
rect 6865 20308 6869 20364
rect 6869 20308 6925 20364
rect 6925 20308 6929 20364
rect 6865 20304 6929 20308
rect 6945 20364 7009 20368
rect 6945 20308 6949 20364
rect 6949 20308 7005 20364
rect 7005 20308 7009 20364
rect 6945 20304 7009 20308
rect 10523 20364 10587 20368
rect 10523 20308 10527 20364
rect 10527 20308 10583 20364
rect 10583 20308 10587 20364
rect 10523 20304 10587 20308
rect 10603 20364 10667 20368
rect 10603 20308 10607 20364
rect 10607 20308 10663 20364
rect 10663 20308 10667 20364
rect 10603 20304 10667 20308
rect 10683 20364 10747 20368
rect 10683 20308 10687 20364
rect 10687 20308 10743 20364
rect 10743 20308 10747 20364
rect 10683 20304 10747 20308
rect 10763 20364 10827 20368
rect 10763 20308 10767 20364
rect 10767 20308 10823 20364
rect 10823 20308 10827 20364
rect 10763 20304 10827 20308
rect 14341 20364 14405 20368
rect 14341 20308 14345 20364
rect 14345 20308 14401 20364
rect 14401 20308 14405 20364
rect 14341 20304 14405 20308
rect 14421 20364 14485 20368
rect 14421 20308 14425 20364
rect 14425 20308 14481 20364
rect 14481 20308 14485 20364
rect 14421 20304 14485 20308
rect 14501 20364 14565 20368
rect 14501 20308 14505 20364
rect 14505 20308 14561 20364
rect 14561 20308 14565 20364
rect 14501 20304 14565 20308
rect 14581 20364 14645 20368
rect 14581 20308 14585 20364
rect 14585 20308 14641 20364
rect 14641 20308 14645 20364
rect 14581 20304 14645 20308
rect 18159 20364 18223 20368
rect 18159 20308 18163 20364
rect 18163 20308 18219 20364
rect 18219 20308 18223 20364
rect 18159 20304 18223 20308
rect 18239 20364 18303 20368
rect 18239 20308 18243 20364
rect 18243 20308 18299 20364
rect 18299 20308 18303 20364
rect 18239 20304 18303 20308
rect 18319 20364 18383 20368
rect 18319 20308 18323 20364
rect 18323 20308 18379 20364
rect 18379 20308 18383 20364
rect 18319 20304 18383 20308
rect 18399 20364 18463 20368
rect 18399 20308 18403 20364
rect 18403 20308 18459 20364
rect 18459 20308 18463 20364
rect 18399 20304 18463 20308
rect 6045 19820 6109 19824
rect 6045 19764 6049 19820
rect 6049 19764 6105 19820
rect 6105 19764 6109 19820
rect 6045 19760 6109 19764
rect 6125 19820 6189 19824
rect 6125 19764 6129 19820
rect 6129 19764 6185 19820
rect 6185 19764 6189 19820
rect 6125 19760 6189 19764
rect 6205 19820 6269 19824
rect 6205 19764 6209 19820
rect 6209 19764 6265 19820
rect 6265 19764 6269 19820
rect 6205 19760 6269 19764
rect 6285 19820 6349 19824
rect 6285 19764 6289 19820
rect 6289 19764 6345 19820
rect 6345 19764 6349 19820
rect 6285 19760 6349 19764
rect 9863 19820 9927 19824
rect 9863 19764 9867 19820
rect 9867 19764 9923 19820
rect 9923 19764 9927 19820
rect 9863 19760 9927 19764
rect 9943 19820 10007 19824
rect 9943 19764 9947 19820
rect 9947 19764 10003 19820
rect 10003 19764 10007 19820
rect 9943 19760 10007 19764
rect 10023 19820 10087 19824
rect 10023 19764 10027 19820
rect 10027 19764 10083 19820
rect 10083 19764 10087 19820
rect 10023 19760 10087 19764
rect 10103 19820 10167 19824
rect 10103 19764 10107 19820
rect 10107 19764 10163 19820
rect 10163 19764 10167 19820
rect 10103 19760 10167 19764
rect 13681 19820 13745 19824
rect 13681 19764 13685 19820
rect 13685 19764 13741 19820
rect 13741 19764 13745 19820
rect 13681 19760 13745 19764
rect 13761 19820 13825 19824
rect 13761 19764 13765 19820
rect 13765 19764 13821 19820
rect 13821 19764 13825 19820
rect 13761 19760 13825 19764
rect 13841 19820 13905 19824
rect 13841 19764 13845 19820
rect 13845 19764 13901 19820
rect 13901 19764 13905 19820
rect 13841 19760 13905 19764
rect 13921 19820 13985 19824
rect 13921 19764 13925 19820
rect 13925 19764 13981 19820
rect 13981 19764 13985 19820
rect 13921 19760 13985 19764
rect 17499 19820 17563 19824
rect 17499 19764 17503 19820
rect 17503 19764 17559 19820
rect 17559 19764 17563 19820
rect 17499 19760 17563 19764
rect 17579 19820 17643 19824
rect 17579 19764 17583 19820
rect 17583 19764 17639 19820
rect 17639 19764 17643 19820
rect 17579 19760 17643 19764
rect 17659 19820 17723 19824
rect 17659 19764 17663 19820
rect 17663 19764 17719 19820
rect 17719 19764 17723 19820
rect 17659 19760 17723 19764
rect 17739 19820 17803 19824
rect 17739 19764 17743 19820
rect 17743 19764 17799 19820
rect 17799 19764 17803 19820
rect 17739 19760 17803 19764
rect 6705 19276 6769 19280
rect 6705 19220 6709 19276
rect 6709 19220 6765 19276
rect 6765 19220 6769 19276
rect 6705 19216 6769 19220
rect 6785 19276 6849 19280
rect 6785 19220 6789 19276
rect 6789 19220 6845 19276
rect 6845 19220 6849 19276
rect 6785 19216 6849 19220
rect 6865 19276 6929 19280
rect 6865 19220 6869 19276
rect 6869 19220 6925 19276
rect 6925 19220 6929 19276
rect 6865 19216 6929 19220
rect 6945 19276 7009 19280
rect 6945 19220 6949 19276
rect 6949 19220 7005 19276
rect 7005 19220 7009 19276
rect 6945 19216 7009 19220
rect 10523 19276 10587 19280
rect 10523 19220 10527 19276
rect 10527 19220 10583 19276
rect 10583 19220 10587 19276
rect 10523 19216 10587 19220
rect 10603 19276 10667 19280
rect 10603 19220 10607 19276
rect 10607 19220 10663 19276
rect 10663 19220 10667 19276
rect 10603 19216 10667 19220
rect 10683 19276 10747 19280
rect 10683 19220 10687 19276
rect 10687 19220 10743 19276
rect 10743 19220 10747 19276
rect 10683 19216 10747 19220
rect 10763 19276 10827 19280
rect 10763 19220 10767 19276
rect 10767 19220 10823 19276
rect 10823 19220 10827 19276
rect 10763 19216 10827 19220
rect 14341 19276 14405 19280
rect 14341 19220 14345 19276
rect 14345 19220 14401 19276
rect 14401 19220 14405 19276
rect 14341 19216 14405 19220
rect 14421 19276 14485 19280
rect 14421 19220 14425 19276
rect 14425 19220 14481 19276
rect 14481 19220 14485 19276
rect 14421 19216 14485 19220
rect 14501 19276 14565 19280
rect 14501 19220 14505 19276
rect 14505 19220 14561 19276
rect 14561 19220 14565 19276
rect 14501 19216 14565 19220
rect 14581 19276 14645 19280
rect 14581 19220 14585 19276
rect 14585 19220 14641 19276
rect 14641 19220 14645 19276
rect 14581 19216 14645 19220
rect 18159 19276 18223 19280
rect 18159 19220 18163 19276
rect 18163 19220 18219 19276
rect 18219 19220 18223 19276
rect 18159 19216 18223 19220
rect 18239 19276 18303 19280
rect 18239 19220 18243 19276
rect 18243 19220 18299 19276
rect 18299 19220 18303 19276
rect 18239 19216 18303 19220
rect 18319 19276 18383 19280
rect 18319 19220 18323 19276
rect 18323 19220 18379 19276
rect 18379 19220 18383 19276
rect 18319 19216 18383 19220
rect 18399 19276 18463 19280
rect 18399 19220 18403 19276
rect 18403 19220 18459 19276
rect 18459 19220 18463 19276
rect 18399 19216 18463 19220
rect 6045 18732 6109 18736
rect 6045 18676 6049 18732
rect 6049 18676 6105 18732
rect 6105 18676 6109 18732
rect 6045 18672 6109 18676
rect 6125 18732 6189 18736
rect 6125 18676 6129 18732
rect 6129 18676 6185 18732
rect 6185 18676 6189 18732
rect 6125 18672 6189 18676
rect 6205 18732 6269 18736
rect 6205 18676 6209 18732
rect 6209 18676 6265 18732
rect 6265 18676 6269 18732
rect 6205 18672 6269 18676
rect 6285 18732 6349 18736
rect 6285 18676 6289 18732
rect 6289 18676 6345 18732
rect 6345 18676 6349 18732
rect 6285 18672 6349 18676
rect 9863 18732 9927 18736
rect 9863 18676 9867 18732
rect 9867 18676 9923 18732
rect 9923 18676 9927 18732
rect 9863 18672 9927 18676
rect 9943 18732 10007 18736
rect 9943 18676 9947 18732
rect 9947 18676 10003 18732
rect 10003 18676 10007 18732
rect 9943 18672 10007 18676
rect 10023 18732 10087 18736
rect 10023 18676 10027 18732
rect 10027 18676 10083 18732
rect 10083 18676 10087 18732
rect 10023 18672 10087 18676
rect 10103 18732 10167 18736
rect 10103 18676 10107 18732
rect 10107 18676 10163 18732
rect 10163 18676 10167 18732
rect 10103 18672 10167 18676
rect 13681 18732 13745 18736
rect 13681 18676 13685 18732
rect 13685 18676 13741 18732
rect 13741 18676 13745 18732
rect 13681 18672 13745 18676
rect 13761 18732 13825 18736
rect 13761 18676 13765 18732
rect 13765 18676 13821 18732
rect 13821 18676 13825 18732
rect 13761 18672 13825 18676
rect 13841 18732 13905 18736
rect 13841 18676 13845 18732
rect 13845 18676 13901 18732
rect 13901 18676 13905 18732
rect 13841 18672 13905 18676
rect 13921 18732 13985 18736
rect 13921 18676 13925 18732
rect 13925 18676 13981 18732
rect 13981 18676 13985 18732
rect 13921 18672 13985 18676
rect 17499 18732 17563 18736
rect 17499 18676 17503 18732
rect 17503 18676 17559 18732
rect 17559 18676 17563 18732
rect 17499 18672 17563 18676
rect 17579 18732 17643 18736
rect 17579 18676 17583 18732
rect 17583 18676 17639 18732
rect 17639 18676 17643 18732
rect 17579 18672 17643 18676
rect 17659 18732 17723 18736
rect 17659 18676 17663 18732
rect 17663 18676 17719 18732
rect 17719 18676 17723 18732
rect 17659 18672 17723 18676
rect 17739 18732 17803 18736
rect 17739 18676 17743 18732
rect 17743 18676 17799 18732
rect 17799 18676 17803 18732
rect 17739 18672 17803 18676
rect 6705 18188 6769 18192
rect 6705 18132 6709 18188
rect 6709 18132 6765 18188
rect 6765 18132 6769 18188
rect 6705 18128 6769 18132
rect 6785 18188 6849 18192
rect 6785 18132 6789 18188
rect 6789 18132 6845 18188
rect 6845 18132 6849 18188
rect 6785 18128 6849 18132
rect 6865 18188 6929 18192
rect 6865 18132 6869 18188
rect 6869 18132 6925 18188
rect 6925 18132 6929 18188
rect 6865 18128 6929 18132
rect 6945 18188 7009 18192
rect 6945 18132 6949 18188
rect 6949 18132 7005 18188
rect 7005 18132 7009 18188
rect 6945 18128 7009 18132
rect 10523 18188 10587 18192
rect 10523 18132 10527 18188
rect 10527 18132 10583 18188
rect 10583 18132 10587 18188
rect 10523 18128 10587 18132
rect 10603 18188 10667 18192
rect 10603 18132 10607 18188
rect 10607 18132 10663 18188
rect 10663 18132 10667 18188
rect 10603 18128 10667 18132
rect 10683 18188 10747 18192
rect 10683 18132 10687 18188
rect 10687 18132 10743 18188
rect 10743 18132 10747 18188
rect 10683 18128 10747 18132
rect 10763 18188 10827 18192
rect 10763 18132 10767 18188
rect 10767 18132 10823 18188
rect 10823 18132 10827 18188
rect 10763 18128 10827 18132
rect 14341 18188 14405 18192
rect 14341 18132 14345 18188
rect 14345 18132 14401 18188
rect 14401 18132 14405 18188
rect 14341 18128 14405 18132
rect 14421 18188 14485 18192
rect 14421 18132 14425 18188
rect 14425 18132 14481 18188
rect 14481 18132 14485 18188
rect 14421 18128 14485 18132
rect 14501 18188 14565 18192
rect 14501 18132 14505 18188
rect 14505 18132 14561 18188
rect 14561 18132 14565 18188
rect 14501 18128 14565 18132
rect 14581 18188 14645 18192
rect 14581 18132 14585 18188
rect 14585 18132 14641 18188
rect 14641 18132 14645 18188
rect 14581 18128 14645 18132
rect 18159 18188 18223 18192
rect 18159 18132 18163 18188
rect 18163 18132 18219 18188
rect 18219 18132 18223 18188
rect 18159 18128 18223 18132
rect 18239 18188 18303 18192
rect 18239 18132 18243 18188
rect 18243 18132 18299 18188
rect 18299 18132 18303 18188
rect 18239 18128 18303 18132
rect 18319 18188 18383 18192
rect 18319 18132 18323 18188
rect 18323 18132 18379 18188
rect 18379 18132 18383 18188
rect 18319 18128 18383 18132
rect 18399 18188 18463 18192
rect 18399 18132 18403 18188
rect 18403 18132 18459 18188
rect 18459 18132 18463 18188
rect 18399 18128 18463 18132
rect 6045 17644 6109 17648
rect 6045 17588 6049 17644
rect 6049 17588 6105 17644
rect 6105 17588 6109 17644
rect 6045 17584 6109 17588
rect 6125 17644 6189 17648
rect 6125 17588 6129 17644
rect 6129 17588 6185 17644
rect 6185 17588 6189 17644
rect 6125 17584 6189 17588
rect 6205 17644 6269 17648
rect 6205 17588 6209 17644
rect 6209 17588 6265 17644
rect 6265 17588 6269 17644
rect 6205 17584 6269 17588
rect 6285 17644 6349 17648
rect 6285 17588 6289 17644
rect 6289 17588 6345 17644
rect 6345 17588 6349 17644
rect 6285 17584 6349 17588
rect 9863 17644 9927 17648
rect 9863 17588 9867 17644
rect 9867 17588 9923 17644
rect 9923 17588 9927 17644
rect 9863 17584 9927 17588
rect 9943 17644 10007 17648
rect 9943 17588 9947 17644
rect 9947 17588 10003 17644
rect 10003 17588 10007 17644
rect 9943 17584 10007 17588
rect 10023 17644 10087 17648
rect 10023 17588 10027 17644
rect 10027 17588 10083 17644
rect 10083 17588 10087 17644
rect 10023 17584 10087 17588
rect 10103 17644 10167 17648
rect 10103 17588 10107 17644
rect 10107 17588 10163 17644
rect 10163 17588 10167 17644
rect 10103 17584 10167 17588
rect 13681 17644 13745 17648
rect 13681 17588 13685 17644
rect 13685 17588 13741 17644
rect 13741 17588 13745 17644
rect 13681 17584 13745 17588
rect 13761 17644 13825 17648
rect 13761 17588 13765 17644
rect 13765 17588 13821 17644
rect 13821 17588 13825 17644
rect 13761 17584 13825 17588
rect 13841 17644 13905 17648
rect 13841 17588 13845 17644
rect 13845 17588 13901 17644
rect 13901 17588 13905 17644
rect 13841 17584 13905 17588
rect 13921 17644 13985 17648
rect 13921 17588 13925 17644
rect 13925 17588 13981 17644
rect 13981 17588 13985 17644
rect 13921 17584 13985 17588
rect 17499 17644 17563 17648
rect 17499 17588 17503 17644
rect 17503 17588 17559 17644
rect 17559 17588 17563 17644
rect 17499 17584 17563 17588
rect 17579 17644 17643 17648
rect 17579 17588 17583 17644
rect 17583 17588 17639 17644
rect 17639 17588 17643 17644
rect 17579 17584 17643 17588
rect 17659 17644 17723 17648
rect 17659 17588 17663 17644
rect 17663 17588 17719 17644
rect 17719 17588 17723 17644
rect 17659 17584 17723 17588
rect 17739 17644 17803 17648
rect 17739 17588 17743 17644
rect 17743 17588 17799 17644
rect 17799 17588 17803 17644
rect 17739 17584 17803 17588
rect 6705 17100 6769 17104
rect 6705 17044 6709 17100
rect 6709 17044 6765 17100
rect 6765 17044 6769 17100
rect 6705 17040 6769 17044
rect 6785 17100 6849 17104
rect 6785 17044 6789 17100
rect 6789 17044 6845 17100
rect 6845 17044 6849 17100
rect 6785 17040 6849 17044
rect 6865 17100 6929 17104
rect 6865 17044 6869 17100
rect 6869 17044 6925 17100
rect 6925 17044 6929 17100
rect 6865 17040 6929 17044
rect 6945 17100 7009 17104
rect 6945 17044 6949 17100
rect 6949 17044 7005 17100
rect 7005 17044 7009 17100
rect 6945 17040 7009 17044
rect 10523 17100 10587 17104
rect 10523 17044 10527 17100
rect 10527 17044 10583 17100
rect 10583 17044 10587 17100
rect 10523 17040 10587 17044
rect 10603 17100 10667 17104
rect 10603 17044 10607 17100
rect 10607 17044 10663 17100
rect 10663 17044 10667 17100
rect 10603 17040 10667 17044
rect 10683 17100 10747 17104
rect 10683 17044 10687 17100
rect 10687 17044 10743 17100
rect 10743 17044 10747 17100
rect 10683 17040 10747 17044
rect 10763 17100 10827 17104
rect 10763 17044 10767 17100
rect 10767 17044 10823 17100
rect 10823 17044 10827 17100
rect 10763 17040 10827 17044
rect 14341 17100 14405 17104
rect 14341 17044 14345 17100
rect 14345 17044 14401 17100
rect 14401 17044 14405 17100
rect 14341 17040 14405 17044
rect 14421 17100 14485 17104
rect 14421 17044 14425 17100
rect 14425 17044 14481 17100
rect 14481 17044 14485 17100
rect 14421 17040 14485 17044
rect 14501 17100 14565 17104
rect 14501 17044 14505 17100
rect 14505 17044 14561 17100
rect 14561 17044 14565 17100
rect 14501 17040 14565 17044
rect 14581 17100 14645 17104
rect 14581 17044 14585 17100
rect 14585 17044 14641 17100
rect 14641 17044 14645 17100
rect 14581 17040 14645 17044
rect 18159 17100 18223 17104
rect 18159 17044 18163 17100
rect 18163 17044 18219 17100
rect 18219 17044 18223 17100
rect 18159 17040 18223 17044
rect 18239 17100 18303 17104
rect 18239 17044 18243 17100
rect 18243 17044 18299 17100
rect 18299 17044 18303 17100
rect 18239 17040 18303 17044
rect 18319 17100 18383 17104
rect 18319 17044 18323 17100
rect 18323 17044 18379 17100
rect 18379 17044 18383 17100
rect 18319 17040 18383 17044
rect 18399 17100 18463 17104
rect 18399 17044 18403 17100
rect 18403 17044 18459 17100
rect 18459 17044 18463 17100
rect 18399 17040 18463 17044
rect 6045 16556 6109 16560
rect 6045 16500 6049 16556
rect 6049 16500 6105 16556
rect 6105 16500 6109 16556
rect 6045 16496 6109 16500
rect 6125 16556 6189 16560
rect 6125 16500 6129 16556
rect 6129 16500 6185 16556
rect 6185 16500 6189 16556
rect 6125 16496 6189 16500
rect 6205 16556 6269 16560
rect 6205 16500 6209 16556
rect 6209 16500 6265 16556
rect 6265 16500 6269 16556
rect 6205 16496 6269 16500
rect 6285 16556 6349 16560
rect 6285 16500 6289 16556
rect 6289 16500 6345 16556
rect 6345 16500 6349 16556
rect 6285 16496 6349 16500
rect 9863 16556 9927 16560
rect 9863 16500 9867 16556
rect 9867 16500 9923 16556
rect 9923 16500 9927 16556
rect 9863 16496 9927 16500
rect 9943 16556 10007 16560
rect 9943 16500 9947 16556
rect 9947 16500 10003 16556
rect 10003 16500 10007 16556
rect 9943 16496 10007 16500
rect 10023 16556 10087 16560
rect 10023 16500 10027 16556
rect 10027 16500 10083 16556
rect 10083 16500 10087 16556
rect 10023 16496 10087 16500
rect 10103 16556 10167 16560
rect 10103 16500 10107 16556
rect 10107 16500 10163 16556
rect 10163 16500 10167 16556
rect 10103 16496 10167 16500
rect 13681 16556 13745 16560
rect 13681 16500 13685 16556
rect 13685 16500 13741 16556
rect 13741 16500 13745 16556
rect 13681 16496 13745 16500
rect 13761 16556 13825 16560
rect 13761 16500 13765 16556
rect 13765 16500 13821 16556
rect 13821 16500 13825 16556
rect 13761 16496 13825 16500
rect 13841 16556 13905 16560
rect 13841 16500 13845 16556
rect 13845 16500 13901 16556
rect 13901 16500 13905 16556
rect 13841 16496 13905 16500
rect 13921 16556 13985 16560
rect 13921 16500 13925 16556
rect 13925 16500 13981 16556
rect 13981 16500 13985 16556
rect 13921 16496 13985 16500
rect 17499 16556 17563 16560
rect 17499 16500 17503 16556
rect 17503 16500 17559 16556
rect 17559 16500 17563 16556
rect 17499 16496 17563 16500
rect 17579 16556 17643 16560
rect 17579 16500 17583 16556
rect 17583 16500 17639 16556
rect 17639 16500 17643 16556
rect 17579 16496 17643 16500
rect 17659 16556 17723 16560
rect 17659 16500 17663 16556
rect 17663 16500 17719 16556
rect 17719 16500 17723 16556
rect 17659 16496 17723 16500
rect 17739 16556 17803 16560
rect 17739 16500 17743 16556
rect 17743 16500 17799 16556
rect 17799 16500 17803 16556
rect 17739 16496 17803 16500
rect 6705 16012 6769 16016
rect 6705 15956 6709 16012
rect 6709 15956 6765 16012
rect 6765 15956 6769 16012
rect 6705 15952 6769 15956
rect 6785 16012 6849 16016
rect 6785 15956 6789 16012
rect 6789 15956 6845 16012
rect 6845 15956 6849 16012
rect 6785 15952 6849 15956
rect 6865 16012 6929 16016
rect 6865 15956 6869 16012
rect 6869 15956 6925 16012
rect 6925 15956 6929 16012
rect 6865 15952 6929 15956
rect 6945 16012 7009 16016
rect 6945 15956 6949 16012
rect 6949 15956 7005 16012
rect 7005 15956 7009 16012
rect 6945 15952 7009 15956
rect 10523 16012 10587 16016
rect 10523 15956 10527 16012
rect 10527 15956 10583 16012
rect 10583 15956 10587 16012
rect 10523 15952 10587 15956
rect 10603 16012 10667 16016
rect 10603 15956 10607 16012
rect 10607 15956 10663 16012
rect 10663 15956 10667 16012
rect 10603 15952 10667 15956
rect 10683 16012 10747 16016
rect 10683 15956 10687 16012
rect 10687 15956 10743 16012
rect 10743 15956 10747 16012
rect 10683 15952 10747 15956
rect 10763 16012 10827 16016
rect 10763 15956 10767 16012
rect 10767 15956 10823 16012
rect 10823 15956 10827 16012
rect 10763 15952 10827 15956
rect 14341 16012 14405 16016
rect 14341 15956 14345 16012
rect 14345 15956 14401 16012
rect 14401 15956 14405 16012
rect 14341 15952 14405 15956
rect 14421 16012 14485 16016
rect 14421 15956 14425 16012
rect 14425 15956 14481 16012
rect 14481 15956 14485 16012
rect 14421 15952 14485 15956
rect 14501 16012 14565 16016
rect 14501 15956 14505 16012
rect 14505 15956 14561 16012
rect 14561 15956 14565 16012
rect 14501 15952 14565 15956
rect 14581 16012 14645 16016
rect 14581 15956 14585 16012
rect 14585 15956 14641 16012
rect 14641 15956 14645 16012
rect 14581 15952 14645 15956
rect 18159 16012 18223 16016
rect 18159 15956 18163 16012
rect 18163 15956 18219 16012
rect 18219 15956 18223 16012
rect 18159 15952 18223 15956
rect 18239 16012 18303 16016
rect 18239 15956 18243 16012
rect 18243 15956 18299 16012
rect 18299 15956 18303 16012
rect 18239 15952 18303 15956
rect 18319 16012 18383 16016
rect 18319 15956 18323 16012
rect 18323 15956 18379 16012
rect 18379 15956 18383 16012
rect 18319 15952 18383 15956
rect 18399 16012 18463 16016
rect 18399 15956 18403 16012
rect 18403 15956 18459 16012
rect 18459 15956 18463 16012
rect 18399 15952 18463 15956
rect 6045 15468 6109 15472
rect 6045 15412 6049 15468
rect 6049 15412 6105 15468
rect 6105 15412 6109 15468
rect 6045 15408 6109 15412
rect 6125 15468 6189 15472
rect 6125 15412 6129 15468
rect 6129 15412 6185 15468
rect 6185 15412 6189 15468
rect 6125 15408 6189 15412
rect 6205 15468 6269 15472
rect 6205 15412 6209 15468
rect 6209 15412 6265 15468
rect 6265 15412 6269 15468
rect 6205 15408 6269 15412
rect 6285 15468 6349 15472
rect 6285 15412 6289 15468
rect 6289 15412 6345 15468
rect 6345 15412 6349 15468
rect 6285 15408 6349 15412
rect 9863 15468 9927 15472
rect 9863 15412 9867 15468
rect 9867 15412 9923 15468
rect 9923 15412 9927 15468
rect 9863 15408 9927 15412
rect 9943 15468 10007 15472
rect 9943 15412 9947 15468
rect 9947 15412 10003 15468
rect 10003 15412 10007 15468
rect 9943 15408 10007 15412
rect 10023 15468 10087 15472
rect 10023 15412 10027 15468
rect 10027 15412 10083 15468
rect 10083 15412 10087 15468
rect 10023 15408 10087 15412
rect 10103 15468 10167 15472
rect 10103 15412 10107 15468
rect 10107 15412 10163 15468
rect 10163 15412 10167 15468
rect 10103 15408 10167 15412
rect 13681 15468 13745 15472
rect 13681 15412 13685 15468
rect 13685 15412 13741 15468
rect 13741 15412 13745 15468
rect 13681 15408 13745 15412
rect 13761 15468 13825 15472
rect 13761 15412 13765 15468
rect 13765 15412 13821 15468
rect 13821 15412 13825 15468
rect 13761 15408 13825 15412
rect 13841 15468 13905 15472
rect 13841 15412 13845 15468
rect 13845 15412 13901 15468
rect 13901 15412 13905 15468
rect 13841 15408 13905 15412
rect 13921 15468 13985 15472
rect 13921 15412 13925 15468
rect 13925 15412 13981 15468
rect 13981 15412 13985 15468
rect 13921 15408 13985 15412
rect 17499 15468 17563 15472
rect 17499 15412 17503 15468
rect 17503 15412 17559 15468
rect 17559 15412 17563 15468
rect 17499 15408 17563 15412
rect 17579 15468 17643 15472
rect 17579 15412 17583 15468
rect 17583 15412 17639 15468
rect 17639 15412 17643 15468
rect 17579 15408 17643 15412
rect 17659 15468 17723 15472
rect 17659 15412 17663 15468
rect 17663 15412 17719 15468
rect 17719 15412 17723 15468
rect 17659 15408 17723 15412
rect 17739 15468 17803 15472
rect 17739 15412 17743 15468
rect 17743 15412 17799 15468
rect 17799 15412 17803 15468
rect 17739 15408 17803 15412
rect 6705 14924 6769 14928
rect 6705 14868 6709 14924
rect 6709 14868 6765 14924
rect 6765 14868 6769 14924
rect 6705 14864 6769 14868
rect 6785 14924 6849 14928
rect 6785 14868 6789 14924
rect 6789 14868 6845 14924
rect 6845 14868 6849 14924
rect 6785 14864 6849 14868
rect 6865 14924 6929 14928
rect 6865 14868 6869 14924
rect 6869 14868 6925 14924
rect 6925 14868 6929 14924
rect 6865 14864 6929 14868
rect 6945 14924 7009 14928
rect 6945 14868 6949 14924
rect 6949 14868 7005 14924
rect 7005 14868 7009 14924
rect 6945 14864 7009 14868
rect 10523 14924 10587 14928
rect 10523 14868 10527 14924
rect 10527 14868 10583 14924
rect 10583 14868 10587 14924
rect 10523 14864 10587 14868
rect 10603 14924 10667 14928
rect 10603 14868 10607 14924
rect 10607 14868 10663 14924
rect 10663 14868 10667 14924
rect 10603 14864 10667 14868
rect 10683 14924 10747 14928
rect 10683 14868 10687 14924
rect 10687 14868 10743 14924
rect 10743 14868 10747 14924
rect 10683 14864 10747 14868
rect 10763 14924 10827 14928
rect 10763 14868 10767 14924
rect 10767 14868 10823 14924
rect 10823 14868 10827 14924
rect 10763 14864 10827 14868
rect 14341 14924 14405 14928
rect 14341 14868 14345 14924
rect 14345 14868 14401 14924
rect 14401 14868 14405 14924
rect 14341 14864 14405 14868
rect 14421 14924 14485 14928
rect 14421 14868 14425 14924
rect 14425 14868 14481 14924
rect 14481 14868 14485 14924
rect 14421 14864 14485 14868
rect 14501 14924 14565 14928
rect 14501 14868 14505 14924
rect 14505 14868 14561 14924
rect 14561 14868 14565 14924
rect 14501 14864 14565 14868
rect 14581 14924 14645 14928
rect 14581 14868 14585 14924
rect 14585 14868 14641 14924
rect 14641 14868 14645 14924
rect 14581 14864 14645 14868
rect 18159 14924 18223 14928
rect 18159 14868 18163 14924
rect 18163 14868 18219 14924
rect 18219 14868 18223 14924
rect 18159 14864 18223 14868
rect 18239 14924 18303 14928
rect 18239 14868 18243 14924
rect 18243 14868 18299 14924
rect 18299 14868 18303 14924
rect 18239 14864 18303 14868
rect 18319 14924 18383 14928
rect 18319 14868 18323 14924
rect 18323 14868 18379 14924
rect 18379 14868 18383 14924
rect 18319 14864 18383 14868
rect 18399 14924 18463 14928
rect 18399 14868 18403 14924
rect 18403 14868 18459 14924
rect 18459 14868 18463 14924
rect 18399 14864 18463 14868
rect 6045 14380 6109 14384
rect 6045 14324 6049 14380
rect 6049 14324 6105 14380
rect 6105 14324 6109 14380
rect 6045 14320 6109 14324
rect 6125 14380 6189 14384
rect 6125 14324 6129 14380
rect 6129 14324 6185 14380
rect 6185 14324 6189 14380
rect 6125 14320 6189 14324
rect 6205 14380 6269 14384
rect 6205 14324 6209 14380
rect 6209 14324 6265 14380
rect 6265 14324 6269 14380
rect 6205 14320 6269 14324
rect 6285 14380 6349 14384
rect 6285 14324 6289 14380
rect 6289 14324 6345 14380
rect 6345 14324 6349 14380
rect 6285 14320 6349 14324
rect 9863 14380 9927 14384
rect 9863 14324 9867 14380
rect 9867 14324 9923 14380
rect 9923 14324 9927 14380
rect 9863 14320 9927 14324
rect 9943 14380 10007 14384
rect 9943 14324 9947 14380
rect 9947 14324 10003 14380
rect 10003 14324 10007 14380
rect 9943 14320 10007 14324
rect 10023 14380 10087 14384
rect 10023 14324 10027 14380
rect 10027 14324 10083 14380
rect 10083 14324 10087 14380
rect 10023 14320 10087 14324
rect 10103 14380 10167 14384
rect 10103 14324 10107 14380
rect 10107 14324 10163 14380
rect 10163 14324 10167 14380
rect 10103 14320 10167 14324
rect 13681 14380 13745 14384
rect 13681 14324 13685 14380
rect 13685 14324 13741 14380
rect 13741 14324 13745 14380
rect 13681 14320 13745 14324
rect 13761 14380 13825 14384
rect 13761 14324 13765 14380
rect 13765 14324 13821 14380
rect 13821 14324 13825 14380
rect 13761 14320 13825 14324
rect 13841 14380 13905 14384
rect 13841 14324 13845 14380
rect 13845 14324 13901 14380
rect 13901 14324 13905 14380
rect 13841 14320 13905 14324
rect 13921 14380 13985 14384
rect 13921 14324 13925 14380
rect 13925 14324 13981 14380
rect 13981 14324 13985 14380
rect 13921 14320 13985 14324
rect 17499 14380 17563 14384
rect 17499 14324 17503 14380
rect 17503 14324 17559 14380
rect 17559 14324 17563 14380
rect 17499 14320 17563 14324
rect 17579 14380 17643 14384
rect 17579 14324 17583 14380
rect 17583 14324 17639 14380
rect 17639 14324 17643 14380
rect 17579 14320 17643 14324
rect 17659 14380 17723 14384
rect 17659 14324 17663 14380
rect 17663 14324 17719 14380
rect 17719 14324 17723 14380
rect 17659 14320 17723 14324
rect 17739 14380 17803 14384
rect 17739 14324 17743 14380
rect 17743 14324 17799 14380
rect 17799 14324 17803 14380
rect 17739 14320 17803 14324
rect 6705 13836 6769 13840
rect 6705 13780 6709 13836
rect 6709 13780 6765 13836
rect 6765 13780 6769 13836
rect 6705 13776 6769 13780
rect 6785 13836 6849 13840
rect 6785 13780 6789 13836
rect 6789 13780 6845 13836
rect 6845 13780 6849 13836
rect 6785 13776 6849 13780
rect 6865 13836 6929 13840
rect 6865 13780 6869 13836
rect 6869 13780 6925 13836
rect 6925 13780 6929 13836
rect 6865 13776 6929 13780
rect 6945 13836 7009 13840
rect 6945 13780 6949 13836
rect 6949 13780 7005 13836
rect 7005 13780 7009 13836
rect 6945 13776 7009 13780
rect 10523 13836 10587 13840
rect 10523 13780 10527 13836
rect 10527 13780 10583 13836
rect 10583 13780 10587 13836
rect 10523 13776 10587 13780
rect 10603 13836 10667 13840
rect 10603 13780 10607 13836
rect 10607 13780 10663 13836
rect 10663 13780 10667 13836
rect 10603 13776 10667 13780
rect 10683 13836 10747 13840
rect 10683 13780 10687 13836
rect 10687 13780 10743 13836
rect 10743 13780 10747 13836
rect 10683 13776 10747 13780
rect 10763 13836 10827 13840
rect 10763 13780 10767 13836
rect 10767 13780 10823 13836
rect 10823 13780 10827 13836
rect 10763 13776 10827 13780
rect 14341 13836 14405 13840
rect 14341 13780 14345 13836
rect 14345 13780 14401 13836
rect 14401 13780 14405 13836
rect 14341 13776 14405 13780
rect 14421 13836 14485 13840
rect 14421 13780 14425 13836
rect 14425 13780 14481 13836
rect 14481 13780 14485 13836
rect 14421 13776 14485 13780
rect 14501 13836 14565 13840
rect 14501 13780 14505 13836
rect 14505 13780 14561 13836
rect 14561 13780 14565 13836
rect 14501 13776 14565 13780
rect 14581 13836 14645 13840
rect 14581 13780 14585 13836
rect 14585 13780 14641 13836
rect 14641 13780 14645 13836
rect 14581 13776 14645 13780
rect 18159 13836 18223 13840
rect 18159 13780 18163 13836
rect 18163 13780 18219 13836
rect 18219 13780 18223 13836
rect 18159 13776 18223 13780
rect 18239 13836 18303 13840
rect 18239 13780 18243 13836
rect 18243 13780 18299 13836
rect 18299 13780 18303 13836
rect 18239 13776 18303 13780
rect 18319 13836 18383 13840
rect 18319 13780 18323 13836
rect 18323 13780 18379 13836
rect 18379 13780 18383 13836
rect 18319 13776 18383 13780
rect 18399 13836 18463 13840
rect 18399 13780 18403 13836
rect 18403 13780 18459 13836
rect 18459 13780 18463 13836
rect 18399 13776 18463 13780
rect 6045 13292 6109 13296
rect 6045 13236 6049 13292
rect 6049 13236 6105 13292
rect 6105 13236 6109 13292
rect 6045 13232 6109 13236
rect 6125 13292 6189 13296
rect 6125 13236 6129 13292
rect 6129 13236 6185 13292
rect 6185 13236 6189 13292
rect 6125 13232 6189 13236
rect 6205 13292 6269 13296
rect 6205 13236 6209 13292
rect 6209 13236 6265 13292
rect 6265 13236 6269 13292
rect 6205 13232 6269 13236
rect 6285 13292 6349 13296
rect 6285 13236 6289 13292
rect 6289 13236 6345 13292
rect 6345 13236 6349 13292
rect 6285 13232 6349 13236
rect 9863 13292 9927 13296
rect 9863 13236 9867 13292
rect 9867 13236 9923 13292
rect 9923 13236 9927 13292
rect 9863 13232 9927 13236
rect 9943 13292 10007 13296
rect 9943 13236 9947 13292
rect 9947 13236 10003 13292
rect 10003 13236 10007 13292
rect 9943 13232 10007 13236
rect 10023 13292 10087 13296
rect 10023 13236 10027 13292
rect 10027 13236 10083 13292
rect 10083 13236 10087 13292
rect 10023 13232 10087 13236
rect 10103 13292 10167 13296
rect 10103 13236 10107 13292
rect 10107 13236 10163 13292
rect 10163 13236 10167 13292
rect 10103 13232 10167 13236
rect 13681 13292 13745 13296
rect 13681 13236 13685 13292
rect 13685 13236 13741 13292
rect 13741 13236 13745 13292
rect 13681 13232 13745 13236
rect 13761 13292 13825 13296
rect 13761 13236 13765 13292
rect 13765 13236 13821 13292
rect 13821 13236 13825 13292
rect 13761 13232 13825 13236
rect 13841 13292 13905 13296
rect 13841 13236 13845 13292
rect 13845 13236 13901 13292
rect 13901 13236 13905 13292
rect 13841 13232 13905 13236
rect 13921 13292 13985 13296
rect 13921 13236 13925 13292
rect 13925 13236 13981 13292
rect 13981 13236 13985 13292
rect 13921 13232 13985 13236
rect 17499 13292 17563 13296
rect 17499 13236 17503 13292
rect 17503 13236 17559 13292
rect 17559 13236 17563 13292
rect 17499 13232 17563 13236
rect 17579 13292 17643 13296
rect 17579 13236 17583 13292
rect 17583 13236 17639 13292
rect 17639 13236 17643 13292
rect 17579 13232 17643 13236
rect 17659 13292 17723 13296
rect 17659 13236 17663 13292
rect 17663 13236 17719 13292
rect 17719 13236 17723 13292
rect 17659 13232 17723 13236
rect 17739 13292 17803 13296
rect 17739 13236 17743 13292
rect 17743 13236 17799 13292
rect 17799 13236 17803 13292
rect 17739 13232 17803 13236
rect 6705 12748 6769 12752
rect 6705 12692 6709 12748
rect 6709 12692 6765 12748
rect 6765 12692 6769 12748
rect 6705 12688 6769 12692
rect 6785 12748 6849 12752
rect 6785 12692 6789 12748
rect 6789 12692 6845 12748
rect 6845 12692 6849 12748
rect 6785 12688 6849 12692
rect 6865 12748 6929 12752
rect 6865 12692 6869 12748
rect 6869 12692 6925 12748
rect 6925 12692 6929 12748
rect 6865 12688 6929 12692
rect 6945 12748 7009 12752
rect 6945 12692 6949 12748
rect 6949 12692 7005 12748
rect 7005 12692 7009 12748
rect 6945 12688 7009 12692
rect 10523 12748 10587 12752
rect 10523 12692 10527 12748
rect 10527 12692 10583 12748
rect 10583 12692 10587 12748
rect 10523 12688 10587 12692
rect 10603 12748 10667 12752
rect 10603 12692 10607 12748
rect 10607 12692 10663 12748
rect 10663 12692 10667 12748
rect 10603 12688 10667 12692
rect 10683 12748 10747 12752
rect 10683 12692 10687 12748
rect 10687 12692 10743 12748
rect 10743 12692 10747 12748
rect 10683 12688 10747 12692
rect 10763 12748 10827 12752
rect 10763 12692 10767 12748
rect 10767 12692 10823 12748
rect 10823 12692 10827 12748
rect 10763 12688 10827 12692
rect 14341 12748 14405 12752
rect 14341 12692 14345 12748
rect 14345 12692 14401 12748
rect 14401 12692 14405 12748
rect 14341 12688 14405 12692
rect 14421 12748 14485 12752
rect 14421 12692 14425 12748
rect 14425 12692 14481 12748
rect 14481 12692 14485 12748
rect 14421 12688 14485 12692
rect 14501 12748 14565 12752
rect 14501 12692 14505 12748
rect 14505 12692 14561 12748
rect 14561 12692 14565 12748
rect 14501 12688 14565 12692
rect 14581 12748 14645 12752
rect 14581 12692 14585 12748
rect 14585 12692 14641 12748
rect 14641 12692 14645 12748
rect 14581 12688 14645 12692
rect 18159 12748 18223 12752
rect 18159 12692 18163 12748
rect 18163 12692 18219 12748
rect 18219 12692 18223 12748
rect 18159 12688 18223 12692
rect 18239 12748 18303 12752
rect 18239 12692 18243 12748
rect 18243 12692 18299 12748
rect 18299 12692 18303 12748
rect 18239 12688 18303 12692
rect 18319 12748 18383 12752
rect 18319 12692 18323 12748
rect 18323 12692 18379 12748
rect 18379 12692 18383 12748
rect 18319 12688 18383 12692
rect 18399 12748 18463 12752
rect 18399 12692 18403 12748
rect 18403 12692 18459 12748
rect 18459 12692 18463 12748
rect 18399 12688 18463 12692
rect 6045 12204 6109 12208
rect 6045 12148 6049 12204
rect 6049 12148 6105 12204
rect 6105 12148 6109 12204
rect 6045 12144 6109 12148
rect 6125 12204 6189 12208
rect 6125 12148 6129 12204
rect 6129 12148 6185 12204
rect 6185 12148 6189 12204
rect 6125 12144 6189 12148
rect 6205 12204 6269 12208
rect 6205 12148 6209 12204
rect 6209 12148 6265 12204
rect 6265 12148 6269 12204
rect 6205 12144 6269 12148
rect 6285 12204 6349 12208
rect 6285 12148 6289 12204
rect 6289 12148 6345 12204
rect 6345 12148 6349 12204
rect 6285 12144 6349 12148
rect 9863 12204 9927 12208
rect 9863 12148 9867 12204
rect 9867 12148 9923 12204
rect 9923 12148 9927 12204
rect 9863 12144 9927 12148
rect 9943 12204 10007 12208
rect 9943 12148 9947 12204
rect 9947 12148 10003 12204
rect 10003 12148 10007 12204
rect 9943 12144 10007 12148
rect 10023 12204 10087 12208
rect 10023 12148 10027 12204
rect 10027 12148 10083 12204
rect 10083 12148 10087 12204
rect 10023 12144 10087 12148
rect 10103 12204 10167 12208
rect 10103 12148 10107 12204
rect 10107 12148 10163 12204
rect 10163 12148 10167 12204
rect 10103 12144 10167 12148
rect 13681 12204 13745 12208
rect 13681 12148 13685 12204
rect 13685 12148 13741 12204
rect 13741 12148 13745 12204
rect 13681 12144 13745 12148
rect 13761 12204 13825 12208
rect 13761 12148 13765 12204
rect 13765 12148 13821 12204
rect 13821 12148 13825 12204
rect 13761 12144 13825 12148
rect 13841 12204 13905 12208
rect 13841 12148 13845 12204
rect 13845 12148 13901 12204
rect 13901 12148 13905 12204
rect 13841 12144 13905 12148
rect 13921 12204 13985 12208
rect 13921 12148 13925 12204
rect 13925 12148 13981 12204
rect 13981 12148 13985 12204
rect 13921 12144 13985 12148
rect 17499 12204 17563 12208
rect 17499 12148 17503 12204
rect 17503 12148 17559 12204
rect 17559 12148 17563 12204
rect 17499 12144 17563 12148
rect 17579 12204 17643 12208
rect 17579 12148 17583 12204
rect 17583 12148 17639 12204
rect 17639 12148 17643 12204
rect 17579 12144 17643 12148
rect 17659 12204 17723 12208
rect 17659 12148 17663 12204
rect 17663 12148 17719 12204
rect 17719 12148 17723 12204
rect 17659 12144 17723 12148
rect 17739 12204 17803 12208
rect 17739 12148 17743 12204
rect 17743 12148 17799 12204
rect 17799 12148 17803 12204
rect 17739 12144 17803 12148
rect 30920 4090 31040 4210
rect 32950 4100 33030 4200
rect 29740 918 29804 3862
<< mimcap >>
rect 29919 3750 34719 3790
rect 29919 1030 29959 3750
rect 34679 1030 34719 3750
rect 29919 990 34719 1030
<< mimcapcontact >>
rect 29959 1030 34679 3750
<< metal4 >>
rect 6037 27440 6357 27456
rect 6037 27376 6045 27440
rect 6109 27376 6125 27440
rect 6189 27376 6205 27440
rect 6269 27376 6285 27440
rect 6349 27376 6357 27440
rect 6037 26352 6357 27376
rect 6037 26288 6045 26352
rect 6109 26288 6125 26352
rect 6189 26288 6205 26352
rect 6269 26288 6285 26352
rect 6349 26288 6357 26352
rect 6037 26282 6357 26288
rect 6037 26046 6079 26282
rect 6315 26046 6357 26282
rect 6037 25264 6357 26046
rect 6037 25200 6045 25264
rect 6109 25200 6125 25264
rect 6189 25200 6205 25264
rect 6269 25200 6285 25264
rect 6349 25200 6357 25264
rect 6037 24176 6357 25200
rect 6037 24112 6045 24176
rect 6109 24112 6125 24176
rect 6189 24112 6205 24176
rect 6269 24112 6285 24176
rect 6349 24112 6357 24176
rect 6037 23088 6357 24112
rect 6037 23024 6045 23088
rect 6109 23024 6125 23088
rect 6189 23024 6205 23088
rect 6269 23024 6285 23088
rect 6349 23024 6357 23088
rect 6037 22474 6357 23024
rect 6037 22238 6079 22474
rect 6315 22238 6357 22474
rect 6037 22000 6357 22238
rect 6037 21936 6045 22000
rect 6109 21936 6125 22000
rect 6189 21936 6205 22000
rect 6269 21936 6285 22000
rect 6349 21936 6357 22000
rect 6037 20912 6357 21936
rect 6037 20848 6045 20912
rect 6109 20848 6125 20912
rect 6189 20848 6205 20912
rect 6269 20848 6285 20912
rect 6349 20848 6357 20912
rect 6037 19824 6357 20848
rect 6037 19760 6045 19824
rect 6109 19760 6125 19824
rect 6189 19760 6205 19824
rect 6269 19760 6285 19824
rect 6349 19760 6357 19824
rect 6037 18736 6357 19760
rect 6037 18672 6045 18736
rect 6109 18672 6125 18736
rect 6189 18672 6205 18736
rect 6269 18672 6285 18736
rect 6349 18672 6357 18736
rect 6037 18666 6357 18672
rect 6037 18430 6079 18666
rect 6315 18430 6357 18666
rect 6037 17648 6357 18430
rect 6037 17584 6045 17648
rect 6109 17584 6125 17648
rect 6189 17584 6205 17648
rect 6269 17584 6285 17648
rect 6349 17584 6357 17648
rect 6037 16560 6357 17584
rect 6037 16496 6045 16560
rect 6109 16496 6125 16560
rect 6189 16496 6205 16560
rect 6269 16496 6285 16560
rect 6349 16496 6357 16560
rect 6037 15472 6357 16496
rect 6037 15408 6045 15472
rect 6109 15408 6125 15472
rect 6189 15408 6205 15472
rect 6269 15408 6285 15472
rect 6349 15408 6357 15472
rect 6037 14858 6357 15408
rect 6037 14622 6079 14858
rect 6315 14622 6357 14858
rect 6037 14384 6357 14622
rect 6037 14320 6045 14384
rect 6109 14320 6125 14384
rect 6189 14320 6205 14384
rect 6269 14320 6285 14384
rect 6349 14320 6357 14384
rect 6037 13296 6357 14320
rect 6037 13232 6045 13296
rect 6109 13232 6125 13296
rect 6189 13232 6205 13296
rect 6269 13232 6285 13296
rect 6349 13232 6357 13296
rect 6037 12208 6357 13232
rect 6037 12144 6045 12208
rect 6109 12144 6125 12208
rect 6189 12144 6205 12208
rect 6269 12144 6285 12208
rect 6349 12144 6357 12208
rect 6037 12128 6357 12144
rect 6697 26896 7017 27456
rect 6697 26832 6705 26896
rect 6769 26832 6785 26896
rect 6849 26832 6865 26896
rect 6929 26832 6945 26896
rect 7009 26832 7017 26896
rect 6697 25808 7017 26832
rect 6697 25744 6705 25808
rect 6769 25744 6785 25808
rect 6849 25744 6865 25808
rect 6929 25744 6945 25808
rect 7009 25744 7017 25808
rect 6697 25622 7017 25744
rect 6697 25386 6739 25622
rect 6975 25386 7017 25622
rect 6697 24720 7017 25386
rect 6697 24656 6705 24720
rect 6769 24656 6785 24720
rect 6849 24656 6865 24720
rect 6929 24656 6945 24720
rect 7009 24656 7017 24720
rect 6697 23632 7017 24656
rect 6697 23568 6705 23632
rect 6769 23568 6785 23632
rect 6849 23568 6865 23632
rect 6929 23568 6945 23632
rect 7009 23568 7017 23632
rect 6697 22544 7017 23568
rect 6697 22480 6705 22544
rect 6769 22480 6785 22544
rect 6849 22480 6865 22544
rect 6929 22480 6945 22544
rect 7009 22480 7017 22544
rect 6697 21814 7017 22480
rect 6697 21578 6739 21814
rect 6975 21578 7017 21814
rect 6697 21456 7017 21578
rect 6697 21392 6705 21456
rect 6769 21392 6785 21456
rect 6849 21392 6865 21456
rect 6929 21392 6945 21456
rect 7009 21392 7017 21456
rect 6697 20368 7017 21392
rect 6697 20304 6705 20368
rect 6769 20304 6785 20368
rect 6849 20304 6865 20368
rect 6929 20304 6945 20368
rect 7009 20304 7017 20368
rect 6697 19280 7017 20304
rect 6697 19216 6705 19280
rect 6769 19216 6785 19280
rect 6849 19216 6865 19280
rect 6929 19216 6945 19280
rect 7009 19216 7017 19280
rect 6697 18192 7017 19216
rect 6697 18128 6705 18192
rect 6769 18128 6785 18192
rect 6849 18128 6865 18192
rect 6929 18128 6945 18192
rect 7009 18128 7017 18192
rect 6697 18006 7017 18128
rect 6697 17770 6739 18006
rect 6975 17770 7017 18006
rect 6697 17104 7017 17770
rect 6697 17040 6705 17104
rect 6769 17040 6785 17104
rect 6849 17040 6865 17104
rect 6929 17040 6945 17104
rect 7009 17040 7017 17104
rect 6697 16016 7017 17040
rect 6697 15952 6705 16016
rect 6769 15952 6785 16016
rect 6849 15952 6865 16016
rect 6929 15952 6945 16016
rect 7009 15952 7017 16016
rect 6697 14928 7017 15952
rect 6697 14864 6705 14928
rect 6769 14864 6785 14928
rect 6849 14864 6865 14928
rect 6929 14864 6945 14928
rect 7009 14864 7017 14928
rect 6697 14198 7017 14864
rect 6697 13962 6739 14198
rect 6975 13962 7017 14198
rect 6697 13840 7017 13962
rect 6697 13776 6705 13840
rect 6769 13776 6785 13840
rect 6849 13776 6865 13840
rect 6929 13776 6945 13840
rect 7009 13776 7017 13840
rect 6697 12752 7017 13776
rect 6697 12688 6705 12752
rect 6769 12688 6785 12752
rect 6849 12688 6865 12752
rect 6929 12688 6945 12752
rect 7009 12688 7017 12752
rect 6697 12128 7017 12688
rect 9855 27440 10175 27456
rect 9855 27376 9863 27440
rect 9927 27376 9943 27440
rect 10007 27376 10023 27440
rect 10087 27376 10103 27440
rect 10167 27376 10175 27440
rect 9855 26352 10175 27376
rect 9855 26288 9863 26352
rect 9927 26288 9943 26352
rect 10007 26288 10023 26352
rect 10087 26288 10103 26352
rect 10167 26288 10175 26352
rect 9855 26282 10175 26288
rect 9855 26046 9897 26282
rect 10133 26046 10175 26282
rect 9855 25264 10175 26046
rect 9855 25200 9863 25264
rect 9927 25200 9943 25264
rect 10007 25200 10023 25264
rect 10087 25200 10103 25264
rect 10167 25200 10175 25264
rect 9855 24176 10175 25200
rect 9855 24112 9863 24176
rect 9927 24112 9943 24176
rect 10007 24112 10023 24176
rect 10087 24112 10103 24176
rect 10167 24112 10175 24176
rect 9855 23088 10175 24112
rect 9855 23024 9863 23088
rect 9927 23024 9943 23088
rect 10007 23024 10023 23088
rect 10087 23024 10103 23088
rect 10167 23024 10175 23088
rect 9855 22474 10175 23024
rect 9855 22238 9897 22474
rect 10133 22238 10175 22474
rect 9855 22000 10175 22238
rect 9855 21936 9863 22000
rect 9927 21936 9943 22000
rect 10007 21936 10023 22000
rect 10087 21936 10103 22000
rect 10167 21936 10175 22000
rect 9855 20912 10175 21936
rect 9855 20848 9863 20912
rect 9927 20848 9943 20912
rect 10007 20848 10023 20912
rect 10087 20848 10103 20912
rect 10167 20848 10175 20912
rect 9855 19824 10175 20848
rect 9855 19760 9863 19824
rect 9927 19760 9943 19824
rect 10007 19760 10023 19824
rect 10087 19760 10103 19824
rect 10167 19760 10175 19824
rect 9855 18736 10175 19760
rect 9855 18672 9863 18736
rect 9927 18672 9943 18736
rect 10007 18672 10023 18736
rect 10087 18672 10103 18736
rect 10167 18672 10175 18736
rect 9855 18666 10175 18672
rect 9855 18430 9897 18666
rect 10133 18430 10175 18666
rect 9855 17648 10175 18430
rect 9855 17584 9863 17648
rect 9927 17584 9943 17648
rect 10007 17584 10023 17648
rect 10087 17584 10103 17648
rect 10167 17584 10175 17648
rect 9855 16560 10175 17584
rect 9855 16496 9863 16560
rect 9927 16496 9943 16560
rect 10007 16496 10023 16560
rect 10087 16496 10103 16560
rect 10167 16496 10175 16560
rect 9855 15472 10175 16496
rect 9855 15408 9863 15472
rect 9927 15408 9943 15472
rect 10007 15408 10023 15472
rect 10087 15408 10103 15472
rect 10167 15408 10175 15472
rect 9855 14858 10175 15408
rect 9855 14622 9897 14858
rect 10133 14622 10175 14858
rect 9855 14384 10175 14622
rect 9855 14320 9863 14384
rect 9927 14320 9943 14384
rect 10007 14320 10023 14384
rect 10087 14320 10103 14384
rect 10167 14320 10175 14384
rect 9855 13296 10175 14320
rect 9855 13232 9863 13296
rect 9927 13232 9943 13296
rect 10007 13232 10023 13296
rect 10087 13232 10103 13296
rect 10167 13232 10175 13296
rect 9855 12208 10175 13232
rect 9855 12144 9863 12208
rect 9927 12144 9943 12208
rect 10007 12144 10023 12208
rect 10087 12144 10103 12208
rect 10167 12144 10175 12208
rect 9855 12128 10175 12144
rect 10515 26896 10835 27456
rect 10515 26832 10523 26896
rect 10587 26832 10603 26896
rect 10667 26832 10683 26896
rect 10747 26832 10763 26896
rect 10827 26832 10835 26896
rect 10515 25808 10835 26832
rect 10515 25744 10523 25808
rect 10587 25744 10603 25808
rect 10667 25744 10683 25808
rect 10747 25744 10763 25808
rect 10827 25744 10835 25808
rect 10515 25622 10835 25744
rect 10515 25386 10557 25622
rect 10793 25386 10835 25622
rect 10515 24720 10835 25386
rect 10515 24656 10523 24720
rect 10587 24656 10603 24720
rect 10667 24656 10683 24720
rect 10747 24656 10763 24720
rect 10827 24656 10835 24720
rect 10515 23632 10835 24656
rect 10515 23568 10523 23632
rect 10587 23568 10603 23632
rect 10667 23568 10683 23632
rect 10747 23568 10763 23632
rect 10827 23568 10835 23632
rect 10515 22544 10835 23568
rect 10515 22480 10523 22544
rect 10587 22480 10603 22544
rect 10667 22480 10683 22544
rect 10747 22480 10763 22544
rect 10827 22480 10835 22544
rect 10515 21814 10835 22480
rect 10515 21578 10557 21814
rect 10793 21578 10835 21814
rect 10515 21456 10835 21578
rect 10515 21392 10523 21456
rect 10587 21392 10603 21456
rect 10667 21392 10683 21456
rect 10747 21392 10763 21456
rect 10827 21392 10835 21456
rect 10515 20368 10835 21392
rect 10515 20304 10523 20368
rect 10587 20304 10603 20368
rect 10667 20304 10683 20368
rect 10747 20304 10763 20368
rect 10827 20304 10835 20368
rect 10515 19280 10835 20304
rect 10515 19216 10523 19280
rect 10587 19216 10603 19280
rect 10667 19216 10683 19280
rect 10747 19216 10763 19280
rect 10827 19216 10835 19280
rect 10515 18192 10835 19216
rect 10515 18128 10523 18192
rect 10587 18128 10603 18192
rect 10667 18128 10683 18192
rect 10747 18128 10763 18192
rect 10827 18128 10835 18192
rect 10515 18006 10835 18128
rect 10515 17770 10557 18006
rect 10793 17770 10835 18006
rect 10515 17104 10835 17770
rect 10515 17040 10523 17104
rect 10587 17040 10603 17104
rect 10667 17040 10683 17104
rect 10747 17040 10763 17104
rect 10827 17040 10835 17104
rect 10515 16016 10835 17040
rect 10515 15952 10523 16016
rect 10587 15952 10603 16016
rect 10667 15952 10683 16016
rect 10747 15952 10763 16016
rect 10827 15952 10835 16016
rect 10515 14928 10835 15952
rect 10515 14864 10523 14928
rect 10587 14864 10603 14928
rect 10667 14864 10683 14928
rect 10747 14864 10763 14928
rect 10827 14864 10835 14928
rect 10515 14198 10835 14864
rect 10515 13962 10557 14198
rect 10793 13962 10835 14198
rect 10515 13840 10835 13962
rect 10515 13776 10523 13840
rect 10587 13776 10603 13840
rect 10667 13776 10683 13840
rect 10747 13776 10763 13840
rect 10827 13776 10835 13840
rect 10515 12752 10835 13776
rect 10515 12688 10523 12752
rect 10587 12688 10603 12752
rect 10667 12688 10683 12752
rect 10747 12688 10763 12752
rect 10827 12688 10835 12752
rect 10515 12128 10835 12688
rect 13673 27440 13993 27456
rect 13673 27376 13681 27440
rect 13745 27376 13761 27440
rect 13825 27376 13841 27440
rect 13905 27376 13921 27440
rect 13985 27376 13993 27440
rect 13673 26352 13993 27376
rect 13673 26288 13681 26352
rect 13745 26288 13761 26352
rect 13825 26288 13841 26352
rect 13905 26288 13921 26352
rect 13985 26288 13993 26352
rect 13673 26282 13993 26288
rect 13673 26046 13715 26282
rect 13951 26046 13993 26282
rect 13673 25264 13993 26046
rect 13673 25200 13681 25264
rect 13745 25200 13761 25264
rect 13825 25200 13841 25264
rect 13905 25200 13921 25264
rect 13985 25200 13993 25264
rect 13673 24176 13993 25200
rect 13673 24112 13681 24176
rect 13745 24112 13761 24176
rect 13825 24112 13841 24176
rect 13905 24112 13921 24176
rect 13985 24112 13993 24176
rect 13673 23088 13993 24112
rect 13673 23024 13681 23088
rect 13745 23024 13761 23088
rect 13825 23024 13841 23088
rect 13905 23024 13921 23088
rect 13985 23024 13993 23088
rect 13673 22474 13993 23024
rect 13673 22238 13715 22474
rect 13951 22238 13993 22474
rect 13673 22000 13993 22238
rect 13673 21936 13681 22000
rect 13745 21936 13761 22000
rect 13825 21936 13841 22000
rect 13905 21936 13921 22000
rect 13985 21936 13993 22000
rect 13673 20912 13993 21936
rect 13673 20848 13681 20912
rect 13745 20848 13761 20912
rect 13825 20848 13841 20912
rect 13905 20848 13921 20912
rect 13985 20848 13993 20912
rect 13673 19824 13993 20848
rect 13673 19760 13681 19824
rect 13745 19760 13761 19824
rect 13825 19760 13841 19824
rect 13905 19760 13921 19824
rect 13985 19760 13993 19824
rect 13673 18736 13993 19760
rect 13673 18672 13681 18736
rect 13745 18672 13761 18736
rect 13825 18672 13841 18736
rect 13905 18672 13921 18736
rect 13985 18672 13993 18736
rect 13673 18666 13993 18672
rect 13673 18430 13715 18666
rect 13951 18430 13993 18666
rect 13673 17648 13993 18430
rect 13673 17584 13681 17648
rect 13745 17584 13761 17648
rect 13825 17584 13841 17648
rect 13905 17584 13921 17648
rect 13985 17584 13993 17648
rect 13673 16560 13993 17584
rect 13673 16496 13681 16560
rect 13745 16496 13761 16560
rect 13825 16496 13841 16560
rect 13905 16496 13921 16560
rect 13985 16496 13993 16560
rect 13673 15472 13993 16496
rect 13673 15408 13681 15472
rect 13745 15408 13761 15472
rect 13825 15408 13841 15472
rect 13905 15408 13921 15472
rect 13985 15408 13993 15472
rect 13673 14858 13993 15408
rect 13673 14622 13715 14858
rect 13951 14622 13993 14858
rect 13673 14384 13993 14622
rect 13673 14320 13681 14384
rect 13745 14320 13761 14384
rect 13825 14320 13841 14384
rect 13905 14320 13921 14384
rect 13985 14320 13993 14384
rect 13673 13296 13993 14320
rect 13673 13232 13681 13296
rect 13745 13232 13761 13296
rect 13825 13232 13841 13296
rect 13905 13232 13921 13296
rect 13985 13232 13993 13296
rect 13673 12208 13993 13232
rect 13673 12144 13681 12208
rect 13745 12144 13761 12208
rect 13825 12144 13841 12208
rect 13905 12144 13921 12208
rect 13985 12144 13993 12208
rect 13673 12128 13993 12144
rect 14333 26896 14653 27456
rect 14333 26832 14341 26896
rect 14405 26832 14421 26896
rect 14485 26832 14501 26896
rect 14565 26832 14581 26896
rect 14645 26832 14653 26896
rect 14333 25808 14653 26832
rect 14333 25744 14341 25808
rect 14405 25744 14421 25808
rect 14485 25744 14501 25808
rect 14565 25744 14581 25808
rect 14645 25744 14653 25808
rect 14333 25622 14653 25744
rect 14333 25386 14375 25622
rect 14611 25386 14653 25622
rect 14333 24720 14653 25386
rect 14333 24656 14341 24720
rect 14405 24656 14421 24720
rect 14485 24656 14501 24720
rect 14565 24656 14581 24720
rect 14645 24656 14653 24720
rect 14333 23632 14653 24656
rect 14333 23568 14341 23632
rect 14405 23568 14421 23632
rect 14485 23568 14501 23632
rect 14565 23568 14581 23632
rect 14645 23568 14653 23632
rect 14333 22544 14653 23568
rect 14333 22480 14341 22544
rect 14405 22480 14421 22544
rect 14485 22480 14501 22544
rect 14565 22480 14581 22544
rect 14645 22480 14653 22544
rect 14333 21814 14653 22480
rect 14333 21578 14375 21814
rect 14611 21578 14653 21814
rect 14333 21456 14653 21578
rect 14333 21392 14341 21456
rect 14405 21392 14421 21456
rect 14485 21392 14501 21456
rect 14565 21392 14581 21456
rect 14645 21392 14653 21456
rect 14333 20368 14653 21392
rect 14333 20304 14341 20368
rect 14405 20304 14421 20368
rect 14485 20304 14501 20368
rect 14565 20304 14581 20368
rect 14645 20304 14653 20368
rect 14333 19280 14653 20304
rect 14333 19216 14341 19280
rect 14405 19216 14421 19280
rect 14485 19216 14501 19280
rect 14565 19216 14581 19280
rect 14645 19216 14653 19280
rect 14333 18192 14653 19216
rect 14333 18128 14341 18192
rect 14405 18128 14421 18192
rect 14485 18128 14501 18192
rect 14565 18128 14581 18192
rect 14645 18128 14653 18192
rect 14333 18006 14653 18128
rect 14333 17770 14375 18006
rect 14611 17770 14653 18006
rect 14333 17104 14653 17770
rect 14333 17040 14341 17104
rect 14405 17040 14421 17104
rect 14485 17040 14501 17104
rect 14565 17040 14581 17104
rect 14645 17040 14653 17104
rect 14333 16016 14653 17040
rect 14333 15952 14341 16016
rect 14405 15952 14421 16016
rect 14485 15952 14501 16016
rect 14565 15952 14581 16016
rect 14645 15952 14653 16016
rect 14333 14928 14653 15952
rect 14333 14864 14341 14928
rect 14405 14864 14421 14928
rect 14485 14864 14501 14928
rect 14565 14864 14581 14928
rect 14645 14864 14653 14928
rect 14333 14198 14653 14864
rect 14333 13962 14375 14198
rect 14611 13962 14653 14198
rect 14333 13840 14653 13962
rect 14333 13776 14341 13840
rect 14405 13776 14421 13840
rect 14485 13776 14501 13840
rect 14565 13776 14581 13840
rect 14645 13776 14653 13840
rect 14333 12752 14653 13776
rect 14333 12688 14341 12752
rect 14405 12688 14421 12752
rect 14485 12688 14501 12752
rect 14565 12688 14581 12752
rect 14645 12688 14653 12752
rect 14333 12128 14653 12688
rect 17491 27440 17811 27456
rect 17491 27376 17499 27440
rect 17563 27376 17579 27440
rect 17643 27376 17659 27440
rect 17723 27376 17739 27440
rect 17803 27376 17811 27440
rect 17491 26352 17811 27376
rect 17491 26288 17499 26352
rect 17563 26288 17579 26352
rect 17643 26288 17659 26352
rect 17723 26288 17739 26352
rect 17803 26288 17811 26352
rect 17491 26282 17811 26288
rect 17491 26046 17533 26282
rect 17769 26046 17811 26282
rect 17491 25264 17811 26046
rect 17491 25200 17499 25264
rect 17563 25200 17579 25264
rect 17643 25200 17659 25264
rect 17723 25200 17739 25264
rect 17803 25200 17811 25264
rect 17491 24176 17811 25200
rect 17491 24112 17499 24176
rect 17563 24112 17579 24176
rect 17643 24112 17659 24176
rect 17723 24112 17739 24176
rect 17803 24112 17811 24176
rect 17491 23088 17811 24112
rect 17491 23024 17499 23088
rect 17563 23024 17579 23088
rect 17643 23024 17659 23088
rect 17723 23024 17739 23088
rect 17803 23024 17811 23088
rect 17491 22474 17811 23024
rect 17491 22238 17533 22474
rect 17769 22238 17811 22474
rect 17491 22000 17811 22238
rect 17491 21936 17499 22000
rect 17563 21936 17579 22000
rect 17643 21936 17659 22000
rect 17723 21936 17739 22000
rect 17803 21936 17811 22000
rect 17491 20912 17811 21936
rect 17491 20848 17499 20912
rect 17563 20848 17579 20912
rect 17643 20848 17659 20912
rect 17723 20848 17739 20912
rect 17803 20848 17811 20912
rect 17491 19824 17811 20848
rect 17491 19760 17499 19824
rect 17563 19760 17579 19824
rect 17643 19760 17659 19824
rect 17723 19760 17739 19824
rect 17803 19760 17811 19824
rect 17491 18736 17811 19760
rect 17491 18672 17499 18736
rect 17563 18672 17579 18736
rect 17643 18672 17659 18736
rect 17723 18672 17739 18736
rect 17803 18672 17811 18736
rect 17491 18666 17811 18672
rect 17491 18430 17533 18666
rect 17769 18430 17811 18666
rect 17491 17648 17811 18430
rect 17491 17584 17499 17648
rect 17563 17584 17579 17648
rect 17643 17584 17659 17648
rect 17723 17584 17739 17648
rect 17803 17584 17811 17648
rect 17491 16560 17811 17584
rect 17491 16496 17499 16560
rect 17563 16496 17579 16560
rect 17643 16496 17659 16560
rect 17723 16496 17739 16560
rect 17803 16496 17811 16560
rect 17491 15472 17811 16496
rect 17491 15408 17499 15472
rect 17563 15408 17579 15472
rect 17643 15408 17659 15472
rect 17723 15408 17739 15472
rect 17803 15408 17811 15472
rect 17491 14858 17811 15408
rect 17491 14622 17533 14858
rect 17769 14622 17811 14858
rect 17491 14384 17811 14622
rect 17491 14320 17499 14384
rect 17563 14320 17579 14384
rect 17643 14320 17659 14384
rect 17723 14320 17739 14384
rect 17803 14320 17811 14384
rect 17491 13296 17811 14320
rect 17491 13232 17499 13296
rect 17563 13232 17579 13296
rect 17643 13232 17659 13296
rect 17723 13232 17739 13296
rect 17803 13232 17811 13296
rect 17491 12208 17811 13232
rect 17491 12144 17499 12208
rect 17563 12144 17579 12208
rect 17643 12144 17659 12208
rect 17723 12144 17739 12208
rect 17803 12144 17811 12208
rect 17491 12128 17811 12144
rect 18151 26896 18471 27456
rect 18151 26832 18159 26896
rect 18223 26832 18239 26896
rect 18303 26832 18319 26896
rect 18383 26832 18399 26896
rect 18463 26832 18471 26896
rect 18151 25808 18471 26832
rect 18151 25744 18159 25808
rect 18223 25744 18239 25808
rect 18303 25744 18319 25808
rect 18383 25744 18399 25808
rect 18463 25744 18471 25808
rect 18151 25622 18471 25744
rect 18151 25386 18193 25622
rect 18429 25386 18471 25622
rect 18151 24720 18471 25386
rect 18151 24656 18159 24720
rect 18223 24656 18239 24720
rect 18303 24656 18319 24720
rect 18383 24656 18399 24720
rect 18463 24656 18471 24720
rect 18151 23632 18471 24656
rect 18151 23568 18159 23632
rect 18223 23568 18239 23632
rect 18303 23568 18319 23632
rect 18383 23568 18399 23632
rect 18463 23568 18471 23632
rect 18151 22544 18471 23568
rect 18151 22480 18159 22544
rect 18223 22480 18239 22544
rect 18303 22480 18319 22544
rect 18383 22480 18399 22544
rect 18463 22480 18471 22544
rect 18151 21814 18471 22480
rect 18151 21578 18193 21814
rect 18429 21578 18471 21814
rect 18151 21456 18471 21578
rect 18151 21392 18159 21456
rect 18223 21392 18239 21456
rect 18303 21392 18319 21456
rect 18383 21392 18399 21456
rect 18463 21392 18471 21456
rect 18151 20368 18471 21392
rect 18151 20304 18159 20368
rect 18223 20304 18239 20368
rect 18303 20304 18319 20368
rect 18383 20304 18399 20368
rect 18463 20304 18471 20368
rect 18151 19280 18471 20304
rect 18151 19216 18159 19280
rect 18223 19216 18239 19280
rect 18303 19216 18319 19280
rect 18383 19216 18399 19280
rect 18463 19216 18471 19280
rect 18151 18192 18471 19216
rect 18151 18128 18159 18192
rect 18223 18128 18239 18192
rect 18303 18128 18319 18192
rect 18383 18128 18399 18192
rect 18463 18128 18471 18192
rect 18151 18006 18471 18128
rect 18151 17770 18193 18006
rect 18429 17770 18471 18006
rect 18151 17104 18471 17770
rect 18151 17040 18159 17104
rect 18223 17040 18239 17104
rect 18303 17040 18319 17104
rect 18383 17040 18399 17104
rect 18463 17040 18471 17104
rect 18151 16016 18471 17040
rect 18151 15952 18159 16016
rect 18223 15952 18239 16016
rect 18303 15952 18319 16016
rect 18383 15952 18399 16016
rect 18463 15952 18471 16016
rect 18151 14928 18471 15952
rect 18151 14864 18159 14928
rect 18223 14864 18239 14928
rect 18303 14864 18319 14928
rect 18383 14864 18399 14928
rect 18463 14864 18471 14928
rect 18151 14198 18471 14864
rect 18151 13962 18193 14198
rect 18429 13962 18471 14198
rect 18151 13840 18471 13962
rect 18151 13776 18159 13840
rect 18223 13776 18239 13840
rect 18303 13776 18319 13840
rect 18383 13776 18399 13840
rect 18463 13776 18471 13840
rect 18151 12752 18471 13776
rect 18151 12688 18159 12752
rect 18223 12688 18239 12752
rect 18303 12688 18319 12752
rect 18383 12688 18399 12752
rect 18463 12688 18471 12752
rect 18151 12128 18471 12688
rect 30900 4210 31050 4220
rect 30900 4090 30920 4210
rect 31040 4090 31050 4210
rect 30900 4040 31050 4090
rect 29665 3950 31050 4040
rect 32940 4200 33040 4210
rect 32940 4100 32950 4200
rect 33030 4100 33040 4200
rect 29665 3878 29800 3950
rect 29665 3862 29820 3878
rect 29665 3675 29740 3862
rect 29724 918 29740 3675
rect 29804 918 29820 3862
rect 32940 3751 33040 4100
rect 29958 3750 34680 3751
rect 29958 1030 29959 3750
rect 34679 1030 34680 3750
rect 29958 1029 34680 1030
rect 29724 902 29820 918
<< via4 >>
rect 6079 26046 6315 26282
rect 6079 22238 6315 22474
rect 6079 18430 6315 18666
rect 6079 14622 6315 14858
rect 6739 25386 6975 25622
rect 6739 21578 6975 21814
rect 6739 17770 6975 18006
rect 6739 13962 6975 14198
rect 9897 26046 10133 26282
rect 9897 22238 10133 22474
rect 9897 18430 10133 18666
rect 9897 14622 10133 14858
rect 10557 25386 10793 25622
rect 10557 21578 10793 21814
rect 10557 17770 10793 18006
rect 10557 13962 10793 14198
rect 13715 26046 13951 26282
rect 13715 22238 13951 22474
rect 13715 18430 13951 18666
rect 13715 14622 13951 14858
rect 14375 25386 14611 25622
rect 14375 21578 14611 21814
rect 14375 17770 14611 18006
rect 14375 13962 14611 14198
rect 17533 26046 17769 26282
rect 17533 22238 17769 22474
rect 17533 18430 17769 18666
rect 17533 14622 17769 14858
rect 18193 25386 18429 25622
rect 18193 21578 18429 21814
rect 18193 17770 18429 18006
rect 18193 13962 18429 14198
<< metal5 >>
rect 4900 26282 20268 26324
rect 4900 26046 6079 26282
rect 6315 26046 9897 26282
rect 10133 26046 13715 26282
rect 13951 26046 17533 26282
rect 17769 26046 20268 26282
rect 4900 26004 20268 26046
rect 4900 25622 20268 25664
rect 4900 25386 6739 25622
rect 6975 25386 10557 25622
rect 10793 25386 14375 25622
rect 14611 25386 18193 25622
rect 18429 25386 20268 25622
rect 4900 25344 20268 25386
rect 4900 22474 20268 22516
rect 4900 22238 6079 22474
rect 6315 22238 9897 22474
rect 10133 22238 13715 22474
rect 13951 22238 17533 22474
rect 17769 22238 20268 22474
rect 4900 22196 20268 22238
rect 4900 21814 20268 21856
rect 4900 21578 6739 21814
rect 6975 21578 10557 21814
rect 10793 21578 14375 21814
rect 14611 21578 18193 21814
rect 18429 21578 20268 21814
rect 4900 21536 20268 21578
rect 4900 18666 20268 18708
rect 4900 18430 6079 18666
rect 6315 18430 9897 18666
rect 10133 18430 13715 18666
rect 13951 18430 17533 18666
rect 17769 18430 20268 18666
rect 4900 18388 20268 18430
rect 4900 18006 20268 18048
rect 4900 17770 6739 18006
rect 6975 17770 10557 18006
rect 10793 17770 14375 18006
rect 14611 17770 18193 18006
rect 18429 17770 20268 18006
rect 4900 17728 20268 17770
rect 4900 14858 20268 14900
rect 4900 14622 6079 14858
rect 6315 14622 9897 14858
rect 10133 14622 13715 14858
rect 13951 14622 17533 14858
rect 17769 14622 20268 14858
rect 4900 14580 20268 14622
rect 4900 14198 20268 14240
rect 4900 13962 6739 14198
rect 6975 13962 10557 14198
rect 10793 13962 14375 14198
rect 14611 13962 18193 14198
rect 18429 13962 20268 14198
rect 4900 13920 20268 13962
<< res0p35 >>
rect 25844 7576 25918 8664
rect 26162 7576 26236 8664
rect 26480 7576 26554 8664
rect 26798 7576 26872 8664
rect 27116 7576 27190 8664
rect 27434 7576 27508 8664
rect 27752 7576 27826 8664
rect 28070 7576 28144 8664
rect 3514 5236 3588 5440
rect 6814 5236 6888 5344
rect 10114 5236 10188 5484
rect 13414 5236 13488 5764
rect 17014 5236 17088 6324
rect 20214 5236 20288 6324
rect 20532 5236 20606 6324
rect 23314 5236 23388 6324
rect 23632 5236 23706 6324
rect 23950 5236 24024 6324
rect 24268 5236 24342 6324
rect 25814 5236 25888 6324
rect 26132 5236 26206 6324
rect 26450 5236 26524 6324
rect 26768 5236 26842 6324
rect 27086 5236 27160 6324
rect 27404 5236 27478 6324
rect 27722 5236 27796 6324
rect 28040 5236 28114 6324
<< labels >>
flabel space 28700 0 28900 190 0 FreeSans 1600 0 0 0 inp
port 3 nsew
flabel metal2 6000 29510 6200 29700 0 FreeSans 1600 0 0 0 reset
port 6 nsew
flabel metal2 10320 29470 10520 29660 0 FreeSans 1600 0 0 0 sdi
port 7 nsew
flabel metal1 -200 3440 0 3640 0 FreeSans 1600 0 0 0 vd
port 14 nsew
flabel metal1 -200 2500 0 2700 0 FreeSans 1600 0 0 0 gnd
port 5 nsew
flabel metal1 14050 -160 14250 40 0 FreeSans 1600 0 0 0 inn
port 15 nsew
flabel metal1 28700 -200 28900 0 0 FreeSans 1600 0 0 0 inp
port 16 nsew
flabel metal1 35430 5790 35630 5990 0 FreeSans 1600 0 0 0 out
port 17 nsew
flabel metal1 29200 9440 29400 9640 0 FreeSans 1600 0 0 0 ib
port 18 nsew
flabel metal1 -200 19690 0 19880 0 FreeSans 1600 0 0 0 gndd
port 9 nsew
flabel metal2 14650 29470 14850 29660 0 FreeSans 1600 0 0 0 sclk
port 19 nsew
flabel metal2 18980 29470 19180 29660 0 FreeSans 1600 0 0 0 ss
port 21 nsew
flabel metal1 -200 19170 0 19360 0 FreeSans 1600 0 0 0 vpwr
port 11 nsew
flabel metal1 1418 19770 1508 19788 0 FreeSans 1600 0 0 0 vgnd
flabel metal4 17491 12128 17811 27456 0 FreeSans 1920 90 0 0 sr_0.VGND
flabel metal4 13673 12128 13993 27456 0 FreeSans 1920 90 0 0 sr_0.VGND
flabel metal4 9855 12128 10175 27456 0 FreeSans 1920 90 0 0 sr_0.VGND
flabel metal4 6037 12128 6357 27456 0 FreeSans 1920 90 0 0 sr_0.VGND
flabel metal5 4900 14580 20268 14900 0 FreeSans 2560 0 0 0 sr_0.VGND
flabel metal5 4900 18388 20268 18708 0 FreeSans 2560 0 0 0 sr_0.VGND
flabel metal5 4900 22196 20268 22516 0 FreeSans 2560 0 0 0 sr_0.VGND
flabel metal5 4900 26004 20268 26324 0 FreeSans 2560 0 0 0 sr_0.VGND
flabel metal4 18151 12128 18471 27456 0 FreeSans 1920 90 0 0 sr_0.VPWR
flabel metal4 14333 12128 14653 27456 0 FreeSans 1920 90 0 0 sr_0.VPWR
flabel metal4 10515 12128 10835 27456 0 FreeSans 1920 90 0 0 sr_0.VPWR
flabel metal4 6697 12128 7017 27456 0 FreeSans 1920 90 0 0 sr_0.VPWR
flabel metal5 4900 13920 20268 14240 0 FreeSans 2560 0 0 0 sr_0.VPWR
flabel metal5 4900 17728 20268 18048 0 FreeSans 2560 0 0 0 sr_0.VPWR
flabel metal5 4900 21536 20268 21856 0 FreeSans 2560 0 0 0 sr_0.VPWR
flabel metal5 4900 25344 20268 25664 0 FreeSans 2560 0 0 0 sr_0.VPWR
flabel metal2 19962 10000 20018 10800 0 FreeSans 224 90 0 0 sr_0.data[0]
flabel metal2 17846 10000 17902 10800 0 FreeSans 224 90 0 0 sr_0.data[1]
flabel metal2 15730 10000 15786 10800 0 FreeSans 224 90 0 0 sr_0.data[2]
flabel metal2 13614 10000 13670 10800 0 FreeSans 224 90 0 0 sr_0.data[3]
flabel metal2 11498 10000 11554 10800 0 FreeSans 224 90 0 0 sr_0.data[4]
flabel metal2 9382 10000 9438 10800 0 FreeSans 224 90 0 0 sr_0.data[5]
flabel metal2 7266 10000 7322 10800 0 FreeSans 224 90 0 0 sr_0.data[6]
flabel metal2 5150 10000 5206 10800 0 FreeSans 224 90 0 0 sr_0.data[7]
flabel metal2 6070 28856 6126 29656 0 FreeSans 224 90 0 0 sr_0.reset
flabel metal2 14718 28856 14774 29656 0 FreeSans 224 90 0 0 sr_0.sclk
flabel metal2 10394 28856 10450 29656 0 FreeSans 224 90 0 0 sr_0.sdi
flabel metal2 19042 28856 19098 29656 0 FreeSans 224 90 0 0 sr_0.ss
rlabel metal1 12584 27408 12584 27408 0 sr_0.VGND
rlabel metal1 12584 26864 12584 26864 0 sr_0.VPWR
rlabel metal1 15804 12958 15804 12958 0 sr_0._00_
rlabel metal1 14056 12618 14056 12618 0 sr_0._01_
rlabel metal2 12538 13162 12538 13162 0 sr_0._02_
rlabel metal1 11250 12958 11250 12958 0 sr_0._03_
rlabel metal1 11710 14046 11710 14046 0 sr_0._04_
rlabel metal1 15574 12482 15574 12482 0 sr_0._05_
rlabel metal2 16034 14386 16034 14386 0 sr_0._06_
rlabel metal1 16540 13706 16540 13706 0 sr_0._07_
rlabel metal1 15298 14250 15298 14250 0 sr_0._08_
rlabel metal1 14194 12890 14194 12890 0 sr_0._09_
rlabel metal1 13642 12414 13642 12414 0 sr_0._10_
rlabel metal1 12446 12618 12446 12618 0 sr_0._11_
rlabel metal1 10100 12550 10100 12550 0 sr_0._12_
rlabel metal1 12032 14114 12032 14114 0 sr_0._13_
rlabel metal2 14746 13706 14746 13706 0 sr_0.clknet_0_sclk
rlabel metal1 16264 13706 16264 13706 0 sr_0.clknet_1_0__leaf_sclk
rlabel metal2 11894 13876 11894 13876 0 sr_0.clknet_1_1__leaf_sclk
rlabel metal2 19990 11554 19990 11554 0 sr_0.data[0]
rlabel metal2 17874 11554 17874 11554 0 sr_0.data[1]
rlabel metal2 15758 10959 15758 10959 0 sr_0.data[2]
rlabel metal2 13642 10959 13642 10959 0 sr_0.data[3]
rlabel metal2 11526 11792 11526 11792 0 sr_0.data[4]
rlabel metal2 9410 11520 9410 11520 0 sr_0.data[5]
rlabel metal2 7294 11520 7294 11520 0 sr_0.data[6]
rlabel metal1 15535 13026 15535 13026 0 sr_0.net1
rlabel metal1 10330 12414 10330 12414 0 sr_0.net10
rlabel metal2 5178 11027 5178 11027 0 sr_0.net11
rlabel metal1 17000 13162 17000 13162 0 sr_0.net12
rlabel metal1 15252 14114 15252 14114 0 sr_0.net13
rlabel metal1 16172 14114 16172 14114 0 sr_0.net14
rlabel metal1 13090 14692 13090 14692 0 sr_0.net15
rlabel metal1 10376 12482 10376 12482 0 sr_0.net16
rlabel metal2 14746 12856 14746 12856 0 sr_0.net17
rlabel metal1 10698 26966 10698 26966 0 sr_0.net2
rlabel metal1 17966 13570 17966 13570 0 sr_0.net3
rlabel metal2 17598 12686 17598 12686 0 sr_0.net4
rlabel metal2 15666 14352 15666 14352 0 sr_0.net5
rlabel metal2 14194 13434 14194 13434 0 sr_0.net6
rlabel metal1 14470 12992 14470 12992 0 sr_0.net7
rlabel metal1 13458 12822 13458 12822 0 sr_0.net8
rlabel metal1 9824 12958 9824 12958 0 sr_0.net9
rlabel metal2 5914 28105 5914 28105 0 sr_0.reset
rlabel metal2 14746 27146 14746 27146 0 sr_0.sclk
rlabel metal1 10192 27170 10192 27170 0 sr_0.sdi
rlabel metal1 18978 27238 18978 27238 0 sr_0.ss
flabel metal1 19329 12159 19363 12193 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_9.VGND
flabel metal1 19329 12703 19363 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_9.VPWR
flabel nwell 19329 12703 19363 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_9.VPB
flabel pwell 19329 12159 19363 12193 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_9.VNB
rlabel comment 19392 12176 19392 12176 6 sr_0.FILLER_0_0_9.decap_12
flabel metal1 19881 13247 19915 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_3.VGND
flabel metal1 19881 12703 19915 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_3.VPWR
flabel nwell 19881 12703 19915 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_3.VPB
flabel pwell 19881 13247 19915 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_3.VNB
rlabel comment 19944 13264 19944 13264 8 sr_0.FILLER_0_1_3.decap_12
flabel metal1 18777 13247 18811 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_15.VGND
flabel metal1 18777 12703 18811 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_15.VPWR
flabel nwell 18777 12703 18811 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_15.VPB
flabel pwell 18777 13247 18811 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_15.VNB
rlabel comment 18840 13264 18840 13264 8 sr_0.FILLER_0_1_15.decap_12
flabel metal1 20157 12703 20191 12737 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_0_Left_28.VPWR
flabel metal1 20157 12159 20191 12193 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_0_Left_28.VGND
flabel nwell 20157 12703 20191 12737 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_0_Left_28.VPB
flabel pwell 20157 12159 20191 12193 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_0_Left_28.VNB
rlabel comment 20220 12176 20220 12176 6 sr_0.PHY_EDGE_ROW_0_Left_28.decap_3
rlabel metal1 19944 12128 20220 12224 1 sr_0.PHY_EDGE_ROW_0_Left_28.VGND
rlabel metal1 19944 12672 20220 12768 1 sr_0.PHY_EDGE_ROW_0_Left_28.VPWR
flabel metal1 20157 12703 20191 12737 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_1_Left_29.VPWR
flabel metal1 20157 13247 20191 13281 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_1_Left_29.VGND
flabel nwell 20157 12703 20191 12737 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_1_Left_29.VPB
flabel pwell 20157 13247 20191 13281 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_1_Left_29.VNB
rlabel comment 20220 13264 20220 13264 8 sr_0.PHY_EDGE_ROW_1_Left_29.decap_3
rlabel metal1 19944 13216 20220 13312 5 sr_0.PHY_EDGE_ROW_1_Left_29.VGND
rlabel metal1 19944 12672 20220 12768 5 sr_0.PHY_EDGE_ROW_1_Left_29.VPWR
flabel locali 19789 12465 19823 12499 0 FreeSans 200 0 0 0 sr_0.output4.X
flabel locali 19513 12329 19547 12363 0 FreeSans 200 0 0 0 sr_0.output4.A
flabel locali 19881 12329 19915 12363 0 FreeSans 200 0 0 0 sr_0.output4.X
flabel locali 19513 12397 19547 12431 0 FreeSans 200 0 0 0 sr_0.output4.A
flabel locali 19881 12397 19915 12431 0 FreeSans 200 0 0 0 sr_0.output4.X
flabel metal1 19421 12159 19455 12193 0 FreeSans 200 0 0 0 sr_0.output4.VGND
flabel metal1 19421 12703 19455 12737 0 FreeSans 200 0 0 0 sr_0.output4.VPWR
flabel nwell 19421 12703 19455 12737 0 FreeSans 200 0 0 0 sr_0.output4.VPB
flabel pwell 19421 12159 19455 12193 0 FreeSans 200 0 0 0 sr_0.output4.VNB
rlabel comment 19392 12176 19392 12176 4 sr_0.output4.clkbuf_4
rlabel metal1 19392 12128 19944 12224 1 sr_0.output4.VGND
rlabel metal1 19392 12672 19944 12768 1 sr_0.output4.VPWR
flabel metal1 18225 12703 18259 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_21.VPWR
flabel metal1 18225 12159 18259 12193 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_21.VGND
flabel nwell 18225 12703 18259 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_21.VPB
flabel pwell 18225 12159 18259 12193 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_21.VNB
rlabel comment 18288 12176 18288 12176 6 sr_0.FILLER_0_0_21.decap_6
rlabel metal1 17736 12128 18288 12224 1 sr_0.FILLER_0_0_21.VGND
rlabel metal1 17736 12672 18288 12768 1 sr_0.FILLER_0_0_21.VPWR
flabel metal1 17678 12703 17714 12733 0 FreeSans 250 0 0 0 sr_0.FILLER_0_0_27.VPWR
flabel metal1 17678 12163 17714 12192 0 FreeSans 250 0 0 0 sr_0.FILLER_0_0_27.VGND
flabel nwell 17685 12710 17705 12727 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_27.VPB
flabel pwell 17684 12165 17708 12187 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_27.VNB
rlabel comment 17736 12176 17736 12176 6 sr_0.FILLER_0_0_27.fill_1
rlabel metal1 17644 12128 17736 12224 1 sr_0.FILLER_0_0_27.VGND
rlabel metal1 17644 12672 17736 12768 1 sr_0.FILLER_0_0_27.VPWR
flabel metal1 16942 12703 16978 12733 0 FreeSans 250 0 0 0 sr_0.FILLER_0_0_35.VPWR
flabel metal1 16942 12163 16978 12192 0 FreeSans 250 0 0 0 sr_0.FILLER_0_0_35.VGND
flabel nwell 16949 12710 16969 12727 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_35.VPB
flabel pwell 16948 12165 16972 12187 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_35.VNB
rlabel comment 17000 12176 17000 12176 6 sr_0.FILLER_0_0_35.fill_1
rlabel metal1 16908 12128 17000 12224 1 sr_0.FILLER_0_0_35.VGND
rlabel metal1 16908 12672 17000 12768 1 sr_0.FILLER_0_0_35.VPWR
flabel metal1 17678 12707 17714 12737 0 FreeSans 250 0 0 0 sr_0.FILLER_0_1_27.VPWR
flabel metal1 17678 13248 17714 13277 0 FreeSans 250 0 0 0 sr_0.FILLER_0_1_27.VGND
flabel nwell 17685 12713 17705 12730 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_27.VPB
flabel pwell 17684 13253 17708 13275 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_27.VNB
rlabel comment 17736 13264 17736 13264 8 sr_0.FILLER_0_1_27.fill_1
rlabel metal1 17644 13216 17736 13312 5 sr_0.FILLER_0_1_27.VGND
rlabel metal1 17644 12672 17736 12768 5 sr_0.FILLER_0_1_27.VPWR
flabel metal1 17569 12700 17622 12729 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_0_56.VPWR
flabel metal1 17572 12158 17623 12196 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_0_56.VGND
rlabel comment 17644 12176 17644 12176 6 sr_0.TAP_TAPCELL_ROW_0_56.tapvpwrvgnd_1
rlabel metal1 17552 12128 17644 12224 1 sr_0.TAP_TAPCELL_ROW_0_56.VGND
rlabel metal1 17552 12672 17644 12768 1 sr_0.TAP_TAPCELL_ROW_0_56.VPWR
flabel locali 16844 12601 16878 12635 0 FreeSans 400 0 0 0 sr_0._28_.Q
flabel locali 16844 12533 16878 12567 0 FreeSans 400 0 0 0 sr_0._28_.Q
flabel locali 16844 12465 16878 12499 0 FreeSans 400 0 0 0 sr_0._28_.Q
flabel locali 16844 12261 16878 12295 0 FreeSans 400 0 0 0 sr_0._28_.Q
flabel locali 16549 12329 16583 12363 0 FreeSans 400 0 0 0 sr_0._28_.RESET_B
flabel locali 15373 12465 15407 12499 0 FreeSans 400 0 0 0 sr_0._28_.D
flabel locali 15098 12465 15132 12499 0 FreeSans 400 0 0 0 sr_0._28_.CLK
flabel locali 15098 12397 15132 12431 0 FreeSans 400 0 0 0 sr_0._28_.CLK
flabel locali 16549 12397 16583 12431 0 FreeSans 400 0 0 0 sr_0._28_.RESET_B
flabel metal1 15097 12159 15131 12193 0 FreeSans 200 0 0 0 sr_0._28_.VGND
flabel metal1 15097 12703 15131 12737 0 FreeSans 200 0 0 0 sr_0._28_.VPWR
flabel nwell 15097 12703 15131 12737 0 FreeSans 200 0 0 0 sr_0._28_.VPB
flabel pwell 15097 12159 15131 12193 0 FreeSans 200 0 0 0 sr_0._28_.VNB
rlabel comment 15068 12176 15068 12176 4 sr_0._28_.dfrtp_1
rlabel locali 16549 12303 16597 12383 1 sr_0._28_.RESET_B
rlabel locali 16489 12383 16597 12457 1 sr_0._28_.RESET_B
rlabel metal1 16537 12323 16595 12332 1 sr_0._28_.RESET_B
rlabel metal1 16477 12369 16535 12432 1 sr_0._28_.RESET_B
rlabel metal1 16477 12360 16595 12369 1 sr_0._28_.RESET_B
rlabel metal1 15817 12360 15947 12369 1 sr_0._28_.RESET_B
rlabel metal1 15817 12332 16595 12360 1 sr_0._28_.RESET_B
rlabel metal1 15817 12323 15947 12332 1 sr_0._28_.RESET_B
rlabel metal1 15068 12128 16908 12224 1 sr_0._28_.VGND
rlabel metal1 15068 12672 16908 12768 1 sr_0._28_.VPWR
flabel locali 15098 12805 15132 12839 0 FreeSans 400 0 0 0 sr_0._30_.Q
flabel locali 15098 12873 15132 12907 0 FreeSans 400 0 0 0 sr_0._30_.Q
flabel locali 15098 12941 15132 12975 0 FreeSans 400 0 0 0 sr_0._30_.Q
flabel locali 15098 13145 15132 13179 0 FreeSans 400 0 0 0 sr_0._30_.Q
flabel locali 15393 13077 15427 13111 0 FreeSans 400 0 0 0 sr_0._30_.RESET_B
flabel locali 16569 12941 16603 12975 0 FreeSans 400 0 0 0 sr_0._30_.D
flabel locali 16844 12941 16878 12975 0 FreeSans 400 0 0 0 sr_0._30_.CLK
flabel locali 16844 13009 16878 13043 0 FreeSans 400 0 0 0 sr_0._30_.CLK
flabel locali 15393 13009 15427 13043 0 FreeSans 400 0 0 0 sr_0._30_.RESET_B
flabel metal1 16845 13247 16879 13281 0 FreeSans 200 0 0 0 sr_0._30_.VGND
flabel metal1 16845 12703 16879 12737 0 FreeSans 200 0 0 0 sr_0._30_.VPWR
flabel nwell 16845 12703 16879 12737 0 FreeSans 200 0 0 0 sr_0._30_.VPB
flabel pwell 16845 13247 16879 13281 0 FreeSans 200 0 0 0 sr_0._30_.VNB
rlabel comment 16908 13264 16908 13264 8 sr_0._30_.dfrtp_1
rlabel locali 15379 13057 15427 13137 5 sr_0._30_.RESET_B
rlabel locali 15379 12983 15487 13057 5 sr_0._30_.RESET_B
rlabel metal1 15381 13108 15439 13117 5 sr_0._30_.RESET_B
rlabel metal1 15441 13008 15499 13071 5 sr_0._30_.RESET_B
rlabel metal1 15381 13071 15499 13080 5 sr_0._30_.RESET_B
rlabel metal1 16029 13071 16159 13080 5 sr_0._30_.RESET_B
rlabel metal1 15381 13080 16159 13108 5 sr_0._30_.RESET_B
rlabel metal1 16029 13108 16159 13117 5 sr_0._30_.RESET_B
rlabel metal1 15068 13216 16908 13312 5 sr_0._30_.VGND
rlabel metal1 15068 12672 16908 12768 5 sr_0._30_.VPWR
flabel locali 17581 13009 17615 13043 0 FreeSans 200 0 0 0 sr_0.hold1.A
flabel locali 16933 13077 16967 13111 0 FreeSans 200 0 0 0 sr_0.hold1.X
flabel locali 17581 12941 17615 12975 0 FreeSans 200 0 0 0 sr_0.hold1.A
flabel locali 16933 13145 16967 13179 0 FreeSans 200 0 0 0 sr_0.hold1.X
flabel locali 17489 13009 17523 13043 0 FreeSans 200 0 0 0 sr_0.hold1.A
flabel locali 17489 12941 17523 12975 0 FreeSans 200 0 0 0 sr_0.hold1.A
flabel locali 16933 12805 16967 12839 0 FreeSans 200 0 0 0 sr_0.hold1.X
flabel locali 16933 12941 16967 12975 0 FreeSans 200 0 0 0 sr_0.hold1.X
flabel locali 16933 12873 16967 12907 0 FreeSans 200 0 0 0 sr_0.hold1.X
flabel locali 16933 13009 16967 13043 0 FreeSans 200 0 0 0 sr_0.hold1.X
flabel nwell 17581 12703 17615 12737 0 FreeSans 200 0 0 0 sr_0.hold1.VPB
flabel pwell 17581 13247 17615 13281 0 FreeSans 200 0 0 0 sr_0.hold1.VNB
flabel metal1 17581 13247 17615 13281 0 FreeSans 200 0 0 0 sr_0.hold1.VGND
flabel metal1 17581 12703 17615 12737 0 FreeSans 200 0 0 0 sr_0.hold1.VPWR
rlabel comment 17644 13264 17644 13264 8 sr_0.hold1.dlygate4sd3_1
rlabel metal1 16908 13216 17644 13312 5 sr_0.hold1.VGND
rlabel metal1 16908 12672 17644 12768 5 sr_0.hold1.VPWR
flabel locali 17397 12465 17431 12499 0 FreeSans 200 0 0 0 sr_0.output5.X
flabel locali 17121 12329 17155 12363 0 FreeSans 200 0 0 0 sr_0.output5.A
flabel locali 17489 12329 17523 12363 0 FreeSans 200 0 0 0 sr_0.output5.X
flabel locali 17121 12397 17155 12431 0 FreeSans 200 0 0 0 sr_0.output5.A
flabel locali 17489 12397 17523 12431 0 FreeSans 200 0 0 0 sr_0.output5.X
flabel metal1 17029 12159 17063 12193 0 FreeSans 200 0 0 0 sr_0.output5.VGND
flabel metal1 17029 12703 17063 12737 0 FreeSans 200 0 0 0 sr_0.output5.VPWR
flabel nwell 17029 12703 17063 12737 0 FreeSans 200 0 0 0 sr_0.output5.VPB
flabel pwell 17029 12159 17063 12193 0 FreeSans 200 0 0 0 sr_0.output5.VNB
rlabel comment 17000 12176 17000 12176 4 sr_0.output5.clkbuf_4
rlabel metal1 17000 12128 17552 12224 1 sr_0.output5.VGND
rlabel metal1 17000 12672 17552 12768 1 sr_0.output5.VPWR
flabel metal1 14903 12162 14956 12194 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_57.VGND
flabel metal1 14903 12706 14955 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_57.VPWR
flabel nwell 14914 12711 14948 12729 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_57.VPB
flabel pwell 14913 12166 14945 12188 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_57.VNB
rlabel comment 14976 12176 14976 12176 6 sr_0.FILLER_0_0_57.fill_2
rlabel metal1 14792 12128 14976 12224 1 sr_0.FILLER_0_0_57.VGND
rlabel metal1 14792 12672 14976 12768 1 sr_0.FILLER_0_0_57.VPWR
flabel metal1 14918 12707 14954 12737 0 FreeSans 250 0 0 0 sr_0.FILLER_0_1_57.VPWR
flabel metal1 14918 13248 14954 13277 0 FreeSans 250 0 0 0 sr_0.FILLER_0_1_57.VGND
flabel nwell 14925 12713 14945 12730 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_57.VPB
flabel pwell 14924 13253 14948 13275 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_57.VNB
rlabel comment 14976 13264 14976 13264 8 sr_0.FILLER_0_1_57.fill_1
rlabel metal1 14884 13216 14976 13312 5 sr_0.FILLER_0_1_57.VGND
rlabel metal1 14884 12672 14976 12768 5 sr_0.FILLER_0_1_57.VPWR
flabel metal1 14993 12700 15046 12729 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_0_57.VPWR
flabel metal1 14996 12158 15047 12196 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_0_57.VGND
rlabel comment 15068 12176 15068 12176 6 sr_0.TAP_TAPCELL_ROW_0_57.tapvpwrvgnd_1
rlabel metal1 14976 12128 15068 12224 1 sr_0.TAP_TAPCELL_ROW_0_57.VGND
rlabel metal1 14976 12672 15068 12768 1 sr_0.TAP_TAPCELL_ROW_0_57.VPWR
flabel metal1 14993 12711 15046 12740 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_1_61.VPWR
flabel metal1 14996 13244 15047 13282 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_1_61.VGND
rlabel comment 15068 13264 15068 13264 8 sr_0.TAP_TAPCELL_ROW_1_61.tapvpwrvgnd_1
rlabel metal1 14976 13216 15068 13312 5 sr_0.TAP_TAPCELL_ROW_1_61.VGND
rlabel metal1 14976 12672 15068 12768 5 sr_0.TAP_TAPCELL_ROW_1_61.VPWR
flabel metal1 14086 13247 14120 13281 0 FreeSans 200 0 0 0 sr_0._18_.VGND
flabel metal1 14086 12703 14120 12737 0 FreeSans 200 0 0 0 sr_0._18_.VPWR
flabel locali 14730 12941 14764 12975 0 FreeSans 250 0 0 0 sr_0._18_.S
flabel locali 14638 12941 14672 12975 0 FreeSans 250 0 0 0 sr_0._18_.S
flabel locali 14546 13077 14580 13111 0 FreeSans 250 0 0 0 sr_0._18_.A1
flabel locali 14546 13009 14580 13043 0 FreeSans 250 0 0 0 sr_0._18_.A1
flabel locali 14454 13009 14488 13043 0 FreeSans 250 0 0 0 sr_0._18_.A0
flabel locali 14086 13145 14120 13179 0 FreeSans 250 0 0 0 sr_0._18_.X
flabel locali 14086 12873 14120 12907 0 FreeSans 250 0 0 0 sr_0._18_.X
flabel locali 14086 12805 14120 12839 0 FreeSans 250 0 0 0 sr_0._18_.X
flabel nwell 14130 12703 14164 12737 0 FreeSans 250 0 0 0 sr_0._18_.VPB
flabel pwell 14140 13247 14174 13281 0 FreeSans 250 0 0 0 sr_0._18_.VNB
rlabel comment 14056 13264 14056 13264 2 sr_0._18_.mux2_1
rlabel metal1 14056 13216 14884 13312 5 sr_0._18_.VGND
rlabel metal1 14056 12672 14884 12768 5 sr_0._18_.VPWR
flabel locali 14085 12397 14119 12431 0 FreeSans 200 0 0 0 sr_0.hold6.A
flabel locali 14733 12329 14767 12363 0 FreeSans 200 0 0 0 sr_0.hold6.X
flabel locali 14085 12465 14119 12499 0 FreeSans 200 0 0 0 sr_0.hold6.A
flabel locali 14733 12261 14767 12295 0 FreeSans 200 0 0 0 sr_0.hold6.X
flabel locali 14177 12397 14211 12431 0 FreeSans 200 0 0 0 sr_0.hold6.A
flabel locali 14177 12465 14211 12499 0 FreeSans 200 0 0 0 sr_0.hold6.A
flabel locali 14733 12601 14767 12635 0 FreeSans 200 0 0 0 sr_0.hold6.X
flabel locali 14733 12465 14767 12499 0 FreeSans 200 0 0 0 sr_0.hold6.X
flabel locali 14733 12533 14767 12567 0 FreeSans 200 0 0 0 sr_0.hold6.X
flabel locali 14733 12397 14767 12431 0 FreeSans 200 0 0 0 sr_0.hold6.X
flabel nwell 14085 12703 14119 12737 0 FreeSans 200 0 0 0 sr_0.hold6.VPB
flabel pwell 14085 12159 14119 12193 0 FreeSans 200 0 0 0 sr_0.hold6.VNB
flabel metal1 14085 12159 14119 12193 0 FreeSans 200 0 0 0 sr_0.hold6.VGND
flabel metal1 14085 12703 14119 12737 0 FreeSans 200 0 0 0 sr_0.hold6.VPWR
rlabel comment 14056 12176 14056 12176 4 sr_0.hold6.dlygate4sd3_1
rlabel metal1 14056 12128 14792 12224 1 sr_0.hold6.VGND
rlabel metal1 14056 12672 14792 12768 1 sr_0.hold6.VPWR
flabel metal1 12603 12162 12656 12194 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_82.VGND
flabel metal1 12603 12706 12655 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_82.VPWR
flabel nwell 12614 12711 12648 12729 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_82.VPB
flabel pwell 12613 12166 12645 12188 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_82.VNB
rlabel comment 12676 12176 12676 12176 6 sr_0.FILLER_0_0_82.fill_2
rlabel metal1 12492 12128 12676 12224 1 sr_0.FILLER_0_0_82.VGND
rlabel metal1 12492 12672 12676 12768 1 sr_0.FILLER_0_0_82.VPWR
flabel metal1 13809 12159 13843 12193 0 FreeSans 200 180 0 0 sr_0._21_.VGND
flabel metal1 13809 12703 13843 12737 0 FreeSans 200 180 0 0 sr_0._21_.VPWR
flabel locali 13993 12261 14027 12295 0 FreeSans 200 180 0 0 sr_0._21_.X
flabel locali 13993 12533 14027 12567 0 FreeSans 200 180 0 0 sr_0._21_.X
flabel locali 13993 12601 14027 12635 0 FreeSans 200 180 0 0 sr_0._21_.X
flabel locali 13809 12397 13843 12431 0 FreeSans 200 180 0 0 sr_0._21_.A
flabel nwell 13809 12703 13843 12737 0 FreeSans 200 180 0 0 sr_0._21_.VPB
flabel pwell 13809 12159 13843 12193 0 FreeSans 200 180 0 0 sr_0._21_.VNB
rlabel comment 14056 12176 14056 12176 6 sr_0._21_.clkbuf_1
rlabel metal1 13780 12128 14056 12224 1 sr_0._21_.VGND
rlabel metal1 13780 12672 14056 12768 1 sr_0._21_.VPWR
flabel locali 13992 12805 14026 12839 0 FreeSans 400 0 0 0 sr_0._32_.Q
flabel locali 13992 12873 14026 12907 0 FreeSans 400 0 0 0 sr_0._32_.Q
flabel locali 13992 12941 14026 12975 0 FreeSans 400 0 0 0 sr_0._32_.Q
flabel locali 13992 13145 14026 13179 0 FreeSans 400 0 0 0 sr_0._32_.Q
flabel locali 13697 13077 13731 13111 0 FreeSans 400 0 0 0 sr_0._32_.RESET_B
flabel locali 12521 12941 12555 12975 0 FreeSans 400 0 0 0 sr_0._32_.D
flabel locali 12246 12941 12280 12975 0 FreeSans 400 0 0 0 sr_0._32_.CLK
flabel locali 12246 13009 12280 13043 0 FreeSans 400 0 0 0 sr_0._32_.CLK
flabel locali 13697 13009 13731 13043 0 FreeSans 400 0 0 0 sr_0._32_.RESET_B
flabel metal1 12245 13247 12279 13281 0 FreeSans 200 0 0 0 sr_0._32_.VGND
flabel metal1 12245 12703 12279 12737 0 FreeSans 200 0 0 0 sr_0._32_.VPWR
flabel nwell 12245 12703 12279 12737 0 FreeSans 200 0 0 0 sr_0._32_.VPB
flabel pwell 12245 13247 12279 13281 0 FreeSans 200 0 0 0 sr_0._32_.VNB
rlabel comment 12216 13264 12216 13264 2 sr_0._32_.dfrtp_1
rlabel locali 13697 13057 13745 13137 5 sr_0._32_.RESET_B
rlabel locali 13637 12983 13745 13057 5 sr_0._32_.RESET_B
rlabel metal1 13685 13108 13743 13117 5 sr_0._32_.RESET_B
rlabel metal1 13625 13008 13683 13071 5 sr_0._32_.RESET_B
rlabel metal1 13625 13071 13743 13080 5 sr_0._32_.RESET_B
rlabel metal1 12965 13071 13095 13080 5 sr_0._32_.RESET_B
rlabel metal1 12965 13080 13743 13108 5 sr_0._32_.RESET_B
rlabel metal1 12965 13108 13095 13117 5 sr_0._32_.RESET_B
rlabel metal1 12216 13216 14056 13312 5 sr_0._32_.VGND
rlabel metal1 12216 12672 14056 12768 5 sr_0._32_.VPWR
flabel locali 12797 12465 12831 12499 0 FreeSans 200 0 0 0 sr_0.output6.X
flabel locali 13073 12329 13107 12363 0 FreeSans 200 0 0 0 sr_0.output6.A
flabel locali 12705 12329 12739 12363 0 FreeSans 200 0 0 0 sr_0.output6.X
flabel locali 13073 12397 13107 12431 0 FreeSans 200 0 0 0 sr_0.output6.A
flabel locali 12705 12397 12739 12431 0 FreeSans 200 0 0 0 sr_0.output6.X
flabel metal1 13165 12159 13199 12193 0 FreeSans 200 0 0 0 sr_0.output6.VGND
flabel metal1 13165 12703 13199 12737 0 FreeSans 200 0 0 0 sr_0.output6.VPWR
flabel nwell 13165 12703 13199 12737 0 FreeSans 200 0 0 0 sr_0.output6.VPB
flabel pwell 13165 12159 13199 12193 0 FreeSans 200 0 0 0 sr_0.output6.VNB
rlabel comment 13228 12176 13228 12176 6 sr_0.output6.clkbuf_4
rlabel metal1 12676 12128 13228 12224 1 sr_0.output6.VGND
rlabel metal1 12676 12672 13228 12768 1 sr_0.output6.VPWR
flabel locali 13625 12465 13659 12499 0 FreeSans 200 0 0 0 sr_0.output7.X
flabel locali 13349 12329 13383 12363 0 FreeSans 200 0 0 0 sr_0.output7.A
flabel locali 13717 12329 13751 12363 0 FreeSans 200 0 0 0 sr_0.output7.X
flabel locali 13349 12397 13383 12431 0 FreeSans 200 0 0 0 sr_0.output7.A
flabel locali 13717 12397 13751 12431 0 FreeSans 200 0 0 0 sr_0.output7.X
flabel metal1 13257 12159 13291 12193 0 FreeSans 200 0 0 0 sr_0.output7.VGND
flabel metal1 13257 12703 13291 12737 0 FreeSans 200 0 0 0 sr_0.output7.VPWR
flabel nwell 13257 12703 13291 12737 0 FreeSans 200 0 0 0 sr_0.output7.VPB
flabel pwell 13257 12159 13291 12193 0 FreeSans 200 0 0 0 sr_0.output7.VNB
rlabel comment 13228 12176 13228 12176 4 sr_0.output7.clkbuf_4
rlabel metal1 13228 12128 13780 12224 1 sr_0.output7.VGND
rlabel metal1 13228 12672 13780 12768 1 sr_0.output7.VPWR
flabel metal1 12327 12162 12380 12194 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_85.VGND
flabel metal1 12327 12706 12379 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_85.VPWR
flabel nwell 12338 12711 12372 12729 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_85.VPB
flabel pwell 12337 12166 12369 12188 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_85.VNB
rlabel comment 12400 12176 12400 12176 6 sr_0.FILLER_0_0_85.fill_2
rlabel metal1 12216 12128 12400 12224 1 sr_0.FILLER_0_0_85.VGND
rlabel metal1 12216 12672 12400 12768 1 sr_0.FILLER_0_0_85.VPWR
flabel metal1 11330 12703 11366 12733 0 FreeSans 250 0 0 0 sr_0.FILLER_0_0_96.VPWR
flabel metal1 11330 12163 11366 12192 0 FreeSans 250 0 0 0 sr_0.FILLER_0_0_96.VGND
flabel nwell 11337 12710 11357 12727 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_96.VPB
flabel pwell 11336 12165 11360 12187 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_96.VNB
rlabel comment 11388 12176 11388 12176 6 sr_0.FILLER_0_0_96.fill_1
rlabel metal1 11296 12128 11388 12224 1 sr_0.FILLER_0_0_96.VGND
rlabel metal1 11296 12672 11388 12768 1 sr_0.FILLER_0_0_96.VPWR
flabel metal1 12417 12700 12470 12729 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_0_58.VPWR
flabel metal1 12420 12158 12471 12196 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_0_58.VGND
rlabel comment 12492 12176 12492 12176 6 sr_0.TAP_TAPCELL_ROW_0_58.tapvpwrvgnd_1
rlabel metal1 12400 12128 12492 12224 1 sr_0.TAP_TAPCELL_ROW_0_58.VGND
rlabel metal1 12400 12672 12492 12768 1 sr_0.TAP_TAPCELL_ROW_0_58.VPWR
flabel metal1 12152 12159 12186 12193 0 FreeSans 200 0 0 0 sr_0._22_.VGND
flabel metal1 12152 12703 12186 12737 0 FreeSans 200 0 0 0 sr_0._22_.VPWR
flabel locali 11508 12465 11542 12499 0 FreeSans 250 0 0 0 sr_0._22_.S
flabel locali 11600 12465 11634 12499 0 FreeSans 250 0 0 0 sr_0._22_.S
flabel locali 11692 12329 11726 12363 0 FreeSans 250 0 0 0 sr_0._22_.A1
flabel locali 11692 12397 11726 12431 0 FreeSans 250 0 0 0 sr_0._22_.A1
flabel locali 11784 12397 11818 12431 0 FreeSans 250 0 0 0 sr_0._22_.A0
flabel locali 12152 12261 12186 12295 0 FreeSans 250 0 0 0 sr_0._22_.X
flabel locali 12152 12533 12186 12567 0 FreeSans 250 0 0 0 sr_0._22_.X
flabel locali 12152 12601 12186 12635 0 FreeSans 250 0 0 0 sr_0._22_.X
flabel nwell 12108 12703 12142 12737 0 FreeSans 250 0 0 0 sr_0._22_.VPB
flabel pwell 12098 12159 12132 12193 0 FreeSans 250 0 0 0 sr_0._22_.VNB
rlabel comment 12216 12176 12216 12176 6 sr_0._22_.mux2_1
rlabel metal1 11388 12128 12216 12224 1 sr_0._22_.VGND
rlabel metal1 11388 12672 12216 12768 1 sr_0._22_.VPWR
flabel metal1 10498 12159 10532 12193 0 FreeSans 200 0 0 0 sr_0._24_.VGND
flabel metal1 10498 12703 10532 12737 0 FreeSans 200 0 0 0 sr_0._24_.VPWR
flabel locali 11142 12465 11176 12499 0 FreeSans 250 0 0 0 sr_0._24_.S
flabel locali 11050 12465 11084 12499 0 FreeSans 250 0 0 0 sr_0._24_.S
flabel locali 10958 12329 10992 12363 0 FreeSans 250 0 0 0 sr_0._24_.A1
flabel locali 10958 12397 10992 12431 0 FreeSans 250 0 0 0 sr_0._24_.A1
flabel locali 10866 12397 10900 12431 0 FreeSans 250 0 0 0 sr_0._24_.A0
flabel locali 10498 12261 10532 12295 0 FreeSans 250 0 0 0 sr_0._24_.X
flabel locali 10498 12533 10532 12567 0 FreeSans 250 0 0 0 sr_0._24_.X
flabel locali 10498 12601 10532 12635 0 FreeSans 250 0 0 0 sr_0._24_.X
flabel nwell 10542 12703 10576 12737 0 FreeSans 250 0 0 0 sr_0._24_.VPB
flabel pwell 10552 12159 10586 12193 0 FreeSans 250 0 0 0 sr_0._24_.VNB
rlabel comment 10468 12176 10468 12176 4 sr_0._24_.mux2_1
rlabel metal1 10468 12128 11296 12224 1 sr_0._24_.VGND
rlabel metal1 10468 12672 11296 12768 1 sr_0._24_.VPWR
flabel locali 10406 12805 10440 12839 0 FreeSans 400 0 0 0 sr_0._33_.Q
flabel locali 10406 12873 10440 12907 0 FreeSans 400 0 0 0 sr_0._33_.Q
flabel locali 10406 12941 10440 12975 0 FreeSans 400 0 0 0 sr_0._33_.Q
flabel locali 10406 13145 10440 13179 0 FreeSans 400 0 0 0 sr_0._33_.Q
flabel locali 10701 13077 10735 13111 0 FreeSans 400 0 0 0 sr_0._33_.RESET_B
flabel locali 11877 12941 11911 12975 0 FreeSans 400 0 0 0 sr_0._33_.D
flabel locali 12152 12941 12186 12975 0 FreeSans 400 0 0 0 sr_0._33_.CLK
flabel locali 12152 13009 12186 13043 0 FreeSans 400 0 0 0 sr_0._33_.CLK
flabel locali 10701 13009 10735 13043 0 FreeSans 400 0 0 0 sr_0._33_.RESET_B
flabel metal1 12153 13247 12187 13281 0 FreeSans 200 0 0 0 sr_0._33_.VGND
flabel metal1 12153 12703 12187 12737 0 FreeSans 200 0 0 0 sr_0._33_.VPWR
flabel nwell 12153 12703 12187 12737 0 FreeSans 200 0 0 0 sr_0._33_.VPB
flabel pwell 12153 13247 12187 13281 0 FreeSans 200 0 0 0 sr_0._33_.VNB
rlabel comment 12216 13264 12216 13264 8 sr_0._33_.dfrtp_1
rlabel locali 10687 13057 10735 13137 5 sr_0._33_.RESET_B
rlabel locali 10687 12983 10795 13057 5 sr_0._33_.RESET_B
rlabel metal1 10689 13108 10747 13117 5 sr_0._33_.RESET_B
rlabel metal1 10749 13008 10807 13071 5 sr_0._33_.RESET_B
rlabel metal1 10689 13071 10807 13080 5 sr_0._33_.RESET_B
rlabel metal1 11337 13071 11467 13080 5 sr_0._33_.RESET_B
rlabel metal1 10689 13080 11467 13108 5 sr_0._33_.RESET_B
rlabel metal1 11337 13108 11467 13117 5 sr_0._33_.RESET_B
rlabel metal1 10376 13216 12216 13312 5 sr_0._33_.VGND
rlabel metal1 10376 12672 12216 12768 5 sr_0._33_.VPWR
flabel locali 10037 12465 10071 12499 0 FreeSans 200 0 0 0 sr_0.output8.X
flabel locali 10313 12329 10347 12363 0 FreeSans 200 0 0 0 sr_0.output8.A
flabel locali 9945 12329 9979 12363 0 FreeSans 200 0 0 0 sr_0.output8.X
flabel locali 10313 12397 10347 12431 0 FreeSans 200 0 0 0 sr_0.output8.A
flabel locali 9945 12397 9979 12431 0 FreeSans 200 0 0 0 sr_0.output8.X
flabel metal1 10405 12159 10439 12193 0 FreeSans 200 0 0 0 sr_0.output8.VGND
flabel metal1 10405 12703 10439 12737 0 FreeSans 200 0 0 0 sr_0.output8.VPWR
flabel nwell 10405 12703 10439 12737 0 FreeSans 200 0 0 0 sr_0.output8.VPB
flabel pwell 10405 12159 10439 12193 0 FreeSans 200 0 0 0 sr_0.output8.VNB
rlabel comment 10468 12176 10468 12176 6 sr_0.output8.clkbuf_4
rlabel metal1 9916 12128 10468 12224 1 sr_0.output8.VGND
rlabel metal1 9916 12672 10468 12768 1 sr_0.output8.VPWR
flabel locali 9117 13009 9151 13043 0 FreeSans 200 0 0 0 sr_0.hold5.A
flabel locali 9765 13077 9799 13111 0 FreeSans 200 0 0 0 sr_0.hold5.X
flabel locali 9117 12941 9151 12975 0 FreeSans 200 0 0 0 sr_0.hold5.A
flabel locali 9765 13145 9799 13179 0 FreeSans 200 0 0 0 sr_0.hold5.X
flabel locali 9209 13009 9243 13043 0 FreeSans 200 0 0 0 sr_0.hold5.A
flabel locali 9209 12941 9243 12975 0 FreeSans 200 0 0 0 sr_0.hold5.A
flabel locali 9765 12805 9799 12839 0 FreeSans 200 0 0 0 sr_0.hold5.X
flabel locali 9765 12941 9799 12975 0 FreeSans 200 0 0 0 sr_0.hold5.X
flabel locali 9765 12873 9799 12907 0 FreeSans 200 0 0 0 sr_0.hold5.X
flabel locali 9765 13009 9799 13043 0 FreeSans 200 0 0 0 sr_0.hold5.X
flabel nwell 9117 12703 9151 12737 0 FreeSans 200 0 0 0 sr_0.hold5.VPB
flabel pwell 9117 13247 9151 13281 0 FreeSans 200 0 0 0 sr_0.hold5.VNB
flabel metal1 9117 13247 9151 13281 0 FreeSans 200 0 0 0 sr_0.hold5.VGND
flabel metal1 9117 12703 9151 12737 0 FreeSans 200 0 0 0 sr_0.hold5.VPWR
rlabel comment 9088 13264 9088 13264 2 sr_0.hold5.dlygate4sd3_1
rlabel metal1 9088 13216 9824 13312 5 sr_0.hold5.VGND
rlabel metal1 9088 12672 9824 12768 5 sr_0.hold5.VPWR
flabel metal1 9841 12711 9894 12740 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_1_62.VPWR
flabel metal1 9844 13244 9895 13282 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_1_62.VGND
rlabel comment 9916 13264 9916 13264 8 sr_0.TAP_TAPCELL_ROW_1_62.tapvpwrvgnd_1
rlabel metal1 9824 13216 9916 13312 5 sr_0.TAP_TAPCELL_ROW_1_62.VGND
rlabel metal1 9824 12672 9916 12768 5 sr_0.TAP_TAPCELL_ROW_1_62.VPWR
flabel metal1 9841 12700 9894 12729 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_0_59.VPWR
flabel metal1 9844 12158 9895 12196 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_0_59.VGND
rlabel comment 9916 12176 9916 12176 6 sr_0.TAP_TAPCELL_ROW_0_59.tapvpwrvgnd_1
rlabel metal1 9824 12128 9916 12224 1 sr_0.TAP_TAPCELL_ROW_0_59.VGND
rlabel metal1 9824 12672 9916 12768 1 sr_0.TAP_TAPCELL_ROW_0_59.VPWR
flabel metal1 9950 12707 9986 12737 0 FreeSans 250 0 0 0 sr_0.FILLER_0_1_111.VPWR
flabel metal1 9950 13248 9986 13277 0 FreeSans 250 0 0 0 sr_0.FILLER_0_1_111.VGND
flabel nwell 9957 12713 9977 12730 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_111.VPB
flabel pwell 9956 13253 9980 13275 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_111.VNB
rlabel comment 10008 13264 10008 13264 8 sr_0.FILLER_0_1_111.fill_1
rlabel metal1 9916 13216 10008 13312 5 sr_0.FILLER_0_1_111.VGND
rlabel metal1 9916 12672 10008 12768 5 sr_0.FILLER_0_1_111.VPWR
flabel metal1 10313 13247 10347 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_107.VGND
flabel metal1 10313 12703 10347 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_107.VPWR
flabel nwell 10313 12703 10347 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_107.VPB
flabel pwell 10313 13247 10347 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_107.VNB
rlabel comment 10376 13264 10376 13264 8 sr_0.FILLER_0_1_107.decap_4
rlabel metal1 10008 13216 10376 13312 5 sr_0.FILLER_0_1_107.VGND
rlabel metal1 10008 12672 10376 12768 5 sr_0.FILLER_0_1_107.VPWR
flabel metal1 9761 12159 9795 12193 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_113.VGND
flabel metal1 9761 12703 9795 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_113.VPWR
flabel nwell 9761 12703 9795 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_113.VPB
flabel pwell 9761 12159 9795 12193 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_113.VNB
rlabel comment 9824 12176 9824 12176 6 sr_0.FILLER_0_0_113.decap_4
rlabel metal1 9456 12128 9824 12224 1 sr_0.FILLER_0_0_113.VGND
rlabel metal1 9456 12672 9824 12768 1 sr_0.FILLER_0_0_113.VPWR
flabel locali 8933 12465 8967 12499 0 FreeSans 200 0 0 0 sr_0.output9.X
flabel locali 9209 12329 9243 12363 0 FreeSans 200 0 0 0 sr_0.output9.A
flabel locali 8841 12329 8875 12363 0 FreeSans 200 0 0 0 sr_0.output9.X
flabel locali 9209 12397 9243 12431 0 FreeSans 200 0 0 0 sr_0.output9.A
flabel locali 8841 12397 8875 12431 0 FreeSans 200 0 0 0 sr_0.output9.X
flabel metal1 9301 12159 9335 12193 0 FreeSans 200 0 0 0 sr_0.output9.VGND
flabel metal1 9301 12703 9335 12737 0 FreeSans 200 0 0 0 sr_0.output9.VPWR
flabel nwell 9301 12703 9335 12737 0 FreeSans 200 0 0 0 sr_0.output9.VPB
flabel pwell 9301 12159 9335 12193 0 FreeSans 200 0 0 0 sr_0.output9.VNB
rlabel comment 9364 12176 9364 12176 6 sr_0.output9.clkbuf_4
rlabel metal1 8812 12128 9364 12224 1 sr_0.output9.VGND
rlabel metal1 8812 12672 9364 12768 1 sr_0.output9.VPWR
flabel metal1 9398 12703 9434 12733 0 FreeSans 250 0 0 0 sr_0.FILLER_0_0_117.VPWR
flabel metal1 9398 12163 9434 12192 0 FreeSans 250 0 0 0 sr_0.FILLER_0_0_117.VGND
flabel nwell 9405 12710 9425 12727 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_117.VPB
flabel pwell 9404 12165 9428 12187 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_117.VNB
rlabel comment 9456 12176 9456 12176 6 sr_0.FILLER_0_0_117.fill_1
rlabel metal1 9364 12128 9456 12224 1 sr_0.FILLER_0_0_117.VGND
rlabel metal1 9364 12672 9456 12768 1 sr_0.FILLER_0_0_117.VPWR
flabel metal1 9025 13247 9059 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_121.VGND
flabel metal1 9025 12703 9059 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_121.VPWR
flabel nwell 9025 12703 9059 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_121.VPB
flabel pwell 9025 13247 9059 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_121.VNB
rlabel comment 9088 13264 9088 13264 8 sr_0.FILLER_0_1_121.decap_12
flabel metal1 8749 12159 8783 12193 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_124.VGND
flabel metal1 8749 12703 8783 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_124.VPWR
flabel nwell 8749 12703 8783 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_124.VPB
flabel pwell 8749 12159 8783 12193 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_124.VNB
rlabel comment 8812 12176 8812 12176 6 sr_0.FILLER_0_0_124.decap_12
flabel metal1 7645 12159 7679 12193 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_136.VGND
flabel metal1 7645 12703 7679 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_136.VPWR
flabel nwell 7645 12703 7679 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_136.VPB
flabel pwell 7645 12159 7679 12193 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_136.VNB
rlabel comment 7708 12176 7708 12176 6 sr_0.FILLER_0_0_136.decap_4
rlabel metal1 7340 12128 7708 12224 1 sr_0.FILLER_0_0_136.VGND
rlabel metal1 7340 12672 7708 12768 1 sr_0.FILLER_0_0_136.VPWR
flabel metal1 7921 13247 7955 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_133.VGND
flabel metal1 7921 12703 7955 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_133.VPWR
flabel nwell 7921 12703 7955 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_133.VPB
flabel pwell 7921 13247 7955 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_133.VNB
rlabel comment 7984 13264 7984 13264 8 sr_0.FILLER_0_1_133.decap_12
flabel metal1 6817 13247 6851 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_145.VGND
flabel metal1 6817 12703 6851 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_145.VPWR
flabel nwell 6817 12703 6851 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_145.VPB
flabel pwell 6817 13247 6851 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_145.VNB
rlabel comment 6880 13264 6880 13264 8 sr_0.FILLER_0_1_145.decap_12
flabel metal1 7265 12700 7318 12729 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_0_60.VPWR
flabel metal1 7268 12158 7319 12196 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_0_60.VGND
rlabel comment 7340 12176 7340 12176 6 sr_0.TAP_TAPCELL_ROW_0_60.tapvpwrvgnd_1
rlabel metal1 7248 12128 7340 12224 1 sr_0.TAP_TAPCELL_ROW_0_60.VGND
rlabel metal1 7248 12672 7340 12768 1 sr_0.TAP_TAPCELL_ROW_0_60.VPWR
flabel locali 6817 12465 6851 12499 0 FreeSans 200 0 0 0 sr_0.output10.X
flabel locali 7093 12329 7127 12363 0 FreeSans 200 0 0 0 sr_0.output10.A
flabel locali 6725 12329 6759 12363 0 FreeSans 200 0 0 0 sr_0.output10.X
flabel locali 7093 12397 7127 12431 0 FreeSans 200 0 0 0 sr_0.output10.A
flabel locali 6725 12397 6759 12431 0 FreeSans 200 0 0 0 sr_0.output10.X
flabel metal1 7185 12159 7219 12193 0 FreeSans 200 0 0 0 sr_0.output10.VGND
flabel metal1 7185 12703 7219 12737 0 FreeSans 200 0 0 0 sr_0.output10.VPWR
flabel nwell 7185 12703 7219 12737 0 FreeSans 200 0 0 0 sr_0.output10.VPB
flabel pwell 7185 12159 7219 12193 0 FreeSans 200 0 0 0 sr_0.output10.VNB
rlabel comment 7248 12176 7248 12176 6 sr_0.output10.clkbuf_4
rlabel metal1 6696 12128 7248 12224 1 sr_0.output10.VGND
rlabel metal1 6696 12672 7248 12768 1 sr_0.output10.VPWR
flabel metal1 6633 12159 6667 12193 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_147.VGND
flabel metal1 6633 12703 6667 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_147.VPWR
flabel nwell 6633 12703 6667 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_147.VPB
flabel pwell 6633 12159 6667 12193 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_147.VNB
rlabel comment 6696 12176 6696 12176 6 sr_0.FILLER_0_0_147.decap_12
flabel metal1 5534 12703 5570 12733 0 FreeSans 250 0 0 0 sr_0.FILLER_0_0_159.VPWR
flabel metal1 5534 12163 5570 12192 0 FreeSans 250 0 0 0 sr_0.FILLER_0_0_159.VGND
flabel nwell 5541 12710 5561 12727 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_159.VPB
flabel pwell 5540 12165 5564 12187 0 FreeSans 200 0 0 0 sr_0.FILLER_0_0_159.VNB
rlabel comment 5592 12176 5592 12176 6 sr_0.FILLER_0_0_159.fill_1
rlabel metal1 5500 12128 5592 12224 1 sr_0.FILLER_0_0_159.VGND
rlabel metal1 5500 12672 5592 12768 1 sr_0.FILLER_0_0_159.VPWR
flabel metal1 5713 12703 5747 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_157.VPWR
flabel metal1 5713 13247 5747 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_157.VGND
flabel nwell 5713 12703 5747 12737 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_157.VPB
flabel pwell 5713 13247 5747 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_1_157.VNB
rlabel comment 5776 13264 5776 13264 8 sr_0.FILLER_0_1_157.decap_6
rlabel metal1 5224 13216 5776 13312 5 sr_0.FILLER_0_1_157.VGND
rlabel metal1 5224 12672 5776 12768 5 sr_0.FILLER_0_1_157.VPWR
flabel metal1 4977 12703 5011 12737 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_0_Right_0.VPWR
flabel metal1 4977 12159 5011 12193 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_0_Right_0.VGND
flabel nwell 4977 12703 5011 12737 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_0_Right_0.VPB
flabel pwell 4977 12159 5011 12193 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_0_Right_0.VNB
rlabel comment 4948 12176 4948 12176 4 sr_0.PHY_EDGE_ROW_0_Right_0.decap_3
rlabel metal1 4948 12128 5224 12224 1 sr_0.PHY_EDGE_ROW_0_Right_0.VGND
rlabel metal1 4948 12672 5224 12768 1 sr_0.PHY_EDGE_ROW_0_Right_0.VPWR
flabel metal1 4977 12703 5011 12737 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_1_Right_1.VPWR
flabel metal1 4977 13247 5011 13281 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_1_Right_1.VGND
flabel nwell 4977 12703 5011 12737 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_1_Right_1.VPB
flabel pwell 4977 13247 5011 13281 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_1_Right_1.VNB
rlabel comment 4948 13264 4948 13264 2 sr_0.PHY_EDGE_ROW_1_Right_1.decap_3
rlabel metal1 4948 13216 5224 13312 5 sr_0.PHY_EDGE_ROW_1_Right_1.VGND
rlabel metal1 4948 12672 5224 12768 5 sr_0.PHY_EDGE_ROW_1_Right_1.VPWR
flabel locali 5272 12465 5306 12499 0 FreeSans 200 0 0 0 sr_0.sr_11.LO
flabel locali 5399 12401 5433 12435 0 FreeSans 200 0 0 0 sr_0.sr_11.HI
flabel nwell 5437 12703 5471 12737 0 FreeSans 200 0 0 0 sr_0.sr_11.VPB
flabel pwell 5437 12159 5471 12193 0 FreeSans 200 0 0 0 sr_0.sr_11.VNB
flabel metal1 5437 12159 5471 12193 0 FreeSans 200 0 0 0 sr_0.sr_11.VGND
flabel metal1 5437 12703 5471 12737 0 FreeSans 200 0 0 0 sr_0.sr_11.VPWR
rlabel comment 5500 12176 5500 12176 6 sr_0.sr_11.conb_1
flabel comment 5455 12449 5455 12449 0 FreeSans 200 90 0 0 sr_0.sr_11.resistive_li1_ok
flabel comment 5267 12449 5267 12449 0 FreeSans 200 90 0 0 sr_0.sr_11.resistive_li1_ok
flabel comment 5314 12434 5314 12434 0 FreeSans 200 90 0 0 sr_0.sr_11.no_jumper_check
flabel comment 5417 12434 5417 12434 0 FreeSans 200 90 0 0 sr_0.sr_11.no_jumper_check
rlabel metal1 5224 12128 5500 12224 1 sr_0.sr_11.VGND
rlabel metal1 5224 12672 5500 12768 1 sr_0.sr_11.VPWR
flabel metal1 19881 13247 19915 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_3.VGND
flabel metal1 19881 13791 19915 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_3.VPWR
flabel nwell 19881 13791 19915 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_3.VPB
flabel pwell 19881 13247 19915 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_3.VNB
rlabel comment 19944 13264 19944 13264 6 sr_0.FILLER_0_2_3.decap_12
flabel metal1 18777 13247 18811 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_15.VGND
flabel metal1 18777 13791 18811 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_15.VPWR
flabel nwell 18777 13791 18811 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_15.VPB
flabel pwell 18777 13247 18811 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_15.VNB
rlabel comment 18840 13264 18840 13264 6 sr_0.FILLER_0_2_15.decap_12
flabel metal1 20157 13791 20191 13825 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_2_Left_30.VPWR
flabel metal1 20157 13247 20191 13281 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_2_Left_30.VGND
flabel nwell 20157 13791 20191 13825 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_2_Left_30.VPB
flabel pwell 20157 13247 20191 13281 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_2_Left_30.VNB
rlabel comment 20220 13264 20220 13264 6 sr_0.PHY_EDGE_ROW_2_Left_30.decap_3
rlabel metal1 19944 13216 20220 13312 1 sr_0.PHY_EDGE_ROW_2_Left_30.VGND
rlabel metal1 19944 13760 20220 13856 1 sr_0.PHY_EDGE_ROW_2_Left_30.VPWR
flabel metal1 17678 13791 17714 13821 0 FreeSans 250 0 0 0 sr_0.FILLER_0_2_27.VPWR
flabel metal1 17678 13251 17714 13280 0 FreeSans 250 0 0 0 sr_0.FILLER_0_2_27.VGND
flabel nwell 17685 13798 17705 13815 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_27.VPB
flabel pwell 17684 13253 17708 13275 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_27.VNB
rlabel comment 17736 13264 17736 13264 6 sr_0.FILLER_0_2_27.fill_1
rlabel metal1 17644 13216 17736 13312 1 sr_0.FILLER_0_2_27.VGND
rlabel metal1 17644 13760 17736 13856 1 sr_0.FILLER_0_2_27.VPWR
flabel metal1 17479 13250 17532 13282 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_29.VGND
flabel metal1 17479 13794 17531 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_29.VPWR
flabel nwell 17490 13799 17524 13817 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_29.VPB
flabel pwell 17489 13254 17521 13276 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_29.VNB
rlabel comment 17552 13264 17552 13264 6 sr_0.FILLER_0_2_29.fill_2
rlabel metal1 17368 13216 17552 13312 1 sr_0.FILLER_0_2_29.VGND
rlabel metal1 17368 13760 17552 13856 1 sr_0.FILLER_0_2_29.VPWR
flabel metal1 17569 13788 17622 13817 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_2_63.VPWR
flabel metal1 17572 13246 17623 13284 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_2_63.VGND
rlabel comment 17644 13264 17644 13264 6 sr_0.TAP_TAPCELL_ROW_2_63.tapvpwrvgnd_1
rlabel metal1 17552 13216 17644 13312 1 sr_0.TAP_TAPCELL_ROW_2_63.VGND
rlabel metal1 17552 13760 17644 13856 1 sr_0.TAP_TAPCELL_ROW_2_63.VPWR
flabel metal1 16570 13247 16604 13281 0 FreeSans 200 0 0 0 sr_0._14_.VGND
flabel metal1 16570 13791 16604 13825 0 FreeSans 200 0 0 0 sr_0._14_.VPWR
flabel locali 17214 13553 17248 13587 0 FreeSans 250 0 0 0 sr_0._14_.S
flabel locali 17122 13553 17156 13587 0 FreeSans 250 0 0 0 sr_0._14_.S
flabel locali 17030 13417 17064 13451 0 FreeSans 250 0 0 0 sr_0._14_.A1
flabel locali 17030 13485 17064 13519 0 FreeSans 250 0 0 0 sr_0._14_.A1
flabel locali 16938 13485 16972 13519 0 FreeSans 250 0 0 0 sr_0._14_.A0
flabel locali 16570 13349 16604 13383 0 FreeSans 250 0 0 0 sr_0._14_.X
flabel locali 16570 13621 16604 13655 0 FreeSans 250 0 0 0 sr_0._14_.X
flabel locali 16570 13689 16604 13723 0 FreeSans 250 0 0 0 sr_0._14_.X
flabel nwell 16614 13791 16648 13825 0 FreeSans 250 0 0 0 sr_0._14_.VPB
flabel pwell 16624 13247 16658 13281 0 FreeSans 250 0 0 0 sr_0._14_.VNB
rlabel comment 16540 13264 16540 13264 4 sr_0._14_.mux2_1
rlabel metal1 16540 13216 17368 13312 1 sr_0._14_.VGND
rlabel metal1 16540 13760 17368 13856 1 sr_0._14_.VPWR
flabel locali 16293 13553 16327 13587 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_0__f_sclk.X
flabel locali 16385 13553 16419 13587 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_0__f_sclk.X
flabel locali 16385 13485 16419 13519 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_0__f_sclk.X
flabel locali 16293 13485 16327 13519 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_0__f_sclk.X
flabel locali 16293 13417 16327 13451 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_0__f_sclk.X
flabel locali 16385 13417 16419 13451 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_0__f_sclk.X
flabel locali 14729 13417 14763 13451 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_0__f_sclk.A
flabel locali 14729 13485 14763 13519 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_0__f_sclk.A
flabel pwell 14729 13247 14763 13281 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_0__f_sclk.VNB
flabel pwell 14746 13264 14746 13264 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_0__f_sclk.VNB
flabel nwell 14729 13791 14763 13825 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_0__f_sclk.VPB
flabel nwell 14746 13808 14746 13808 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_0__f_sclk.VPB
flabel metal1 14729 13247 14763 13281 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_0__f_sclk.VGND
flabel metal1 14729 13791 14763 13825 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_0__f_sclk.VPWR
rlabel comment 14700 13264 14700 13264 4 sr_0.clkbuf_1_0__f_sclk.clkbuf_16
rlabel metal1 14700 13216 16540 13312 1 sr_0.clkbuf_1_0__f_sclk.VGND
rlabel metal1 14700 13760 16540 13856 1 sr_0.clkbuf_1_0__f_sclk.VPWR
flabel locali 12890 13689 12924 13723 0 FreeSans 400 0 0 0 sr_0._31_.Q
flabel locali 12890 13621 12924 13655 0 FreeSans 400 0 0 0 sr_0._31_.Q
flabel locali 12890 13553 12924 13587 0 FreeSans 400 0 0 0 sr_0._31_.Q
flabel locali 12890 13349 12924 13383 0 FreeSans 400 0 0 0 sr_0._31_.Q
flabel locali 13185 13417 13219 13451 0 FreeSans 400 0 0 0 sr_0._31_.RESET_B
flabel locali 14361 13553 14395 13587 0 FreeSans 400 0 0 0 sr_0._31_.D
flabel locali 14636 13553 14670 13587 0 FreeSans 400 0 0 0 sr_0._31_.CLK
flabel locali 14636 13485 14670 13519 0 FreeSans 400 0 0 0 sr_0._31_.CLK
flabel locali 13185 13485 13219 13519 0 FreeSans 400 0 0 0 sr_0._31_.RESET_B
flabel metal1 14637 13247 14671 13281 0 FreeSans 200 0 0 0 sr_0._31_.VGND
flabel metal1 14637 13791 14671 13825 0 FreeSans 200 0 0 0 sr_0._31_.VPWR
flabel nwell 14637 13791 14671 13825 0 FreeSans 200 0 0 0 sr_0._31_.VPB
flabel pwell 14637 13247 14671 13281 0 FreeSans 200 0 0 0 sr_0._31_.VNB
rlabel comment 14700 13264 14700 13264 6 sr_0._31_.dfrtp_1
rlabel locali 13171 13391 13219 13471 1 sr_0._31_.RESET_B
rlabel locali 13171 13471 13279 13545 1 sr_0._31_.RESET_B
rlabel metal1 13173 13411 13231 13420 1 sr_0._31_.RESET_B
rlabel metal1 13233 13457 13291 13520 1 sr_0._31_.RESET_B
rlabel metal1 13173 13448 13291 13457 1 sr_0._31_.RESET_B
rlabel metal1 13821 13448 13951 13457 1 sr_0._31_.RESET_B
rlabel metal1 13173 13420 13951 13448 1 sr_0._31_.RESET_B
rlabel metal1 13821 13411 13951 13420 1 sr_0._31_.RESET_B
rlabel metal1 12860 13216 14700 13312 1 sr_0._31_.VGND
rlabel metal1 12860 13760 14700 13856 1 sr_0._31_.VPWR
flabel metal1 12802 13791 12838 13821 0 FreeSans 250 0 0 0 sr_0.FILLER_0_2_80.VPWR
flabel metal1 12802 13251 12838 13280 0 FreeSans 250 0 0 0 sr_0.FILLER_0_2_80.VGND
flabel nwell 12809 13798 12829 13815 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_80.VPB
flabel pwell 12808 13253 12832 13275 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_80.VNB
rlabel comment 12860 13264 12860 13264 6 sr_0.FILLER_0_2_80.fill_1
rlabel metal1 12768 13216 12860 13312 1 sr_0.FILLER_0_2_80.VGND
rlabel metal1 12768 13760 12860 13856 1 sr_0.FILLER_0_2_80.VPWR
flabel metal1 12705 13247 12739 13281 0 FreeSans 200 180 0 0 sr_0._23_.VGND
flabel metal1 12705 13791 12739 13825 0 FreeSans 200 180 0 0 sr_0._23_.VPWR
flabel locali 12521 13349 12555 13383 0 FreeSans 200 180 0 0 sr_0._23_.X
flabel locali 12521 13621 12555 13655 0 FreeSans 200 180 0 0 sr_0._23_.X
flabel locali 12521 13689 12555 13723 0 FreeSans 200 180 0 0 sr_0._23_.X
flabel locali 12705 13485 12739 13519 0 FreeSans 200 180 0 0 sr_0._23_.A
flabel nwell 12705 13791 12739 13825 0 FreeSans 200 180 0 0 sr_0._23_.VPB
flabel pwell 12705 13247 12739 13281 0 FreeSans 200 180 0 0 sr_0._23_.VNB
rlabel comment 12492 13264 12492 13264 4 sr_0._23_.clkbuf_1
rlabel metal1 12492 13216 12768 13312 1 sr_0._23_.VGND
rlabel metal1 12492 13760 12768 13856 1 sr_0._23_.VPWR
flabel metal1 12337 13791 12371 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_85.VPWR
flabel metal1 12337 13247 12371 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_85.VGND
flabel nwell 12337 13791 12371 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_85.VPB
flabel pwell 12337 13247 12371 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_85.VNB
rlabel comment 12400 13264 12400 13264 6 sr_0.FILLER_0_2_85.decap_6
rlabel metal1 11848 13216 12400 13312 1 sr_0.FILLER_0_2_85.VGND
rlabel metal1 11848 13760 12400 13856 1 sr_0.FILLER_0_2_85.VPWR
flabel metal1 11790 13791 11826 13821 0 FreeSans 250 0 0 0 sr_0.FILLER_0_2_91.VPWR
flabel metal1 11790 13251 11826 13280 0 FreeSans 250 0 0 0 sr_0.FILLER_0_2_91.VGND
flabel nwell 11797 13798 11817 13815 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_91.VPB
flabel pwell 11796 13253 11820 13275 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_91.VNB
rlabel comment 11848 13264 11848 13264 6 sr_0.FILLER_0_2_91.fill_1
rlabel metal1 11756 13216 11848 13312 1 sr_0.FILLER_0_2_91.VGND
rlabel metal1 11756 13760 11848 13856 1 sr_0.FILLER_0_2_91.VPWR
flabel metal1 12417 13788 12470 13817 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_2_64.VPWR
flabel metal1 12420 13246 12471 13284 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_2_64.VGND
rlabel comment 12492 13264 12492 13264 6 sr_0.TAP_TAPCELL_ROW_2_64.tapvpwrvgnd_1
rlabel metal1 12400 13216 12492 13312 1 sr_0.TAP_TAPCELL_ROW_2_64.VGND
rlabel metal1 12400 13760 12492 13856 1 sr_0.TAP_TAPCELL_ROW_2_64.VPWR
flabel locali 10129 13553 10163 13587 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_1__f_sclk.X
flabel locali 10037 13553 10071 13587 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_1__f_sclk.X
flabel locali 10037 13485 10071 13519 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_1__f_sclk.X
flabel locali 10129 13485 10163 13519 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_1__f_sclk.X
flabel locali 10129 13417 10163 13451 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_1__f_sclk.X
flabel locali 10037 13417 10071 13451 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_1__f_sclk.X
flabel locali 11693 13417 11727 13451 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_1__f_sclk.A
flabel locali 11693 13485 11727 13519 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_1__f_sclk.A
flabel pwell 11693 13247 11727 13281 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_1__f_sclk.VNB
flabel pwell 11710 13264 11710 13264 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_1__f_sclk.VNB
flabel nwell 11693 13791 11727 13825 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_1__f_sclk.VPB
flabel nwell 11710 13808 11710 13808 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_1__f_sclk.VPB
flabel metal1 11693 13247 11727 13281 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_1__f_sclk.VGND
flabel metal1 11693 13791 11727 13825 0 FreeSans 200 0 0 0 sr_0.clkbuf_1_1__f_sclk.VPWR
rlabel comment 11756 13264 11756 13264 6 sr_0.clkbuf_1_1__f_sclk.clkbuf_16
rlabel metal1 9916 13216 11756 13312 1 sr_0.clkbuf_1_1__f_sclk.VGND
rlabel metal1 9916 13760 11756 13856 1 sr_0.clkbuf_1_1__f_sclk.VPWR
flabel metal1 9577 13247 9611 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_115.VGND
flabel metal1 9577 13791 9611 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_115.VPWR
flabel nwell 9577 13791 9611 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_115.VPB
flabel pwell 9577 13247 9611 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_115.VNB
rlabel comment 9640 13264 9640 13264 6 sr_0.FILLER_0_2_115.decap_12
flabel metal1 9669 13247 9703 13281 0 FreeSans 200 180 0 0 sr_0._25_.VGND
flabel metal1 9669 13791 9703 13825 0 FreeSans 200 180 0 0 sr_0._25_.VPWR
flabel locali 9853 13349 9887 13383 0 FreeSans 200 180 0 0 sr_0._25_.X
flabel locali 9853 13621 9887 13655 0 FreeSans 200 180 0 0 sr_0._25_.X
flabel locali 9853 13689 9887 13723 0 FreeSans 200 180 0 0 sr_0._25_.X
flabel locali 9669 13485 9703 13519 0 FreeSans 200 180 0 0 sr_0._25_.A
flabel nwell 9669 13791 9703 13825 0 FreeSans 200 180 0 0 sr_0._25_.VPB
flabel pwell 9669 13247 9703 13281 0 FreeSans 200 180 0 0 sr_0._25_.VNB
rlabel comment 9916 13264 9916 13264 6 sr_0._25_.clkbuf_1
rlabel metal1 9640 13216 9916 13312 1 sr_0._25_.VGND
rlabel metal1 9640 13760 9916 13856 1 sr_0._25_.VPWR
flabel metal1 8473 13247 8507 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_127.VGND
flabel metal1 8473 13791 8507 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_127.VPWR
flabel nwell 8473 13791 8507 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_127.VPB
flabel pwell 8473 13247 8507 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_127.VNB
rlabel comment 8536 13264 8536 13264 6 sr_0.FILLER_0_2_127.decap_12
flabel metal1 7374 13791 7410 13821 0 FreeSans 250 0 0 0 sr_0.FILLER_0_2_139.VPWR
flabel metal1 7374 13251 7410 13280 0 FreeSans 250 0 0 0 sr_0.FILLER_0_2_139.VGND
flabel nwell 7381 13798 7401 13815 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_139.VPB
flabel pwell 7380 13253 7404 13275 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_139.VNB
rlabel comment 7432 13264 7432 13264 6 sr_0.FILLER_0_2_139.fill_1
rlabel metal1 7340 13216 7432 13312 1 sr_0.FILLER_0_2_139.VGND
rlabel metal1 7340 13760 7432 13856 1 sr_0.FILLER_0_2_139.VPWR
flabel metal1 7185 13247 7219 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_141.VGND
flabel metal1 7185 13791 7219 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_141.VPWR
flabel nwell 7185 13791 7219 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_141.VPB
flabel pwell 7185 13247 7219 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_141.VNB
rlabel comment 7248 13264 7248 13264 6 sr_0.FILLER_0_2_141.decap_12
flabel metal1 7265 13788 7318 13817 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_2_65.VPWR
flabel metal1 7268 13246 7319 13284 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_2_65.VGND
rlabel comment 7340 13264 7340 13264 6 sr_0.TAP_TAPCELL_ROW_2_65.tapvpwrvgnd_1
rlabel metal1 7248 13216 7340 13312 1 sr_0.TAP_TAPCELL_ROW_2_65.VGND
rlabel metal1 7248 13760 7340 13856 1 sr_0.TAP_TAPCELL_ROW_2_65.VPWR
flabel metal1 6081 13791 6115 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_153.VPWR
flabel metal1 6081 13247 6115 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_153.VGND
flabel nwell 6081 13791 6115 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_153.VPB
flabel pwell 6081 13247 6115 13281 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_153.VNB
rlabel comment 6144 13264 6144 13264 6 sr_0.FILLER_0_2_153.decap_8
rlabel metal1 5408 13216 6144 13312 1 sr_0.FILLER_0_2_153.VGND
rlabel metal1 5408 13760 6144 13856 1 sr_0.FILLER_0_2_153.VPWR
flabel metal1 5335 13250 5388 13282 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_161.VGND
flabel metal1 5335 13794 5387 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_161.VPWR
flabel nwell 5346 13799 5380 13817 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_161.VPB
flabel pwell 5345 13254 5377 13276 0 FreeSans 200 0 0 0 sr_0.FILLER_0_2_161.VNB
rlabel comment 5408 13264 5408 13264 6 sr_0.FILLER_0_2_161.fill_2
rlabel metal1 5224 13216 5408 13312 1 sr_0.FILLER_0_2_161.VGND
rlabel metal1 5224 13760 5408 13856 1 sr_0.FILLER_0_2_161.VPWR
flabel metal1 4977 13791 5011 13825 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_2_Right_2.VPWR
flabel metal1 4977 13247 5011 13281 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_2_Right_2.VGND
flabel nwell 4977 13791 5011 13825 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_2_Right_2.VPB
flabel pwell 4977 13247 5011 13281 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_2_Right_2.VNB
rlabel comment 4948 13264 4948 13264 4 sr_0.PHY_EDGE_ROW_2_Right_2.decap_3
rlabel metal1 4948 13216 5224 13312 1 sr_0.PHY_EDGE_ROW_2_Right_2.VGND
rlabel metal1 4948 13760 5224 13856 1 sr_0.PHY_EDGE_ROW_2_Right_2.VPWR
flabel metal1 19881 14335 19915 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_3.VGND
flabel metal1 19881 13791 19915 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_3.VPWR
flabel nwell 19881 13791 19915 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_3.VPB
flabel pwell 19881 14335 19915 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_3.VNB
rlabel comment 19944 14352 19944 14352 8 sr_0.FILLER_0_3_3.decap_12
flabel metal1 18777 14335 18811 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_15.VGND
flabel metal1 18777 13791 18811 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_15.VPWR
flabel nwell 18777 13791 18811 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_15.VPB
flabel pwell 18777 14335 18811 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_15.VNB
rlabel comment 18840 14352 18840 14352 8 sr_0.FILLER_0_3_15.decap_12
flabel metal1 20157 13791 20191 13825 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_3_Left_31.VPWR
flabel metal1 20157 14335 20191 14369 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_3_Left_31.VGND
flabel nwell 20157 13791 20191 13825 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_3_Left_31.VPB
flabel pwell 20157 14335 20191 14369 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_3_Left_31.VNB
rlabel comment 20220 14352 20220 14352 8 sr_0.PHY_EDGE_ROW_3_Left_31.decap_3
rlabel metal1 19944 14304 20220 14400 5 sr_0.PHY_EDGE_ROW_3_Left_31.VGND
rlabel metal1 19944 13760 20220 13856 5 sr_0.PHY_EDGE_ROW_3_Left_31.VPWR
flabel metal1 17673 14335 17707 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_27.VGND
flabel metal1 17673 13791 17707 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_27.VPWR
flabel nwell 17673 13791 17707 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_27.VPB
flabel pwell 17673 14335 17707 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_27.VNB
rlabel comment 17736 14352 17736 14352 8 sr_0.FILLER_0_3_27.decap_12
flabel metal1 16574 13795 16610 13825 0 FreeSans 250 0 0 0 sr_0.FILLER_0_3_39.VPWR
flabel metal1 16574 14336 16610 14365 0 FreeSans 250 0 0 0 sr_0.FILLER_0_3_39.VGND
flabel nwell 16581 13801 16601 13818 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_39.VPB
flabel pwell 16580 14341 16604 14363 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_39.VNB
rlabel comment 16632 14352 16632 14352 8 sr_0.FILLER_0_3_39.fill_1
rlabel metal1 16540 14304 16632 14400 5 sr_0.FILLER_0_3_39.VGND
rlabel metal1 16540 13760 16632 13856 5 sr_0.FILLER_0_3_39.VPWR
flabel metal1 16477 14335 16511 14369 0 FreeSans 200 180 0 0 sr_0._15_.VGND
flabel metal1 16477 13791 16511 13825 0 FreeSans 200 180 0 0 sr_0._15_.VPWR
flabel locali 16293 14233 16327 14267 0 FreeSans 200 180 0 0 sr_0._15_.X
flabel locali 16293 13961 16327 13995 0 FreeSans 200 180 0 0 sr_0._15_.X
flabel locali 16293 13893 16327 13927 0 FreeSans 200 180 0 0 sr_0._15_.X
flabel locali 16477 14097 16511 14131 0 FreeSans 200 180 0 0 sr_0._15_.A
flabel nwell 16477 13791 16511 13825 0 FreeSans 200 180 0 0 sr_0._15_.VPB
flabel pwell 16477 14335 16511 14369 0 FreeSans 200 180 0 0 sr_0._15_.VNB
rlabel comment 16264 14352 16264 14352 2 sr_0._15_.clkbuf_1
rlabel metal1 16264 14304 16540 14400 5 sr_0._15_.VGND
rlabel metal1 16264 13760 16540 13856 5 sr_0._15_.VPWR
flabel metal1 15102 13795 15138 13825 0 FreeSans 250 0 0 0 sr_0.FILLER_0_3_55.VPWR
flabel metal1 15102 14336 15138 14365 0 FreeSans 250 0 0 0 sr_0.FILLER_0_3_55.VGND
flabel nwell 15109 13801 15129 13818 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_55.VPB
flabel pwell 15108 14341 15132 14363 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_55.VNB
rlabel comment 15160 14352 15160 14352 8 sr_0.FILLER_0_3_55.fill_1
rlabel metal1 15068 14304 15160 14400 5 sr_0.FILLER_0_3_55.VGND
rlabel metal1 15068 13760 15160 13856 5 sr_0.FILLER_0_3_55.VPWR
flabel metal1 14993 13799 15046 13828 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_3_66.VPWR
flabel metal1 14996 14332 15047 14370 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_3_66.VGND
rlabel comment 15068 14352 15068 14352 8 sr_0.TAP_TAPCELL_ROW_3_66.tapvpwrvgnd_1
rlabel metal1 14976 14304 15068 14400 5 sr_0.TAP_TAPCELL_ROW_3_66.VGND
rlabel metal1 14976 13760 15068 13856 5 sr_0.TAP_TAPCELL_ROW_3_66.VPWR
flabel metal1 15190 14335 15224 14369 0 FreeSans 200 0 0 0 sr_0._16_.VGND
flabel metal1 15190 13791 15224 13825 0 FreeSans 200 0 0 0 sr_0._16_.VPWR
flabel locali 15834 14029 15868 14063 0 FreeSans 250 0 0 0 sr_0._16_.S
flabel locali 15742 14029 15776 14063 0 FreeSans 250 0 0 0 sr_0._16_.S
flabel locali 15650 14165 15684 14199 0 FreeSans 250 0 0 0 sr_0._16_.A1
flabel locali 15650 14097 15684 14131 0 FreeSans 250 0 0 0 sr_0._16_.A1
flabel locali 15558 14097 15592 14131 0 FreeSans 250 0 0 0 sr_0._16_.A0
flabel locali 15190 14233 15224 14267 0 FreeSans 250 0 0 0 sr_0._16_.X
flabel locali 15190 13961 15224 13995 0 FreeSans 250 0 0 0 sr_0._16_.X
flabel locali 15190 13893 15224 13927 0 FreeSans 250 0 0 0 sr_0._16_.X
flabel nwell 15234 13791 15268 13825 0 FreeSans 250 0 0 0 sr_0._16_.VPB
flabel pwell 15244 14335 15278 14369 0 FreeSans 250 0 0 0 sr_0._16_.VNB
rlabel comment 15160 14352 15160 14352 2 sr_0._16_.mux2_1
rlabel metal1 15160 14304 15988 14400 5 sr_0._16_.VGND
rlabel metal1 15160 13760 15988 13856 5 sr_0._16_.VPWR
flabel metal1 16201 14335 16235 14369 0 FreeSans 200 180 0 0 sr_0._17_.VGND
flabel metal1 16201 13791 16235 13825 0 FreeSans 200 180 0 0 sr_0._17_.VPWR
flabel locali 16017 14233 16051 14267 0 FreeSans 200 180 0 0 sr_0._17_.X
flabel locali 16017 13961 16051 13995 0 FreeSans 200 180 0 0 sr_0._17_.X
flabel locali 16017 13893 16051 13927 0 FreeSans 200 180 0 0 sr_0._17_.X
flabel locali 16201 14097 16235 14131 0 FreeSans 200 180 0 0 sr_0._17_.A
flabel nwell 16201 13791 16235 13825 0 FreeSans 200 180 0 0 sr_0._17_.VPB
flabel pwell 16201 14335 16235 14369 0 FreeSans 200 180 0 0 sr_0._17_.VNB
rlabel comment 15988 14352 15988 14352 2 sr_0._17_.clkbuf_1
rlabel metal1 15988 14304 16264 14400 5 sr_0._17_.VGND
rlabel metal1 15988 13760 16264 13856 5 sr_0._17_.VPWR
flabel locali 14269 14097 14303 14131 0 FreeSans 200 0 0 0 sr_0.hold2.A
flabel locali 14917 14165 14951 14199 0 FreeSans 200 0 0 0 sr_0.hold2.X
flabel locali 14269 14029 14303 14063 0 FreeSans 200 0 0 0 sr_0.hold2.A
flabel locali 14917 14233 14951 14267 0 FreeSans 200 0 0 0 sr_0.hold2.X
flabel locali 14361 14097 14395 14131 0 FreeSans 200 0 0 0 sr_0.hold2.A
flabel locali 14361 14029 14395 14063 0 FreeSans 200 0 0 0 sr_0.hold2.A
flabel locali 14917 13893 14951 13927 0 FreeSans 200 0 0 0 sr_0.hold2.X
flabel locali 14917 14029 14951 14063 0 FreeSans 200 0 0 0 sr_0.hold2.X
flabel locali 14917 13961 14951 13995 0 FreeSans 200 0 0 0 sr_0.hold2.X
flabel locali 14917 14097 14951 14131 0 FreeSans 200 0 0 0 sr_0.hold2.X
flabel nwell 14269 13791 14303 13825 0 FreeSans 200 0 0 0 sr_0.hold2.VPB
flabel pwell 14269 14335 14303 14369 0 FreeSans 200 0 0 0 sr_0.hold2.VNB
flabel metal1 14269 14335 14303 14369 0 FreeSans 200 0 0 0 sr_0.hold2.VGND
flabel metal1 14269 13791 14303 13825 0 FreeSans 200 0 0 0 sr_0.hold2.VPWR
rlabel comment 14240 14352 14240 14352 2 sr_0.hold2.dlygate4sd3_1
rlabel metal1 14240 14304 14976 14400 5 sr_0.hold2.VGND
rlabel metal1 14240 13760 14976 13856 5 sr_0.hold2.VPWR
flabel metal1 14167 14334 14220 14366 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_65.VGND
flabel metal1 14167 13791 14219 13822 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_65.VPWR
flabel nwell 14178 13799 14212 13817 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_65.VPB
flabel pwell 14177 14340 14209 14362 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_65.VNB
rlabel comment 14240 14352 14240 14352 8 sr_0.FILLER_0_3_65.fill_2
rlabel metal1 14056 14304 14240 14400 5 sr_0.FILLER_0_3_65.VGND
rlabel metal1 14056 13760 14240 13856 5 sr_0.FILLER_0_3_65.VPWR
flabel locali 12429 14029 12463 14063 0 FreeSans 200 0 0 0 sr_0.clkbuf_0_sclk.X
flabel locali 12337 14029 12371 14063 0 FreeSans 200 0 0 0 sr_0.clkbuf_0_sclk.X
flabel locali 12337 14097 12371 14131 0 FreeSans 200 0 0 0 sr_0.clkbuf_0_sclk.X
flabel locali 12429 14097 12463 14131 0 FreeSans 200 0 0 0 sr_0.clkbuf_0_sclk.X
flabel locali 12429 14165 12463 14199 0 FreeSans 200 0 0 0 sr_0.clkbuf_0_sclk.X
flabel locali 12337 14165 12371 14199 0 FreeSans 200 0 0 0 sr_0.clkbuf_0_sclk.X
flabel locali 13993 14165 14027 14199 0 FreeSans 200 0 0 0 sr_0.clkbuf_0_sclk.A
flabel locali 13993 14097 14027 14131 0 FreeSans 200 0 0 0 sr_0.clkbuf_0_sclk.A
flabel pwell 13993 14335 14027 14369 0 FreeSans 200 0 0 0 sr_0.clkbuf_0_sclk.VNB
flabel pwell 14010 14352 14010 14352 0 FreeSans 200 0 0 0 sr_0.clkbuf_0_sclk.VNB
flabel nwell 13993 13791 14027 13825 0 FreeSans 200 0 0 0 sr_0.clkbuf_0_sclk.VPB
flabel nwell 14010 13808 14010 13808 0 FreeSans 200 0 0 0 sr_0.clkbuf_0_sclk.VPB
flabel metal1 13993 14335 14027 14369 0 FreeSans 200 0 0 0 sr_0.clkbuf_0_sclk.VGND
flabel metal1 13993 13791 14027 13825 0 FreeSans 200 0 0 0 sr_0.clkbuf_0_sclk.VPWR
rlabel comment 14056 14352 14056 14352 8 sr_0.clkbuf_0_sclk.clkbuf_16
rlabel metal1 12216 14304 14056 14400 5 sr_0.clkbuf_0_sclk.VGND
rlabel metal1 12216 13760 14056 13856 5 sr_0.clkbuf_0_sclk.VPWR
flabel metal1 12153 14335 12187 14369 0 FreeSans 200 180 0 0 sr_0._27_.VGND
flabel metal1 12153 13791 12187 13825 0 FreeSans 200 180 0 0 sr_0._27_.VPWR
flabel locali 11969 14233 12003 14267 0 FreeSans 200 180 0 0 sr_0._27_.X
flabel locali 11969 13961 12003 13995 0 FreeSans 200 180 0 0 sr_0._27_.X
flabel locali 11969 13893 12003 13927 0 FreeSans 200 180 0 0 sr_0._27_.X
flabel locali 12153 14097 12187 14131 0 FreeSans 200 180 0 0 sr_0._27_.A
flabel nwell 12153 13791 12187 13825 0 FreeSans 200 180 0 0 sr_0._27_.VPB
flabel pwell 12153 14335 12187 14369 0 FreeSans 200 180 0 0 sr_0._27_.VNB
rlabel comment 11940 14352 11940 14352 2 sr_0._27_.clkbuf_1
rlabel metal1 11940 14304 12216 14400 5 sr_0._27_.VGND
rlabel metal1 11940 13760 12216 13856 5 sr_0._27_.VPWR
flabel locali 10130 13893 10164 13927 0 FreeSans 400 0 0 0 sr_0._34_.Q
flabel locali 10130 13961 10164 13995 0 FreeSans 400 0 0 0 sr_0._34_.Q
flabel locali 10130 14029 10164 14063 0 FreeSans 400 0 0 0 sr_0._34_.Q
flabel locali 10130 14233 10164 14267 0 FreeSans 400 0 0 0 sr_0._34_.Q
flabel locali 10425 14165 10459 14199 0 FreeSans 400 0 0 0 sr_0._34_.RESET_B
flabel locali 11601 14029 11635 14063 0 FreeSans 400 0 0 0 sr_0._34_.D
flabel locali 11876 14029 11910 14063 0 FreeSans 400 0 0 0 sr_0._34_.CLK
flabel locali 11876 14097 11910 14131 0 FreeSans 400 0 0 0 sr_0._34_.CLK
flabel locali 10425 14097 10459 14131 0 FreeSans 400 0 0 0 sr_0._34_.RESET_B
flabel metal1 11877 14335 11911 14369 0 FreeSans 200 0 0 0 sr_0._34_.VGND
flabel metal1 11877 13791 11911 13825 0 FreeSans 200 0 0 0 sr_0._34_.VPWR
flabel nwell 11877 13791 11911 13825 0 FreeSans 200 0 0 0 sr_0._34_.VPB
flabel pwell 11877 14335 11911 14369 0 FreeSans 200 0 0 0 sr_0._34_.VNB
rlabel comment 11940 14352 11940 14352 8 sr_0._34_.dfrtp_1
rlabel locali 10411 14145 10459 14225 5 sr_0._34_.RESET_B
rlabel locali 10411 14071 10519 14145 5 sr_0._34_.RESET_B
rlabel metal1 10413 14196 10471 14205 5 sr_0._34_.RESET_B
rlabel metal1 10473 14096 10531 14159 5 sr_0._34_.RESET_B
rlabel metal1 10413 14159 10531 14168 5 sr_0._34_.RESET_B
rlabel metal1 11061 14159 11191 14168 5 sr_0._34_.RESET_B
rlabel metal1 10413 14168 11191 14196 5 sr_0._34_.RESET_B
rlabel metal1 11061 14196 11191 14205 5 sr_0._34_.RESET_B
rlabel metal1 10100 14304 11940 14400 5 sr_0._34_.VGND
rlabel metal1 10100 13760 11940 13856 5 sr_0._34_.VPWR
flabel metal1 10027 14334 10080 14366 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_110.VGND
flabel metal1 10027 13791 10079 13822 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_110.VPWR
flabel nwell 10038 13799 10072 13817 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_110.VPB
flabel pwell 10037 14340 10069 14362 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_110.VNB
rlabel comment 10100 14352 10100 14352 8 sr_0.FILLER_0_3_110.fill_2
rlabel metal1 9916 14304 10100 14400 5 sr_0.FILLER_0_3_110.VGND
rlabel metal1 9916 13760 10100 13856 5 sr_0.FILLER_0_3_110.VPWR
flabel metal1 9761 14335 9795 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_113.VGND
flabel metal1 9761 13791 9795 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_113.VPWR
flabel nwell 9761 13791 9795 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_113.VPB
flabel pwell 9761 14335 9795 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_113.VNB
rlabel comment 9824 14352 9824 14352 8 sr_0.FILLER_0_3_113.decap_12
flabel metal1 8657 14335 8691 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_125.VGND
flabel metal1 8657 13791 8691 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_125.VPWR
flabel nwell 8657 13791 8691 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_125.VPB
flabel pwell 8657 14335 8691 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_125.VNB
rlabel comment 8720 14352 8720 14352 8 sr_0.FILLER_0_3_125.decap_12
flabel metal1 9841 13799 9894 13828 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_3_67.VPWR
flabel metal1 9844 14332 9895 14370 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_3_67.VGND
rlabel comment 9916 14352 9916 14352 8 sr_0.TAP_TAPCELL_ROW_3_67.tapvpwrvgnd_1
rlabel metal1 9824 14304 9916 14400 5 sr_0.TAP_TAPCELL_ROW_3_67.VGND
rlabel metal1 9824 13760 9916 13856 5 sr_0.TAP_TAPCELL_ROW_3_67.VPWR
flabel metal1 7553 14335 7587 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_137.VGND
flabel metal1 7553 13791 7587 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_137.VPWR
flabel nwell 7553 13791 7587 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_137.VPB
flabel pwell 7553 14335 7587 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_137.VNB
rlabel comment 7616 14352 7616 14352 8 sr_0.FILLER_0_3_137.decap_12
flabel metal1 6449 14335 6483 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_149.VGND
flabel metal1 6449 13791 6483 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_149.VPWR
flabel nwell 6449 13791 6483 13825 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_149.VPB
flabel pwell 6449 14335 6483 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_149.VNB
rlabel comment 6512 14352 6512 14352 8 sr_0.FILLER_0_3_149.decap_12
flabel metal1 5335 14334 5388 14366 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_161.VGND
flabel metal1 5335 13791 5387 13822 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_161.VPWR
flabel nwell 5346 13799 5380 13817 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_161.VPB
flabel pwell 5345 14340 5377 14362 0 FreeSans 200 0 0 0 sr_0.FILLER_0_3_161.VNB
rlabel comment 5408 14352 5408 14352 8 sr_0.FILLER_0_3_161.fill_2
rlabel metal1 5224 14304 5408 14400 5 sr_0.FILLER_0_3_161.VGND
rlabel metal1 5224 13760 5408 13856 5 sr_0.FILLER_0_3_161.VPWR
flabel metal1 4977 13791 5011 13825 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_3_Right_3.VPWR
flabel metal1 4977 14335 5011 14369 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_3_Right_3.VGND
flabel nwell 4977 13791 5011 13825 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_3_Right_3.VPB
flabel pwell 4977 14335 5011 14369 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_3_Right_3.VNB
rlabel comment 4948 14352 4948 14352 2 sr_0.PHY_EDGE_ROW_3_Right_3.decap_3
rlabel metal1 4948 14304 5224 14400 5 sr_0.PHY_EDGE_ROW_3_Right_3.VGND
rlabel metal1 4948 13760 5224 13856 5 sr_0.PHY_EDGE_ROW_3_Right_3.VPWR
flabel metal1 19881 14335 19915 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_3.VGND
flabel metal1 19881 14879 19915 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_3.VPWR
flabel nwell 19881 14879 19915 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_3.VPB
flabel pwell 19881 14335 19915 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_3.VNB
rlabel comment 19944 14352 19944 14352 6 sr_0.FILLER_0_4_3.decap_12
flabel metal1 18777 14335 18811 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_15.VGND
flabel metal1 18777 14879 18811 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_15.VPWR
flabel nwell 18777 14879 18811 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_15.VPB
flabel pwell 18777 14335 18811 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_15.VNB
rlabel comment 18840 14352 18840 14352 6 sr_0.FILLER_0_4_15.decap_12
flabel metal1 20157 14879 20191 14913 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_4_Left_32.VPWR
flabel metal1 20157 14335 20191 14369 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_4_Left_32.VGND
flabel nwell 20157 14879 20191 14913 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_4_Left_32.VPB
flabel pwell 20157 14335 20191 14369 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_4_Left_32.VNB
rlabel comment 20220 14352 20220 14352 6 sr_0.PHY_EDGE_ROW_4_Left_32.decap_3
rlabel metal1 19944 14304 20220 14400 1 sr_0.PHY_EDGE_ROW_4_Left_32.VGND
rlabel metal1 19944 14848 20220 14944 1 sr_0.PHY_EDGE_ROW_4_Left_32.VPWR
flabel metal1 17678 14879 17714 14909 0 FreeSans 250 0 0 0 sr_0.FILLER_0_4_27.VPWR
flabel metal1 17678 14339 17714 14368 0 FreeSans 250 0 0 0 sr_0.FILLER_0_4_27.VGND
flabel nwell 17685 14886 17705 14903 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_27.VPB
flabel pwell 17684 14341 17708 14363 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_27.VNB
rlabel comment 17736 14352 17736 14352 6 sr_0.FILLER_0_4_27.fill_1
rlabel metal1 17644 14304 17736 14400 1 sr_0.FILLER_0_4_27.VGND
rlabel metal1 17644 14848 17736 14944 1 sr_0.FILLER_0_4_27.VPWR
flabel metal1 17489 14335 17523 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_29.VGND
flabel metal1 17489 14879 17523 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_29.VPWR
flabel nwell 17489 14879 17523 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_29.VPB
flabel pwell 17489 14335 17523 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_29.VNB
rlabel comment 17552 14352 17552 14352 6 sr_0.FILLER_0_4_29.decap_12
flabel metal1 16390 14879 16426 14909 0 FreeSans 250 0 0 0 sr_0.FILLER_0_4_41.VPWR
flabel metal1 16390 14339 16426 14368 0 FreeSans 250 0 0 0 sr_0.FILLER_0_4_41.VGND
flabel nwell 16397 14886 16417 14903 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_41.VPB
flabel pwell 16396 14341 16420 14363 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_41.VNB
rlabel comment 16448 14352 16448 14352 6 sr_0.FILLER_0_4_41.fill_1
rlabel metal1 16356 14304 16448 14400 1 sr_0.FILLER_0_4_41.VGND
rlabel metal1 16356 14848 16448 14944 1 sr_0.FILLER_0_4_41.VPWR
flabel metal1 17569 14876 17622 14905 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_4_68.VPWR
flabel metal1 17572 14334 17623 14372 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_4_68.VGND
rlabel comment 17644 14352 17644 14352 6 sr_0.TAP_TAPCELL_ROW_4_68.tapvpwrvgnd_1
rlabel metal1 17552 14304 17644 14400 1 sr_0.TAP_TAPCELL_ROW_4_68.VGND
rlabel metal1 17552 14848 17644 14944 1 sr_0.TAP_TAPCELL_ROW_4_68.VPWR
flabel metal1 14269 14335 14303 14369 0 FreeSans 200 180 0 0 sr_0._19_.VGND
flabel metal1 14269 14879 14303 14913 0 FreeSans 200 180 0 0 sr_0._19_.VPWR
flabel locali 14453 14437 14487 14471 0 FreeSans 200 180 0 0 sr_0._19_.X
flabel locali 14453 14709 14487 14743 0 FreeSans 200 180 0 0 sr_0._19_.X
flabel locali 14453 14777 14487 14811 0 FreeSans 200 180 0 0 sr_0._19_.X
flabel locali 14269 14573 14303 14607 0 FreeSans 200 180 0 0 sr_0._19_.A
flabel nwell 14269 14879 14303 14913 0 FreeSans 200 180 0 0 sr_0._19_.VPB
flabel pwell 14269 14335 14303 14369 0 FreeSans 200 180 0 0 sr_0._19_.VNB
rlabel comment 14516 14352 14516 14352 6 sr_0._19_.clkbuf_1
rlabel metal1 14240 14304 14516 14400 1 sr_0._19_.VGND
rlabel metal1 14240 14848 14516 14944 1 sr_0._19_.VPWR
flabel locali 14546 14777 14580 14811 0 FreeSans 400 0 0 0 sr_0._29_.Q
flabel locali 14546 14709 14580 14743 0 FreeSans 400 0 0 0 sr_0._29_.Q
flabel locali 14546 14641 14580 14675 0 FreeSans 400 0 0 0 sr_0._29_.Q
flabel locali 14546 14437 14580 14471 0 FreeSans 400 0 0 0 sr_0._29_.Q
flabel locali 14841 14505 14875 14539 0 FreeSans 400 0 0 0 sr_0._29_.RESET_B
flabel locali 16017 14641 16051 14675 0 FreeSans 400 0 0 0 sr_0._29_.D
flabel locali 16292 14641 16326 14675 0 FreeSans 400 0 0 0 sr_0._29_.CLK
flabel locali 16292 14573 16326 14607 0 FreeSans 400 0 0 0 sr_0._29_.CLK
flabel locali 14841 14573 14875 14607 0 FreeSans 400 0 0 0 sr_0._29_.RESET_B
flabel metal1 16293 14335 16327 14369 0 FreeSans 200 0 0 0 sr_0._29_.VGND
flabel metal1 16293 14879 16327 14913 0 FreeSans 200 0 0 0 sr_0._29_.VPWR
flabel nwell 16293 14879 16327 14913 0 FreeSans 200 0 0 0 sr_0._29_.VPB
flabel pwell 16293 14335 16327 14369 0 FreeSans 200 0 0 0 sr_0._29_.VNB
rlabel comment 16356 14352 16356 14352 6 sr_0._29_.dfrtp_1
rlabel locali 14827 14479 14875 14559 1 sr_0._29_.RESET_B
rlabel locali 14827 14559 14935 14633 1 sr_0._29_.RESET_B
rlabel metal1 14829 14499 14887 14508 1 sr_0._29_.RESET_B
rlabel metal1 14889 14545 14947 14608 1 sr_0._29_.RESET_B
rlabel metal1 14829 14536 14947 14545 1 sr_0._29_.RESET_B
rlabel metal1 15477 14536 15607 14545 1 sr_0._29_.RESET_B
rlabel metal1 14829 14508 15607 14536 1 sr_0._29_.RESET_B
rlabel metal1 15477 14499 15607 14508 1 sr_0._29_.RESET_B
rlabel metal1 14516 14304 16356 14400 1 sr_0._29_.VGND
rlabel metal1 14516 14848 16356 14944 1 sr_0._29_.VPWR
flabel metal1 14177 14879 14211 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_65.VPWR
flabel metal1 14177 14335 14211 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_65.VGND
flabel nwell 14177 14879 14211 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_65.VPB
flabel pwell 14177 14335 14211 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_65.VNB
rlabel comment 14240 14352 14240 14352 6 sr_0.FILLER_0_4_65.decap_8
rlabel metal1 13504 14304 14240 14400 1 sr_0.FILLER_0_4_65.VGND
rlabel metal1 13504 14848 14240 14944 1 sr_0.FILLER_0_4_65.VPWR
flabel metal1 12603 14338 12656 14370 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_82.VGND
flabel metal1 12603 14882 12655 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_82.VPWR
flabel nwell 12614 14887 12648 14905 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_82.VPB
flabel pwell 12613 14342 12645 14364 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_82.VNB
rlabel comment 12676 14352 12676 14352 6 sr_0.FILLER_0_4_82.fill_2
rlabel metal1 12492 14304 12676 14400 1 sr_0.FILLER_0_4_82.VGND
rlabel metal1 12492 14848 12676 14944 1 sr_0.FILLER_0_4_82.VPWR
flabel metal1 13440 14335 13474 14369 0 FreeSans 200 0 0 0 sr_0._20_.VGND
flabel metal1 13440 14879 13474 14913 0 FreeSans 200 0 0 0 sr_0._20_.VPWR
flabel locali 12796 14641 12830 14675 0 FreeSans 250 0 0 0 sr_0._20_.S
flabel locali 12888 14641 12922 14675 0 FreeSans 250 0 0 0 sr_0._20_.S
flabel locali 12980 14505 13014 14539 0 FreeSans 250 0 0 0 sr_0._20_.A1
flabel locali 12980 14573 13014 14607 0 FreeSans 250 0 0 0 sr_0._20_.A1
flabel locali 13072 14573 13106 14607 0 FreeSans 250 0 0 0 sr_0._20_.A0
flabel locali 13440 14437 13474 14471 0 FreeSans 250 0 0 0 sr_0._20_.X
flabel locali 13440 14709 13474 14743 0 FreeSans 250 0 0 0 sr_0._20_.X
flabel locali 13440 14777 13474 14811 0 FreeSans 250 0 0 0 sr_0._20_.X
flabel nwell 13396 14879 13430 14913 0 FreeSans 250 0 0 0 sr_0._20_.VPB
flabel pwell 13386 14335 13420 14369 0 FreeSans 250 0 0 0 sr_0._20_.VNB
rlabel comment 13504 14352 13504 14352 6 sr_0._20_.mux2_1
rlabel metal1 12676 14304 13504 14400 1 sr_0._20_.VGND
rlabel metal1 12676 14848 13504 14944 1 sr_0._20_.VPWR
flabel metal1 12337 14879 12371 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_85.VPWR
flabel metal1 12337 14335 12371 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_85.VGND
flabel nwell 12337 14879 12371 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_85.VPB
flabel pwell 12337 14335 12371 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_85.VNB
rlabel comment 12400 14352 12400 14352 6 sr_0.FILLER_0_4_85.decap_8
rlabel metal1 11664 14304 12400 14400 1 sr_0.FILLER_0_4_85.VGND
rlabel metal1 11664 14848 12400 14944 1 sr_0.FILLER_0_4_85.VPWR
flabel metal1 11591 14338 11644 14370 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_93.VGND
flabel metal1 11591 14882 11643 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_93.VPWR
flabel nwell 11602 14887 11636 14905 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_93.VPB
flabel pwell 11601 14342 11633 14364 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_93.VNB
rlabel comment 11664 14352 11664 14352 6 sr_0.FILLER_0_4_93.fill_2
rlabel metal1 11480 14304 11664 14400 1 sr_0.FILLER_0_4_93.VGND
rlabel metal1 11480 14848 11664 14944 1 sr_0.FILLER_0_4_93.VPWR
flabel metal1 10589 14335 10623 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_104.VGND
flabel metal1 10589 14879 10623 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_104.VPWR
flabel nwell 10589 14879 10623 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_104.VPB
flabel pwell 10589 14335 10623 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_104.VNB
rlabel comment 10652 14352 10652 14352 6 sr_0.FILLER_0_4_104.decap_12
flabel metal1 12417 14876 12470 14905 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_4_69.VPWR
flabel metal1 12420 14334 12471 14372 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_4_69.VGND
rlabel comment 12492 14352 12492 14352 6 sr_0.TAP_TAPCELL_ROW_4_69.tapvpwrvgnd_1
rlabel metal1 12400 14304 12492 14400 1 sr_0.TAP_TAPCELL_ROW_4_69.VGND
rlabel metal1 12400 14848 12492 14944 1 sr_0.TAP_TAPCELL_ROW_4_69.VPWR
flabel metal1 11416 14335 11450 14369 0 FreeSans 200 0 0 0 sr_0._26_.VGND
flabel metal1 11416 14879 11450 14913 0 FreeSans 200 0 0 0 sr_0._26_.VPWR
flabel locali 10772 14641 10806 14675 0 FreeSans 250 0 0 0 sr_0._26_.S
flabel locali 10864 14641 10898 14675 0 FreeSans 250 0 0 0 sr_0._26_.S
flabel locali 10956 14505 10990 14539 0 FreeSans 250 0 0 0 sr_0._26_.A1
flabel locali 10956 14573 10990 14607 0 FreeSans 250 0 0 0 sr_0._26_.A1
flabel locali 11048 14573 11082 14607 0 FreeSans 250 0 0 0 sr_0._26_.A0
flabel locali 11416 14437 11450 14471 0 FreeSans 250 0 0 0 sr_0._26_.X
flabel locali 11416 14709 11450 14743 0 FreeSans 250 0 0 0 sr_0._26_.X
flabel locali 11416 14777 11450 14811 0 FreeSans 250 0 0 0 sr_0._26_.X
flabel nwell 11372 14879 11406 14913 0 FreeSans 250 0 0 0 sr_0._26_.VPB
flabel pwell 11362 14335 11396 14369 0 FreeSans 250 0 0 0 sr_0._26_.VNB
rlabel comment 11480 14352 11480 14352 6 sr_0._26_.mux2_1
rlabel metal1 10652 14304 11480 14400 1 sr_0._26_.VGND
rlabel metal1 10652 14848 11480 14944 1 sr_0._26_.VPWR
flabel metal1 9485 14335 9519 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_116.VGND
flabel metal1 9485 14879 9519 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_116.VPWR
flabel nwell 9485 14879 9519 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_116.VPB
flabel pwell 9485 14335 9519 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_116.VNB
rlabel comment 9548 14352 9548 14352 6 sr_0.FILLER_0_4_116.decap_12
flabel metal1 8381 14335 8415 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_128.VGND
flabel metal1 8381 14879 8415 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_128.VPWR
flabel nwell 8381 14879 8415 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_128.VPB
flabel pwell 8381 14335 8415 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_128.VNB
rlabel comment 8444 14352 8444 14352 6 sr_0.FILLER_0_4_128.decap_12
flabel metal1 7185 14335 7219 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_141.VGND
flabel metal1 7185 14879 7219 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_141.VPWR
flabel nwell 7185 14879 7219 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_141.VPB
flabel pwell 7185 14335 7219 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_141.VNB
rlabel comment 7248 14352 7248 14352 6 sr_0.FILLER_0_4_141.decap_12
flabel metal1 7265 14876 7318 14905 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_4_70.VPWR
flabel metal1 7268 14334 7319 14372 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_4_70.VGND
rlabel comment 7340 14352 7340 14352 6 sr_0.TAP_TAPCELL_ROW_4_70.tapvpwrvgnd_1
rlabel metal1 7248 14304 7340 14400 1 sr_0.TAP_TAPCELL_ROW_4_70.VGND
rlabel metal1 7248 14848 7340 14944 1 sr_0.TAP_TAPCELL_ROW_4_70.VPWR
flabel metal1 6081 14879 6115 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_153.VPWR
flabel metal1 6081 14335 6115 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_153.VGND
flabel nwell 6081 14879 6115 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_153.VPB
flabel pwell 6081 14335 6115 14369 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_153.VNB
rlabel comment 6144 14352 6144 14352 6 sr_0.FILLER_0_4_153.decap_8
rlabel metal1 5408 14304 6144 14400 1 sr_0.FILLER_0_4_153.VGND
rlabel metal1 5408 14848 6144 14944 1 sr_0.FILLER_0_4_153.VPWR
flabel metal1 5335 14338 5388 14370 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_161.VGND
flabel metal1 5335 14882 5387 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_161.VPWR
flabel nwell 5346 14887 5380 14905 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_161.VPB
flabel pwell 5345 14342 5377 14364 0 FreeSans 200 0 0 0 sr_0.FILLER_0_4_161.VNB
rlabel comment 5408 14352 5408 14352 6 sr_0.FILLER_0_4_161.fill_2
rlabel metal1 5224 14304 5408 14400 1 sr_0.FILLER_0_4_161.VGND
rlabel metal1 5224 14848 5408 14944 1 sr_0.FILLER_0_4_161.VPWR
flabel metal1 4977 14879 5011 14913 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_4_Right_4.VPWR
flabel metal1 4977 14335 5011 14369 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_4_Right_4.VGND
flabel nwell 4977 14879 5011 14913 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_4_Right_4.VPB
flabel pwell 4977 14335 5011 14369 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_4_Right_4.VNB
rlabel comment 4948 14352 4948 14352 4 sr_0.PHY_EDGE_ROW_4_Right_4.decap_3
rlabel metal1 4948 14304 5224 14400 1 sr_0.PHY_EDGE_ROW_4_Right_4.VGND
rlabel metal1 4948 14848 5224 14944 1 sr_0.PHY_EDGE_ROW_4_Right_4.VPWR
flabel metal1 19881 15423 19915 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_3.VGND
flabel metal1 19881 14879 19915 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_3.VPWR
flabel nwell 19881 14879 19915 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_3.VPB
flabel pwell 19881 15423 19915 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_3.VNB
rlabel comment 19944 15440 19944 15440 8 sr_0.FILLER_0_5_3.decap_12
flabel metal1 18777 15423 18811 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_15.VGND
flabel metal1 18777 14879 18811 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_15.VPWR
flabel nwell 18777 14879 18811 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_15.VPB
flabel pwell 18777 15423 18811 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_15.VNB
rlabel comment 18840 15440 18840 15440 8 sr_0.FILLER_0_5_15.decap_12
flabel metal1 20157 14879 20191 14913 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_5_Left_33.VPWR
flabel metal1 20157 15423 20191 15457 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_5_Left_33.VGND
flabel nwell 20157 14879 20191 14913 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_5_Left_33.VPB
flabel pwell 20157 15423 20191 15457 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_5_Left_33.VNB
rlabel comment 20220 15440 20220 15440 8 sr_0.PHY_EDGE_ROW_5_Left_33.decap_3
rlabel metal1 19944 15392 20220 15488 5 sr_0.PHY_EDGE_ROW_5_Left_33.VGND
rlabel metal1 19944 14848 20220 14944 5 sr_0.PHY_EDGE_ROW_5_Left_33.VPWR
flabel metal1 17673 15423 17707 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_27.VGND
flabel metal1 17673 14879 17707 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_27.VPWR
flabel nwell 17673 14879 17707 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_27.VPB
flabel pwell 17673 15423 17707 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_27.VNB
rlabel comment 17736 15440 17736 15440 8 sr_0.FILLER_0_5_27.decap_12
flabel metal1 16569 14879 16603 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_39.VPWR
flabel metal1 16569 15423 16603 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_39.VGND
flabel nwell 16569 14879 16603 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_39.VPB
flabel pwell 16569 15423 16603 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_39.VNB
rlabel comment 16632 15440 16632 15440 8 sr_0.FILLER_0_5_39.decap_6
rlabel metal1 16080 15392 16632 15488 5 sr_0.FILLER_0_5_39.VGND
rlabel metal1 16080 14848 16632 14944 5 sr_0.FILLER_0_5_39.VPWR
flabel metal1 15281 14879 15315 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_53.VPWR
flabel metal1 15281 15423 15315 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_53.VGND
flabel nwell 15281 14879 15315 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_53.VPB
flabel pwell 15281 15423 15315 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_53.VNB
rlabel comment 15344 15440 15344 15440 8 sr_0.FILLER_0_5_53.decap_3
rlabel metal1 15068 15392 15344 15488 5 sr_0.FILLER_0_5_53.VGND
rlabel metal1 15068 14848 15344 14944 5 sr_0.FILLER_0_5_53.VPWR
flabel metal1 14913 15423 14947 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_57.VGND
flabel metal1 14913 14879 14947 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_57.VPWR
flabel nwell 14913 14879 14947 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_57.VPB
flabel pwell 14913 15423 14947 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_57.VNB
rlabel comment 14976 15440 14976 15440 8 sr_0.FILLER_0_5_57.decap_12
flabel metal1 14993 14887 15046 14916 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_5_71.VPWR
flabel metal1 14996 15420 15047 15458 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_5_71.VGND
rlabel comment 15068 15440 15068 15440 8 sr_0.TAP_TAPCELL_ROW_5_71.tapvpwrvgnd_1
rlabel metal1 14976 15392 15068 15488 5 sr_0.TAP_TAPCELL_ROW_5_71.VGND
rlabel metal1 14976 14848 15068 14944 5 sr_0.TAP_TAPCELL_ROW_5_71.VPWR
flabel locali 15373 15185 15407 15219 0 FreeSans 200 0 0 0 sr_0.hold3.A
flabel locali 16021 15253 16055 15287 0 FreeSans 200 0 0 0 sr_0.hold3.X
flabel locali 15373 15117 15407 15151 0 FreeSans 200 0 0 0 sr_0.hold3.A
flabel locali 16021 15321 16055 15355 0 FreeSans 200 0 0 0 sr_0.hold3.X
flabel locali 15465 15185 15499 15219 0 FreeSans 200 0 0 0 sr_0.hold3.A
flabel locali 15465 15117 15499 15151 0 FreeSans 200 0 0 0 sr_0.hold3.A
flabel locali 16021 14981 16055 15015 0 FreeSans 200 0 0 0 sr_0.hold3.X
flabel locali 16021 15117 16055 15151 0 FreeSans 200 0 0 0 sr_0.hold3.X
flabel locali 16021 15049 16055 15083 0 FreeSans 200 0 0 0 sr_0.hold3.X
flabel locali 16021 15185 16055 15219 0 FreeSans 200 0 0 0 sr_0.hold3.X
flabel nwell 15373 14879 15407 14913 0 FreeSans 200 0 0 0 sr_0.hold3.VPB
flabel pwell 15373 15423 15407 15457 0 FreeSans 200 0 0 0 sr_0.hold3.VNB
flabel metal1 15373 15423 15407 15457 0 FreeSans 200 0 0 0 sr_0.hold3.VGND
flabel metal1 15373 14879 15407 14913 0 FreeSans 200 0 0 0 sr_0.hold3.VPWR
rlabel comment 15344 15440 15344 15440 2 sr_0.hold3.dlygate4sd3_1
rlabel metal1 15344 15392 16080 15488 5 sr_0.hold3.VGND
rlabel metal1 15344 14848 16080 14944 5 sr_0.hold3.VPWR
flabel metal1 13809 15423 13843 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_69.VGND
flabel metal1 13809 14879 13843 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_69.VPWR
flabel nwell 13809 14879 13843 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_69.VPB
flabel pwell 13809 15423 13843 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_69.VNB
rlabel comment 13872 15440 13872 15440 8 sr_0.FILLER_0_5_69.decap_4
rlabel metal1 13504 15392 13872 15488 5 sr_0.FILLER_0_5_69.VGND
rlabel metal1 13504 14848 13872 14944 5 sr_0.FILLER_0_5_69.VPWR
flabel metal1 12705 15423 12739 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_81.VGND
flabel metal1 12705 14879 12739 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_81.VPWR
flabel nwell 12705 14879 12739 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_81.VPB
flabel pwell 12705 15423 12739 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_81.VNB
rlabel comment 12768 15440 12768 15440 8 sr_0.FILLER_0_5_81.decap_12
flabel locali 12797 15185 12831 15219 0 FreeSans 200 0 0 0 sr_0.hold4.A
flabel locali 13445 15253 13479 15287 0 FreeSans 200 0 0 0 sr_0.hold4.X
flabel locali 12797 15117 12831 15151 0 FreeSans 200 0 0 0 sr_0.hold4.A
flabel locali 13445 15321 13479 15355 0 FreeSans 200 0 0 0 sr_0.hold4.X
flabel locali 12889 15185 12923 15219 0 FreeSans 200 0 0 0 sr_0.hold4.A
flabel locali 12889 15117 12923 15151 0 FreeSans 200 0 0 0 sr_0.hold4.A
flabel locali 13445 14981 13479 15015 0 FreeSans 200 0 0 0 sr_0.hold4.X
flabel locali 13445 15117 13479 15151 0 FreeSans 200 0 0 0 sr_0.hold4.X
flabel locali 13445 15049 13479 15083 0 FreeSans 200 0 0 0 sr_0.hold4.X
flabel locali 13445 15185 13479 15219 0 FreeSans 200 0 0 0 sr_0.hold4.X
flabel nwell 12797 14879 12831 14913 0 FreeSans 200 0 0 0 sr_0.hold4.VPB
flabel pwell 12797 15423 12831 15457 0 FreeSans 200 0 0 0 sr_0.hold4.VNB
flabel metal1 12797 15423 12831 15457 0 FreeSans 200 0 0 0 sr_0.hold4.VGND
flabel metal1 12797 14879 12831 14913 0 FreeSans 200 0 0 0 sr_0.hold4.VPWR
rlabel comment 12768 15440 12768 15440 2 sr_0.hold4.dlygate4sd3_1
rlabel metal1 12768 15392 13504 15488 5 sr_0.hold4.VGND
rlabel metal1 12768 14848 13504 14944 5 sr_0.hold4.VPWR
flabel metal1 11601 15423 11635 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_93.VGND
flabel metal1 11601 14879 11635 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_93.VPWR
flabel nwell 11601 14879 11635 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_93.VPB
flabel pwell 11601 15423 11635 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_93.VNB
rlabel comment 11664 15440 11664 15440 8 sr_0.FILLER_0_5_93.decap_12
flabel metal1 10497 14879 10531 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_105.VPWR
flabel metal1 10497 15423 10531 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_105.VGND
flabel nwell 10497 14879 10531 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_105.VPB
flabel pwell 10497 15423 10531 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_105.VNB
rlabel comment 10560 15440 10560 15440 8 sr_0.FILLER_0_5_105.decap_6
rlabel metal1 10008 15392 10560 15488 5 sr_0.FILLER_0_5_105.VGND
rlabel metal1 10008 14848 10560 14944 5 sr_0.FILLER_0_5_105.VPWR
flabel metal1 9950 14883 9986 14913 0 FreeSans 250 0 0 0 sr_0.FILLER_0_5_111.VPWR
flabel metal1 9950 15424 9986 15453 0 FreeSans 250 0 0 0 sr_0.FILLER_0_5_111.VGND
flabel nwell 9957 14889 9977 14906 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_111.VPB
flabel pwell 9956 15429 9980 15451 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_111.VNB
rlabel comment 10008 15440 10008 15440 8 sr_0.FILLER_0_5_111.fill_1
rlabel metal1 9916 15392 10008 15488 5 sr_0.FILLER_0_5_111.VGND
rlabel metal1 9916 14848 10008 14944 5 sr_0.FILLER_0_5_111.VPWR
flabel metal1 9761 15423 9795 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_113.VGND
flabel metal1 9761 14879 9795 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_113.VPWR
flabel nwell 9761 14879 9795 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_113.VPB
flabel pwell 9761 15423 9795 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_113.VNB
rlabel comment 9824 15440 9824 15440 8 sr_0.FILLER_0_5_113.decap_12
flabel metal1 8657 15423 8691 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_125.VGND
flabel metal1 8657 14879 8691 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_125.VPWR
flabel nwell 8657 14879 8691 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_125.VPB
flabel pwell 8657 15423 8691 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_125.VNB
rlabel comment 8720 15440 8720 15440 8 sr_0.FILLER_0_5_125.decap_12
flabel metal1 9841 14887 9894 14916 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_5_72.VPWR
flabel metal1 9844 15420 9895 15458 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_5_72.VGND
rlabel comment 9916 15440 9916 15440 8 sr_0.TAP_TAPCELL_ROW_5_72.tapvpwrvgnd_1
rlabel metal1 9824 15392 9916 15488 5 sr_0.TAP_TAPCELL_ROW_5_72.VGND
rlabel metal1 9824 14848 9916 14944 5 sr_0.TAP_TAPCELL_ROW_5_72.VPWR
flabel metal1 7553 15423 7587 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_137.VGND
flabel metal1 7553 14879 7587 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_137.VPWR
flabel nwell 7553 14879 7587 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_137.VPB
flabel pwell 7553 15423 7587 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_137.VNB
rlabel comment 7616 15440 7616 15440 8 sr_0.FILLER_0_5_137.decap_12
flabel metal1 6449 15423 6483 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_149.VGND
flabel metal1 6449 14879 6483 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_149.VPWR
flabel nwell 6449 14879 6483 14913 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_149.VPB
flabel pwell 6449 15423 6483 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_149.VNB
rlabel comment 6512 15440 6512 15440 8 sr_0.FILLER_0_5_149.decap_12
flabel metal1 5335 15422 5388 15454 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_161.VGND
flabel metal1 5335 14879 5387 14910 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_161.VPWR
flabel nwell 5346 14887 5380 14905 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_161.VPB
flabel pwell 5345 15428 5377 15450 0 FreeSans 200 0 0 0 sr_0.FILLER_0_5_161.VNB
rlabel comment 5408 15440 5408 15440 8 sr_0.FILLER_0_5_161.fill_2
rlabel metal1 5224 15392 5408 15488 5 sr_0.FILLER_0_5_161.VGND
rlabel metal1 5224 14848 5408 14944 5 sr_0.FILLER_0_5_161.VPWR
flabel metal1 4977 14879 5011 14913 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_5_Right_5.VPWR
flabel metal1 4977 15423 5011 15457 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_5_Right_5.VGND
flabel nwell 4977 14879 5011 14913 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_5_Right_5.VPB
flabel pwell 4977 15423 5011 15457 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_5_Right_5.VNB
rlabel comment 4948 15440 4948 15440 2 sr_0.PHY_EDGE_ROW_5_Right_5.decap_3
rlabel metal1 4948 15392 5224 15488 5 sr_0.PHY_EDGE_ROW_5_Right_5.VGND
rlabel metal1 4948 14848 5224 14944 5 sr_0.PHY_EDGE_ROW_5_Right_5.VPWR
flabel metal1 19881 15423 19915 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_3.VGND
flabel metal1 19881 15967 19915 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_3.VPWR
flabel nwell 19881 15967 19915 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_3.VPB
flabel pwell 19881 15423 19915 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_3.VNB
rlabel comment 19944 15440 19944 15440 6 sr_0.FILLER_0_6_3.decap_12
flabel metal1 18777 15423 18811 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_15.VGND
flabel metal1 18777 15967 18811 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_15.VPWR
flabel nwell 18777 15967 18811 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_15.VPB
flabel pwell 18777 15423 18811 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_15.VNB
rlabel comment 18840 15440 18840 15440 6 sr_0.FILLER_0_6_15.decap_12
flabel metal1 19881 16511 19915 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_3.VGND
flabel metal1 19881 15967 19915 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_3.VPWR
flabel nwell 19881 15967 19915 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_3.VPB
flabel pwell 19881 16511 19915 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_3.VNB
rlabel comment 19944 16528 19944 16528 8 sr_0.FILLER_0_7_3.decap_12
flabel metal1 18777 16511 18811 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_15.VGND
flabel metal1 18777 15967 18811 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_15.VPWR
flabel nwell 18777 15967 18811 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_15.VPB
flabel pwell 18777 16511 18811 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_15.VNB
rlabel comment 18840 16528 18840 16528 8 sr_0.FILLER_0_7_15.decap_12
flabel metal1 20157 15967 20191 16001 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_6_Left_34.VPWR
flabel metal1 20157 15423 20191 15457 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_6_Left_34.VGND
flabel nwell 20157 15967 20191 16001 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_6_Left_34.VPB
flabel pwell 20157 15423 20191 15457 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_6_Left_34.VNB
rlabel comment 20220 15440 20220 15440 6 sr_0.PHY_EDGE_ROW_6_Left_34.decap_3
rlabel metal1 19944 15392 20220 15488 1 sr_0.PHY_EDGE_ROW_6_Left_34.VGND
rlabel metal1 19944 15936 20220 16032 1 sr_0.PHY_EDGE_ROW_6_Left_34.VPWR
flabel metal1 20157 15967 20191 16001 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_7_Left_35.VPWR
flabel metal1 20157 16511 20191 16545 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_7_Left_35.VGND
flabel nwell 20157 15967 20191 16001 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_7_Left_35.VPB
flabel pwell 20157 16511 20191 16545 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_7_Left_35.VNB
rlabel comment 20220 16528 20220 16528 8 sr_0.PHY_EDGE_ROW_7_Left_35.decap_3
rlabel metal1 19944 16480 20220 16576 5 sr_0.PHY_EDGE_ROW_7_Left_35.VGND
rlabel metal1 19944 15936 20220 16032 5 sr_0.PHY_EDGE_ROW_7_Left_35.VPWR
flabel metal1 17678 15967 17714 15997 0 FreeSans 250 0 0 0 sr_0.FILLER_0_6_27.VPWR
flabel metal1 17678 15427 17714 15456 0 FreeSans 250 0 0 0 sr_0.FILLER_0_6_27.VGND
flabel nwell 17685 15974 17705 15991 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_27.VPB
flabel pwell 17684 15429 17708 15451 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_27.VNB
rlabel comment 17736 15440 17736 15440 6 sr_0.FILLER_0_6_27.fill_1
rlabel metal1 17644 15392 17736 15488 1 sr_0.FILLER_0_6_27.VGND
rlabel metal1 17644 15936 17736 16032 1 sr_0.FILLER_0_6_27.VPWR
flabel metal1 17489 15423 17523 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_29.VGND
flabel metal1 17489 15967 17523 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_29.VPWR
flabel nwell 17489 15967 17523 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_29.VPB
flabel pwell 17489 15423 17523 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_29.VNB
rlabel comment 17552 15440 17552 15440 6 sr_0.FILLER_0_6_29.decap_12
flabel metal1 16385 15423 16419 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_41.VGND
flabel metal1 16385 15967 16419 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_41.VPWR
flabel nwell 16385 15967 16419 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_41.VPB
flabel pwell 16385 15423 16419 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_41.VNB
rlabel comment 16448 15440 16448 15440 6 sr_0.FILLER_0_6_41.decap_12
flabel metal1 17673 16511 17707 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_27.VGND
flabel metal1 17673 15967 17707 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_27.VPWR
flabel nwell 17673 15967 17707 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_27.VPB
flabel pwell 17673 16511 17707 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_27.VNB
rlabel comment 17736 16528 17736 16528 8 sr_0.FILLER_0_7_27.decap_12
flabel metal1 16569 16511 16603 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_39.VGND
flabel metal1 16569 15967 16603 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_39.VPWR
flabel nwell 16569 15967 16603 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_39.VPB
flabel pwell 16569 16511 16603 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_39.VNB
rlabel comment 16632 16528 16632 16528 8 sr_0.FILLER_0_7_39.decap_12
flabel metal1 17569 15964 17622 15993 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_6_73.VPWR
flabel metal1 17572 15422 17623 15460 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_6_73.VGND
rlabel comment 17644 15440 17644 15440 6 sr_0.TAP_TAPCELL_ROW_6_73.tapvpwrvgnd_1
rlabel metal1 17552 15392 17644 15488 1 sr_0.TAP_TAPCELL_ROW_6_73.VGND
rlabel metal1 17552 15936 17644 16032 1 sr_0.TAP_TAPCELL_ROW_6_73.VPWR
flabel metal1 15281 15423 15315 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_53.VGND
flabel metal1 15281 15967 15315 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_53.VPWR
flabel nwell 15281 15967 15315 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_53.VPB
flabel pwell 15281 15423 15315 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_53.VNB
rlabel comment 15344 15440 15344 15440 6 sr_0.FILLER_0_6_53.decap_12
flabel metal1 15465 16511 15499 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_51.VGND
flabel metal1 15465 15967 15499 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_51.VPWR
flabel nwell 15465 15967 15499 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_51.VPB
flabel pwell 15465 16511 15499 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_51.VNB
rlabel comment 15528 16528 15528 16528 8 sr_0.FILLER_0_7_51.decap_4
rlabel metal1 15160 16480 15528 16576 5 sr_0.FILLER_0_7_51.VGND
rlabel metal1 15160 15936 15528 16032 5 sr_0.FILLER_0_7_51.VPWR
flabel metal1 15102 15971 15138 16001 0 FreeSans 250 0 0 0 sr_0.FILLER_0_7_55.VPWR
flabel metal1 15102 16512 15138 16541 0 FreeSans 250 0 0 0 sr_0.FILLER_0_7_55.VGND
flabel nwell 15109 15977 15129 15994 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_55.VPB
flabel pwell 15108 16517 15132 16539 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_55.VNB
rlabel comment 15160 16528 15160 16528 8 sr_0.FILLER_0_7_55.fill_1
rlabel metal1 15068 16480 15160 16576 5 sr_0.FILLER_0_7_55.VGND
rlabel metal1 15068 15936 15160 16032 5 sr_0.FILLER_0_7_55.VPWR
flabel metal1 14913 16511 14947 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_57.VGND
flabel metal1 14913 15967 14947 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_57.VPWR
flabel nwell 14913 15967 14947 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_57.VPB
flabel pwell 14913 16511 14947 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_57.VNB
rlabel comment 14976 16528 14976 16528 8 sr_0.FILLER_0_7_57.decap_12
flabel metal1 14993 15975 15046 16004 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_7_76.VPWR
flabel metal1 14996 16508 15047 16546 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_7_76.VGND
rlabel comment 15068 16528 15068 16528 8 sr_0.TAP_TAPCELL_ROW_7_76.tapvpwrvgnd_1
rlabel metal1 14976 16480 15068 16576 5 sr_0.TAP_TAPCELL_ROW_7_76.VGND
rlabel metal1 14976 15936 15068 16032 5 sr_0.TAP_TAPCELL_ROW_7_76.VPWR
flabel metal1 14177 15423 14211 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_65.VGND
flabel metal1 14177 15967 14211 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_65.VPWR
flabel nwell 14177 15967 14211 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_65.VPB
flabel pwell 14177 15423 14211 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_65.VNB
rlabel comment 14240 15440 14240 15440 6 sr_0.FILLER_0_6_65.decap_12
flabel metal1 13073 15967 13107 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_77.VPWR
flabel metal1 13073 15423 13107 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_77.VGND
flabel nwell 13073 15967 13107 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_77.VPB
flabel pwell 13073 15423 13107 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_77.VNB
rlabel comment 13136 15440 13136 15440 6 sr_0.FILLER_0_6_77.decap_6
rlabel metal1 12584 15392 13136 15488 1 sr_0.FILLER_0_6_77.VGND
rlabel metal1 12584 15936 13136 16032 1 sr_0.FILLER_0_6_77.VPWR
flabel metal1 12526 15967 12562 15997 0 FreeSans 250 0 0 0 sr_0.FILLER_0_6_83.VPWR
flabel metal1 12526 15427 12562 15456 0 FreeSans 250 0 0 0 sr_0.FILLER_0_6_83.VGND
flabel nwell 12533 15974 12553 15991 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_83.VPB
flabel pwell 12532 15429 12556 15451 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_83.VNB
rlabel comment 12584 15440 12584 15440 6 sr_0.FILLER_0_6_83.fill_1
rlabel metal1 12492 15392 12584 15488 1 sr_0.FILLER_0_6_83.VGND
rlabel metal1 12492 15936 12584 16032 1 sr_0.FILLER_0_6_83.VPWR
flabel metal1 13809 16511 13843 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_69.VGND
flabel metal1 13809 15967 13843 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_69.VPWR
flabel nwell 13809 15967 13843 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_69.VPB
flabel pwell 13809 16511 13843 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_69.VNB
rlabel comment 13872 16528 13872 16528 8 sr_0.FILLER_0_7_69.decap_12
flabel metal1 12705 16511 12739 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_81.VGND
flabel metal1 12705 15967 12739 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_81.VPWR
flabel nwell 12705 15967 12739 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_81.VPB
flabel pwell 12705 16511 12739 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_81.VNB
rlabel comment 12768 16528 12768 16528 8 sr_0.FILLER_0_7_81.decap_12
flabel metal1 12337 15423 12371 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_85.VGND
flabel metal1 12337 15967 12371 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_85.VPWR
flabel nwell 12337 15967 12371 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_85.VPB
flabel pwell 12337 15423 12371 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_85.VNB
rlabel comment 12400 15440 12400 15440 6 sr_0.FILLER_0_6_85.decap_12
flabel metal1 11233 15423 11267 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_97.VGND
flabel metal1 11233 15967 11267 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_97.VPWR
flabel nwell 11233 15967 11267 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_97.VPB
flabel pwell 11233 15423 11267 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_97.VNB
rlabel comment 11296 15440 11296 15440 6 sr_0.FILLER_0_6_97.decap_12
flabel metal1 11601 16511 11635 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_93.VGND
flabel metal1 11601 15967 11635 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_93.VPWR
flabel nwell 11601 15967 11635 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_93.VPB
flabel pwell 11601 16511 11635 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_93.VNB
rlabel comment 11664 16528 11664 16528 8 sr_0.FILLER_0_7_93.decap_12
flabel metal1 12417 15964 12470 15993 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_6_74.VPWR
flabel metal1 12420 15422 12471 15460 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_6_74.VGND
rlabel comment 12492 15440 12492 15440 6 sr_0.TAP_TAPCELL_ROW_6_74.tapvpwrvgnd_1
rlabel metal1 12400 15392 12492 15488 1 sr_0.TAP_TAPCELL_ROW_6_74.VGND
rlabel metal1 12400 15936 12492 16032 1 sr_0.TAP_TAPCELL_ROW_6_74.VPWR
flabel metal1 10129 15423 10163 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_109.VGND
flabel metal1 10129 15967 10163 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_109.VPWR
flabel nwell 10129 15967 10163 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_109.VPB
flabel pwell 10129 15423 10163 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_109.VNB
rlabel comment 10192 15440 10192 15440 6 sr_0.FILLER_0_6_109.decap_12
flabel metal1 9025 15423 9059 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_121.VGND
flabel metal1 9025 15967 9059 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_121.VPWR
flabel nwell 9025 15967 9059 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_121.VPB
flabel pwell 9025 15423 9059 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_121.VNB
rlabel comment 9088 15440 9088 15440 6 sr_0.FILLER_0_6_121.decap_12
flabel metal1 10497 15967 10531 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_105.VPWR
flabel metal1 10497 16511 10531 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_105.VGND
flabel nwell 10497 15967 10531 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_105.VPB
flabel pwell 10497 16511 10531 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_105.VNB
rlabel comment 10560 16528 10560 16528 8 sr_0.FILLER_0_7_105.decap_6
rlabel metal1 10008 16480 10560 16576 5 sr_0.FILLER_0_7_105.VGND
rlabel metal1 10008 15936 10560 16032 5 sr_0.FILLER_0_7_105.VPWR
flabel metal1 9950 15971 9986 16001 0 FreeSans 250 0 0 0 sr_0.FILLER_0_7_111.VPWR
flabel metal1 9950 16512 9986 16541 0 FreeSans 250 0 0 0 sr_0.FILLER_0_7_111.VGND
flabel nwell 9957 15977 9977 15994 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_111.VPB
flabel pwell 9956 16517 9980 16539 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_111.VNB
rlabel comment 10008 16528 10008 16528 8 sr_0.FILLER_0_7_111.fill_1
rlabel metal1 9916 16480 10008 16576 5 sr_0.FILLER_0_7_111.VGND
rlabel metal1 9916 15936 10008 16032 5 sr_0.FILLER_0_7_111.VPWR
flabel metal1 9761 16511 9795 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_113.VGND
flabel metal1 9761 15967 9795 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_113.VPWR
flabel nwell 9761 15967 9795 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_113.VPB
flabel pwell 9761 16511 9795 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_113.VNB
rlabel comment 9824 16528 9824 16528 8 sr_0.FILLER_0_7_113.decap_12
flabel metal1 8657 16511 8691 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_125.VGND
flabel metal1 8657 15967 8691 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_125.VPWR
flabel nwell 8657 15967 8691 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_125.VPB
flabel pwell 8657 16511 8691 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_125.VNB
rlabel comment 8720 16528 8720 16528 8 sr_0.FILLER_0_7_125.decap_12
flabel metal1 9841 15975 9894 16004 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_7_77.VPWR
flabel metal1 9844 16508 9895 16546 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_7_77.VGND
rlabel comment 9916 16528 9916 16528 8 sr_0.TAP_TAPCELL_ROW_7_77.tapvpwrvgnd_1
rlabel metal1 9824 16480 9916 16576 5 sr_0.TAP_TAPCELL_ROW_7_77.VGND
rlabel metal1 9824 15936 9916 16032 5 sr_0.TAP_TAPCELL_ROW_7_77.VPWR
flabel metal1 7921 15967 7955 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_133.VPWR
flabel metal1 7921 15423 7955 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_133.VGND
flabel nwell 7921 15967 7955 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_133.VPB
flabel pwell 7921 15423 7955 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_133.VNB
rlabel comment 7984 15440 7984 15440 6 sr_0.FILLER_0_6_133.decap_6
rlabel metal1 7432 15392 7984 15488 1 sr_0.FILLER_0_6_133.VGND
rlabel metal1 7432 15936 7984 16032 1 sr_0.FILLER_0_6_133.VPWR
flabel metal1 7374 15967 7410 15997 0 FreeSans 250 0 0 0 sr_0.FILLER_0_6_139.VPWR
flabel metal1 7374 15427 7410 15456 0 FreeSans 250 0 0 0 sr_0.FILLER_0_6_139.VGND
flabel nwell 7381 15974 7401 15991 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_139.VPB
flabel pwell 7380 15429 7404 15451 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_139.VNB
rlabel comment 7432 15440 7432 15440 6 sr_0.FILLER_0_6_139.fill_1
rlabel metal1 7340 15392 7432 15488 1 sr_0.FILLER_0_6_139.VGND
rlabel metal1 7340 15936 7432 16032 1 sr_0.FILLER_0_6_139.VPWR
flabel metal1 7185 15423 7219 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_141.VGND
flabel metal1 7185 15967 7219 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_141.VPWR
flabel nwell 7185 15967 7219 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_141.VPB
flabel pwell 7185 15423 7219 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_141.VNB
rlabel comment 7248 15440 7248 15440 6 sr_0.FILLER_0_6_141.decap_12
flabel metal1 7553 16511 7587 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_137.VGND
flabel metal1 7553 15967 7587 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_137.VPWR
flabel nwell 7553 15967 7587 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_137.VPB
flabel pwell 7553 16511 7587 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_137.VNB
rlabel comment 7616 16528 7616 16528 8 sr_0.FILLER_0_7_137.decap_12
flabel metal1 7265 15964 7318 15993 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_6_75.VPWR
flabel metal1 7268 15422 7319 15460 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_6_75.VGND
rlabel comment 7340 15440 7340 15440 6 sr_0.TAP_TAPCELL_ROW_6_75.tapvpwrvgnd_1
rlabel metal1 7248 15392 7340 15488 1 sr_0.TAP_TAPCELL_ROW_6_75.VGND
rlabel metal1 7248 15936 7340 16032 1 sr_0.TAP_TAPCELL_ROW_6_75.VPWR
flabel metal1 6081 15967 6115 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_153.VPWR
flabel metal1 6081 15423 6115 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_153.VGND
flabel nwell 6081 15967 6115 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_153.VPB
flabel pwell 6081 15423 6115 15457 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_153.VNB
rlabel comment 6144 15440 6144 15440 6 sr_0.FILLER_0_6_153.decap_8
rlabel metal1 5408 15392 6144 15488 1 sr_0.FILLER_0_6_153.VGND
rlabel metal1 5408 15936 6144 16032 1 sr_0.FILLER_0_6_153.VPWR
flabel metal1 5335 15426 5388 15458 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_161.VGND
flabel metal1 5335 15970 5387 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_161.VPWR
flabel nwell 5346 15975 5380 15993 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_161.VPB
flabel pwell 5345 15430 5377 15452 0 FreeSans 200 0 0 0 sr_0.FILLER_0_6_161.VNB
rlabel comment 5408 15440 5408 15440 6 sr_0.FILLER_0_6_161.fill_2
rlabel metal1 5224 15392 5408 15488 1 sr_0.FILLER_0_6_161.VGND
rlabel metal1 5224 15936 5408 16032 1 sr_0.FILLER_0_6_161.VPWR
flabel metal1 6449 16511 6483 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_149.VGND
flabel metal1 6449 15967 6483 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_149.VPWR
flabel nwell 6449 15967 6483 16001 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_149.VPB
flabel pwell 6449 16511 6483 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_149.VNB
rlabel comment 6512 16528 6512 16528 8 sr_0.FILLER_0_7_149.decap_12
flabel metal1 5335 16510 5388 16542 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_161.VGND
flabel metal1 5335 15967 5387 15998 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_161.VPWR
flabel nwell 5346 15975 5380 15993 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_161.VPB
flabel pwell 5345 16516 5377 16538 0 FreeSans 200 0 0 0 sr_0.FILLER_0_7_161.VNB
rlabel comment 5408 16528 5408 16528 8 sr_0.FILLER_0_7_161.fill_2
rlabel metal1 5224 16480 5408 16576 5 sr_0.FILLER_0_7_161.VGND
rlabel metal1 5224 15936 5408 16032 5 sr_0.FILLER_0_7_161.VPWR
flabel metal1 4977 15967 5011 16001 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_6_Right_6.VPWR
flabel metal1 4977 15423 5011 15457 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_6_Right_6.VGND
flabel nwell 4977 15967 5011 16001 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_6_Right_6.VPB
flabel pwell 4977 15423 5011 15457 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_6_Right_6.VNB
rlabel comment 4948 15440 4948 15440 4 sr_0.PHY_EDGE_ROW_6_Right_6.decap_3
rlabel metal1 4948 15392 5224 15488 1 sr_0.PHY_EDGE_ROW_6_Right_6.VGND
rlabel metal1 4948 15936 5224 16032 1 sr_0.PHY_EDGE_ROW_6_Right_6.VPWR
flabel metal1 4977 15967 5011 16001 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_7_Right_7.VPWR
flabel metal1 4977 16511 5011 16545 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_7_Right_7.VGND
flabel nwell 4977 15967 5011 16001 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_7_Right_7.VPB
flabel pwell 4977 16511 5011 16545 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_7_Right_7.VNB
rlabel comment 4948 16528 4948 16528 2 sr_0.PHY_EDGE_ROW_7_Right_7.decap_3
rlabel metal1 4948 16480 5224 16576 5 sr_0.PHY_EDGE_ROW_7_Right_7.VGND
rlabel metal1 4948 15936 5224 16032 5 sr_0.PHY_EDGE_ROW_7_Right_7.VPWR
flabel metal1 19881 16511 19915 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_3.VGND
flabel metal1 19881 17055 19915 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_3.VPWR
flabel nwell 19881 17055 19915 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_3.VPB
flabel pwell 19881 16511 19915 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_3.VNB
rlabel comment 19944 16528 19944 16528 6 sr_0.FILLER_0_8_3.decap_12
flabel metal1 18777 16511 18811 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_15.VGND
flabel metal1 18777 17055 18811 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_15.VPWR
flabel nwell 18777 17055 18811 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_15.VPB
flabel pwell 18777 16511 18811 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_15.VNB
rlabel comment 18840 16528 18840 16528 6 sr_0.FILLER_0_8_15.decap_12
flabel metal1 20157 17055 20191 17089 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_8_Left_36.VPWR
flabel metal1 20157 16511 20191 16545 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_8_Left_36.VGND
flabel nwell 20157 17055 20191 17089 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_8_Left_36.VPB
flabel pwell 20157 16511 20191 16545 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_8_Left_36.VNB
rlabel comment 20220 16528 20220 16528 6 sr_0.PHY_EDGE_ROW_8_Left_36.decap_3
rlabel metal1 19944 16480 20220 16576 1 sr_0.PHY_EDGE_ROW_8_Left_36.VGND
rlabel metal1 19944 17024 20220 17120 1 sr_0.PHY_EDGE_ROW_8_Left_36.VPWR
flabel metal1 17678 17055 17714 17085 0 FreeSans 250 0 0 0 sr_0.FILLER_0_8_27.VPWR
flabel metal1 17678 16515 17714 16544 0 FreeSans 250 0 0 0 sr_0.FILLER_0_8_27.VGND
flabel nwell 17685 17062 17705 17079 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_27.VPB
flabel pwell 17684 16517 17708 16539 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_27.VNB
rlabel comment 17736 16528 17736 16528 6 sr_0.FILLER_0_8_27.fill_1
rlabel metal1 17644 16480 17736 16576 1 sr_0.FILLER_0_8_27.VGND
rlabel metal1 17644 17024 17736 17120 1 sr_0.FILLER_0_8_27.VPWR
flabel metal1 17489 16511 17523 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_29.VGND
flabel metal1 17489 17055 17523 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_29.VPWR
flabel nwell 17489 17055 17523 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_29.VPB
flabel pwell 17489 16511 17523 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_29.VNB
rlabel comment 17552 16528 17552 16528 6 sr_0.FILLER_0_8_29.decap_12
flabel metal1 16385 16511 16419 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_41.VGND
flabel metal1 16385 17055 16419 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_41.VPWR
flabel nwell 16385 17055 16419 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_41.VPB
flabel pwell 16385 16511 16419 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_41.VNB
rlabel comment 16448 16528 16448 16528 6 sr_0.FILLER_0_8_41.decap_12
flabel metal1 17569 17052 17622 17081 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_8_78.VPWR
flabel metal1 17572 16510 17623 16548 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_8_78.VGND
rlabel comment 17644 16528 17644 16528 6 sr_0.TAP_TAPCELL_ROW_8_78.tapvpwrvgnd_1
rlabel metal1 17552 16480 17644 16576 1 sr_0.TAP_TAPCELL_ROW_8_78.VGND
rlabel metal1 17552 17024 17644 17120 1 sr_0.TAP_TAPCELL_ROW_8_78.VPWR
flabel metal1 15281 16511 15315 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_53.VGND
flabel metal1 15281 17055 15315 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_53.VPWR
flabel nwell 15281 17055 15315 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_53.VPB
flabel pwell 15281 16511 15315 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_53.VNB
rlabel comment 15344 16528 15344 16528 6 sr_0.FILLER_0_8_53.decap_12
flabel metal1 14177 16511 14211 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_65.VGND
flabel metal1 14177 17055 14211 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_65.VPWR
flabel nwell 14177 17055 14211 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_65.VPB
flabel pwell 14177 16511 14211 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_65.VNB
rlabel comment 14240 16528 14240 16528 6 sr_0.FILLER_0_8_65.decap_12
flabel metal1 13073 17055 13107 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_77.VPWR
flabel metal1 13073 16511 13107 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_77.VGND
flabel nwell 13073 17055 13107 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_77.VPB
flabel pwell 13073 16511 13107 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_77.VNB
rlabel comment 13136 16528 13136 16528 6 sr_0.FILLER_0_8_77.decap_6
rlabel metal1 12584 16480 13136 16576 1 sr_0.FILLER_0_8_77.VGND
rlabel metal1 12584 17024 13136 17120 1 sr_0.FILLER_0_8_77.VPWR
flabel metal1 12526 17055 12562 17085 0 FreeSans 250 0 0 0 sr_0.FILLER_0_8_83.VPWR
flabel metal1 12526 16515 12562 16544 0 FreeSans 250 0 0 0 sr_0.FILLER_0_8_83.VGND
flabel nwell 12533 17062 12553 17079 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_83.VPB
flabel pwell 12532 16517 12556 16539 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_83.VNB
rlabel comment 12584 16528 12584 16528 6 sr_0.FILLER_0_8_83.fill_1
rlabel metal1 12492 16480 12584 16576 1 sr_0.FILLER_0_8_83.VGND
rlabel metal1 12492 17024 12584 17120 1 sr_0.FILLER_0_8_83.VPWR
flabel metal1 12337 16511 12371 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_85.VGND
flabel metal1 12337 17055 12371 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_85.VPWR
flabel nwell 12337 17055 12371 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_85.VPB
flabel pwell 12337 16511 12371 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_85.VNB
rlabel comment 12400 16528 12400 16528 6 sr_0.FILLER_0_8_85.decap_12
flabel metal1 11233 16511 11267 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_97.VGND
flabel metal1 11233 17055 11267 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_97.VPWR
flabel nwell 11233 17055 11267 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_97.VPB
flabel pwell 11233 16511 11267 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_97.VNB
rlabel comment 11296 16528 11296 16528 6 sr_0.FILLER_0_8_97.decap_12
flabel metal1 12417 17052 12470 17081 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_8_79.VPWR
flabel metal1 12420 16510 12471 16548 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_8_79.VGND
rlabel comment 12492 16528 12492 16528 6 sr_0.TAP_TAPCELL_ROW_8_79.tapvpwrvgnd_1
rlabel metal1 12400 16480 12492 16576 1 sr_0.TAP_TAPCELL_ROW_8_79.VGND
rlabel metal1 12400 17024 12492 17120 1 sr_0.TAP_TAPCELL_ROW_8_79.VPWR
flabel metal1 10129 16511 10163 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_109.VGND
flabel metal1 10129 17055 10163 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_109.VPWR
flabel nwell 10129 17055 10163 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_109.VPB
flabel pwell 10129 16511 10163 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_109.VNB
rlabel comment 10192 16528 10192 16528 6 sr_0.FILLER_0_8_109.decap_12
flabel metal1 9025 16511 9059 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_121.VGND
flabel metal1 9025 17055 9059 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_121.VPWR
flabel nwell 9025 17055 9059 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_121.VPB
flabel pwell 9025 16511 9059 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_121.VNB
rlabel comment 9088 16528 9088 16528 6 sr_0.FILLER_0_8_121.decap_12
flabel metal1 7921 17055 7955 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_133.VPWR
flabel metal1 7921 16511 7955 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_133.VGND
flabel nwell 7921 17055 7955 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_133.VPB
flabel pwell 7921 16511 7955 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_133.VNB
rlabel comment 7984 16528 7984 16528 6 sr_0.FILLER_0_8_133.decap_6
rlabel metal1 7432 16480 7984 16576 1 sr_0.FILLER_0_8_133.VGND
rlabel metal1 7432 17024 7984 17120 1 sr_0.FILLER_0_8_133.VPWR
flabel metal1 7374 17055 7410 17085 0 FreeSans 250 0 0 0 sr_0.FILLER_0_8_139.VPWR
flabel metal1 7374 16515 7410 16544 0 FreeSans 250 0 0 0 sr_0.FILLER_0_8_139.VGND
flabel nwell 7381 17062 7401 17079 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_139.VPB
flabel pwell 7380 16517 7404 16539 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_139.VNB
rlabel comment 7432 16528 7432 16528 6 sr_0.FILLER_0_8_139.fill_1
rlabel metal1 7340 16480 7432 16576 1 sr_0.FILLER_0_8_139.VGND
rlabel metal1 7340 17024 7432 17120 1 sr_0.FILLER_0_8_139.VPWR
flabel metal1 7185 16511 7219 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_141.VGND
flabel metal1 7185 17055 7219 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_141.VPWR
flabel nwell 7185 17055 7219 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_141.VPB
flabel pwell 7185 16511 7219 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_141.VNB
rlabel comment 7248 16528 7248 16528 6 sr_0.FILLER_0_8_141.decap_12
flabel metal1 7265 17052 7318 17081 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_8_80.VPWR
flabel metal1 7268 16510 7319 16548 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_8_80.VGND
rlabel comment 7340 16528 7340 16528 6 sr_0.TAP_TAPCELL_ROW_8_80.tapvpwrvgnd_1
rlabel metal1 7248 16480 7340 16576 1 sr_0.TAP_TAPCELL_ROW_8_80.VGND
rlabel metal1 7248 17024 7340 17120 1 sr_0.TAP_TAPCELL_ROW_8_80.VPWR
flabel metal1 6081 17055 6115 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_153.VPWR
flabel metal1 6081 16511 6115 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_153.VGND
flabel nwell 6081 17055 6115 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_153.VPB
flabel pwell 6081 16511 6115 16545 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_153.VNB
rlabel comment 6144 16528 6144 16528 6 sr_0.FILLER_0_8_153.decap_8
rlabel metal1 5408 16480 6144 16576 1 sr_0.FILLER_0_8_153.VGND
rlabel metal1 5408 17024 6144 17120 1 sr_0.FILLER_0_8_153.VPWR
flabel metal1 5335 16514 5388 16546 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_161.VGND
flabel metal1 5335 17058 5387 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_161.VPWR
flabel nwell 5346 17063 5380 17081 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_161.VPB
flabel pwell 5345 16518 5377 16540 0 FreeSans 200 0 0 0 sr_0.FILLER_0_8_161.VNB
rlabel comment 5408 16528 5408 16528 6 sr_0.FILLER_0_8_161.fill_2
rlabel metal1 5224 16480 5408 16576 1 sr_0.FILLER_0_8_161.VGND
rlabel metal1 5224 17024 5408 17120 1 sr_0.FILLER_0_8_161.VPWR
flabel metal1 4977 17055 5011 17089 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_8_Right_8.VPWR
flabel metal1 4977 16511 5011 16545 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_8_Right_8.VGND
flabel nwell 4977 17055 5011 17089 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_8_Right_8.VPB
flabel pwell 4977 16511 5011 16545 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_8_Right_8.VNB
rlabel comment 4948 16528 4948 16528 4 sr_0.PHY_EDGE_ROW_8_Right_8.decap_3
rlabel metal1 4948 16480 5224 16576 1 sr_0.PHY_EDGE_ROW_8_Right_8.VGND
rlabel metal1 4948 17024 5224 17120 1 sr_0.PHY_EDGE_ROW_8_Right_8.VPWR
flabel metal1 19881 17599 19915 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_3.VGND
flabel metal1 19881 17055 19915 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_3.VPWR
flabel nwell 19881 17055 19915 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_3.VPB
flabel pwell 19881 17599 19915 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_3.VNB
rlabel comment 19944 17616 19944 17616 8 sr_0.FILLER_0_9_3.decap_12
flabel metal1 18777 17599 18811 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_15.VGND
flabel metal1 18777 17055 18811 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_15.VPWR
flabel nwell 18777 17055 18811 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_15.VPB
flabel pwell 18777 17599 18811 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_15.VNB
rlabel comment 18840 17616 18840 17616 8 sr_0.FILLER_0_9_15.decap_12
flabel metal1 20157 17055 20191 17089 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_9_Left_37.VPWR
flabel metal1 20157 17599 20191 17633 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_9_Left_37.VGND
flabel nwell 20157 17055 20191 17089 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_9_Left_37.VPB
flabel pwell 20157 17599 20191 17633 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_9_Left_37.VNB
rlabel comment 20220 17616 20220 17616 8 sr_0.PHY_EDGE_ROW_9_Left_37.decap_3
rlabel metal1 19944 17568 20220 17664 5 sr_0.PHY_EDGE_ROW_9_Left_37.VGND
rlabel metal1 19944 17024 20220 17120 5 sr_0.PHY_EDGE_ROW_9_Left_37.VPWR
flabel metal1 17673 17599 17707 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_27.VGND
flabel metal1 17673 17055 17707 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_27.VPWR
flabel nwell 17673 17055 17707 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_27.VPB
flabel pwell 17673 17599 17707 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_27.VNB
rlabel comment 17736 17616 17736 17616 8 sr_0.FILLER_0_9_27.decap_12
flabel metal1 16569 17599 16603 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_39.VGND
flabel metal1 16569 17055 16603 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_39.VPWR
flabel nwell 16569 17055 16603 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_39.VPB
flabel pwell 16569 17599 16603 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_39.VNB
rlabel comment 16632 17616 16632 17616 8 sr_0.FILLER_0_9_39.decap_12
flabel metal1 15465 17599 15499 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_51.VGND
flabel metal1 15465 17055 15499 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_51.VPWR
flabel nwell 15465 17055 15499 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_51.VPB
flabel pwell 15465 17599 15499 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_51.VNB
rlabel comment 15528 17616 15528 17616 8 sr_0.FILLER_0_9_51.decap_4
rlabel metal1 15160 17568 15528 17664 5 sr_0.FILLER_0_9_51.VGND
rlabel metal1 15160 17024 15528 17120 5 sr_0.FILLER_0_9_51.VPWR
flabel metal1 15102 17059 15138 17089 0 FreeSans 250 0 0 0 sr_0.FILLER_0_9_55.VPWR
flabel metal1 15102 17600 15138 17629 0 FreeSans 250 0 0 0 sr_0.FILLER_0_9_55.VGND
flabel nwell 15109 17065 15129 17082 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_55.VPB
flabel pwell 15108 17605 15132 17627 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_55.VNB
rlabel comment 15160 17616 15160 17616 8 sr_0.FILLER_0_9_55.fill_1
rlabel metal1 15068 17568 15160 17664 5 sr_0.FILLER_0_9_55.VGND
rlabel metal1 15068 17024 15160 17120 5 sr_0.FILLER_0_9_55.VPWR
flabel metal1 14913 17599 14947 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_57.VGND
flabel metal1 14913 17055 14947 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_57.VPWR
flabel nwell 14913 17055 14947 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_57.VPB
flabel pwell 14913 17599 14947 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_57.VNB
rlabel comment 14976 17616 14976 17616 8 sr_0.FILLER_0_9_57.decap_12
flabel metal1 14993 17063 15046 17092 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_9_81.VPWR
flabel metal1 14996 17596 15047 17634 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_9_81.VGND
rlabel comment 15068 17616 15068 17616 8 sr_0.TAP_TAPCELL_ROW_9_81.tapvpwrvgnd_1
rlabel metal1 14976 17568 15068 17664 5 sr_0.TAP_TAPCELL_ROW_9_81.VGND
rlabel metal1 14976 17024 15068 17120 5 sr_0.TAP_TAPCELL_ROW_9_81.VPWR
flabel metal1 13809 17599 13843 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_69.VGND
flabel metal1 13809 17055 13843 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_69.VPWR
flabel nwell 13809 17055 13843 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_69.VPB
flabel pwell 13809 17599 13843 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_69.VNB
rlabel comment 13872 17616 13872 17616 8 sr_0.FILLER_0_9_69.decap_12
flabel metal1 12705 17599 12739 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_81.VGND
flabel metal1 12705 17055 12739 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_81.VPWR
flabel nwell 12705 17055 12739 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_81.VPB
flabel pwell 12705 17599 12739 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_81.VNB
rlabel comment 12768 17616 12768 17616 8 sr_0.FILLER_0_9_81.decap_12
flabel metal1 11601 17599 11635 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_93.VGND
flabel metal1 11601 17055 11635 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_93.VPWR
flabel nwell 11601 17055 11635 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_93.VPB
flabel pwell 11601 17599 11635 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_93.VNB
rlabel comment 11664 17616 11664 17616 8 sr_0.FILLER_0_9_93.decap_12
flabel metal1 10497 17055 10531 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_105.VPWR
flabel metal1 10497 17599 10531 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_105.VGND
flabel nwell 10497 17055 10531 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_105.VPB
flabel pwell 10497 17599 10531 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_105.VNB
rlabel comment 10560 17616 10560 17616 8 sr_0.FILLER_0_9_105.decap_6
rlabel metal1 10008 17568 10560 17664 5 sr_0.FILLER_0_9_105.VGND
rlabel metal1 10008 17024 10560 17120 5 sr_0.FILLER_0_9_105.VPWR
flabel metal1 9950 17059 9986 17089 0 FreeSans 250 0 0 0 sr_0.FILLER_0_9_111.VPWR
flabel metal1 9950 17600 9986 17629 0 FreeSans 250 0 0 0 sr_0.FILLER_0_9_111.VGND
flabel nwell 9957 17065 9977 17082 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_111.VPB
flabel pwell 9956 17605 9980 17627 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_111.VNB
rlabel comment 10008 17616 10008 17616 8 sr_0.FILLER_0_9_111.fill_1
rlabel metal1 9916 17568 10008 17664 5 sr_0.FILLER_0_9_111.VGND
rlabel metal1 9916 17024 10008 17120 5 sr_0.FILLER_0_9_111.VPWR
flabel metal1 9761 17599 9795 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_113.VGND
flabel metal1 9761 17055 9795 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_113.VPWR
flabel nwell 9761 17055 9795 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_113.VPB
flabel pwell 9761 17599 9795 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_113.VNB
rlabel comment 9824 17616 9824 17616 8 sr_0.FILLER_0_9_113.decap_12
flabel metal1 8657 17599 8691 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_125.VGND
flabel metal1 8657 17055 8691 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_125.VPWR
flabel nwell 8657 17055 8691 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_125.VPB
flabel pwell 8657 17599 8691 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_125.VNB
rlabel comment 8720 17616 8720 17616 8 sr_0.FILLER_0_9_125.decap_12
flabel metal1 9841 17063 9894 17092 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_9_82.VPWR
flabel metal1 9844 17596 9895 17634 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_9_82.VGND
rlabel comment 9916 17616 9916 17616 8 sr_0.TAP_TAPCELL_ROW_9_82.tapvpwrvgnd_1
rlabel metal1 9824 17568 9916 17664 5 sr_0.TAP_TAPCELL_ROW_9_82.VGND
rlabel metal1 9824 17024 9916 17120 5 sr_0.TAP_TAPCELL_ROW_9_82.VPWR
flabel metal1 7553 17599 7587 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_137.VGND
flabel metal1 7553 17055 7587 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_137.VPWR
flabel nwell 7553 17055 7587 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_137.VPB
flabel pwell 7553 17599 7587 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_137.VNB
rlabel comment 7616 17616 7616 17616 8 sr_0.FILLER_0_9_137.decap_12
flabel metal1 6449 17599 6483 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_149.VGND
flabel metal1 6449 17055 6483 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_149.VPWR
flabel nwell 6449 17055 6483 17089 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_149.VPB
flabel pwell 6449 17599 6483 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_149.VNB
rlabel comment 6512 17616 6512 17616 8 sr_0.FILLER_0_9_149.decap_12
flabel metal1 5335 17598 5388 17630 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_161.VGND
flabel metal1 5335 17055 5387 17086 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_161.VPWR
flabel nwell 5346 17063 5380 17081 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_161.VPB
flabel pwell 5345 17604 5377 17626 0 FreeSans 200 0 0 0 sr_0.FILLER_0_9_161.VNB
rlabel comment 5408 17616 5408 17616 8 sr_0.FILLER_0_9_161.fill_2
rlabel metal1 5224 17568 5408 17664 5 sr_0.FILLER_0_9_161.VGND
rlabel metal1 5224 17024 5408 17120 5 sr_0.FILLER_0_9_161.VPWR
flabel metal1 4977 17055 5011 17089 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_9_Right_9.VPWR
flabel metal1 4977 17599 5011 17633 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_9_Right_9.VGND
flabel nwell 4977 17055 5011 17089 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_9_Right_9.VPB
flabel pwell 4977 17599 5011 17633 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_9_Right_9.VNB
rlabel comment 4948 17616 4948 17616 2 sr_0.PHY_EDGE_ROW_9_Right_9.decap_3
rlabel metal1 4948 17568 5224 17664 5 sr_0.PHY_EDGE_ROW_9_Right_9.VGND
rlabel metal1 4948 17024 5224 17120 5 sr_0.PHY_EDGE_ROW_9_Right_9.VPWR
flabel metal1 19881 17599 19915 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_3.VGND
flabel metal1 19881 18143 19915 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_3.VPWR
flabel nwell 19881 18143 19915 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_3.VPB
flabel pwell 19881 17599 19915 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_3.VNB
rlabel comment 19944 17616 19944 17616 6 sr_0.FILLER_0_10_3.decap_12
flabel metal1 18777 17599 18811 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_15.VGND
flabel metal1 18777 18143 18811 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_15.VPWR
flabel nwell 18777 18143 18811 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_15.VPB
flabel pwell 18777 17599 18811 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_15.VNB
rlabel comment 18840 17616 18840 17616 6 sr_0.FILLER_0_10_15.decap_12
flabel metal1 20157 18143 20191 18177 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_10_Left_38.VPWR
flabel metal1 20157 17599 20191 17633 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_10_Left_38.VGND
flabel nwell 20157 18143 20191 18177 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_10_Left_38.VPB
flabel pwell 20157 17599 20191 17633 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_10_Left_38.VNB
rlabel comment 20220 17616 20220 17616 6 sr_0.PHY_EDGE_ROW_10_Left_38.decap_3
rlabel metal1 19944 17568 20220 17664 1 sr_0.PHY_EDGE_ROW_10_Left_38.VGND
rlabel metal1 19944 18112 20220 18208 1 sr_0.PHY_EDGE_ROW_10_Left_38.VPWR
flabel metal1 17678 18143 17714 18173 0 FreeSans 250 0 0 0 sr_0.FILLER_0_10_27.VPWR
flabel metal1 17678 17603 17714 17632 0 FreeSans 250 0 0 0 sr_0.FILLER_0_10_27.VGND
flabel nwell 17685 18150 17705 18167 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_27.VPB
flabel pwell 17684 17605 17708 17627 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_27.VNB
rlabel comment 17736 17616 17736 17616 6 sr_0.FILLER_0_10_27.fill_1
rlabel metal1 17644 17568 17736 17664 1 sr_0.FILLER_0_10_27.VGND
rlabel metal1 17644 18112 17736 18208 1 sr_0.FILLER_0_10_27.VPWR
flabel metal1 17489 17599 17523 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_29.VGND
flabel metal1 17489 18143 17523 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_29.VPWR
flabel nwell 17489 18143 17523 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_29.VPB
flabel pwell 17489 17599 17523 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_29.VNB
rlabel comment 17552 17616 17552 17616 6 sr_0.FILLER_0_10_29.decap_12
flabel metal1 16385 17599 16419 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_41.VGND
flabel metal1 16385 18143 16419 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_41.VPWR
flabel nwell 16385 18143 16419 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_41.VPB
flabel pwell 16385 17599 16419 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_41.VNB
rlabel comment 16448 17616 16448 17616 6 sr_0.FILLER_0_10_41.decap_12
flabel metal1 17569 18140 17622 18169 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_10_83.VPWR
flabel metal1 17572 17598 17623 17636 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_10_83.VGND
rlabel comment 17644 17616 17644 17616 6 sr_0.TAP_TAPCELL_ROW_10_83.tapvpwrvgnd_1
rlabel metal1 17552 17568 17644 17664 1 sr_0.TAP_TAPCELL_ROW_10_83.VGND
rlabel metal1 17552 18112 17644 18208 1 sr_0.TAP_TAPCELL_ROW_10_83.VPWR
flabel metal1 15281 17599 15315 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_53.VGND
flabel metal1 15281 18143 15315 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_53.VPWR
flabel nwell 15281 18143 15315 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_53.VPB
flabel pwell 15281 17599 15315 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_53.VNB
rlabel comment 15344 17616 15344 17616 6 sr_0.FILLER_0_10_53.decap_12
flabel metal1 14177 17599 14211 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_65.VGND
flabel metal1 14177 18143 14211 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_65.VPWR
flabel nwell 14177 18143 14211 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_65.VPB
flabel pwell 14177 17599 14211 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_65.VNB
rlabel comment 14240 17616 14240 17616 6 sr_0.FILLER_0_10_65.decap_12
flabel metal1 13073 18143 13107 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_77.VPWR
flabel metal1 13073 17599 13107 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_77.VGND
flabel nwell 13073 18143 13107 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_77.VPB
flabel pwell 13073 17599 13107 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_77.VNB
rlabel comment 13136 17616 13136 17616 6 sr_0.FILLER_0_10_77.decap_6
rlabel metal1 12584 17568 13136 17664 1 sr_0.FILLER_0_10_77.VGND
rlabel metal1 12584 18112 13136 18208 1 sr_0.FILLER_0_10_77.VPWR
flabel metal1 12526 18143 12562 18173 0 FreeSans 250 0 0 0 sr_0.FILLER_0_10_83.VPWR
flabel metal1 12526 17603 12562 17632 0 FreeSans 250 0 0 0 sr_0.FILLER_0_10_83.VGND
flabel nwell 12533 18150 12553 18167 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_83.VPB
flabel pwell 12532 17605 12556 17627 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_83.VNB
rlabel comment 12584 17616 12584 17616 6 sr_0.FILLER_0_10_83.fill_1
rlabel metal1 12492 17568 12584 17664 1 sr_0.FILLER_0_10_83.VGND
rlabel metal1 12492 18112 12584 18208 1 sr_0.FILLER_0_10_83.VPWR
flabel metal1 12337 17599 12371 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_85.VGND
flabel metal1 12337 18143 12371 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_85.VPWR
flabel nwell 12337 18143 12371 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_85.VPB
flabel pwell 12337 17599 12371 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_85.VNB
rlabel comment 12400 17616 12400 17616 6 sr_0.FILLER_0_10_85.decap_12
flabel metal1 11233 17599 11267 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_97.VGND
flabel metal1 11233 18143 11267 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_97.VPWR
flabel nwell 11233 18143 11267 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_97.VPB
flabel pwell 11233 17599 11267 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_97.VNB
rlabel comment 11296 17616 11296 17616 6 sr_0.FILLER_0_10_97.decap_12
flabel metal1 12417 18140 12470 18169 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_10_84.VPWR
flabel metal1 12420 17598 12471 17636 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_10_84.VGND
rlabel comment 12492 17616 12492 17616 6 sr_0.TAP_TAPCELL_ROW_10_84.tapvpwrvgnd_1
rlabel metal1 12400 17568 12492 17664 1 sr_0.TAP_TAPCELL_ROW_10_84.VGND
rlabel metal1 12400 18112 12492 18208 1 sr_0.TAP_TAPCELL_ROW_10_84.VPWR
flabel metal1 10129 17599 10163 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_109.VGND
flabel metal1 10129 18143 10163 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_109.VPWR
flabel nwell 10129 18143 10163 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_109.VPB
flabel pwell 10129 17599 10163 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_109.VNB
rlabel comment 10192 17616 10192 17616 6 sr_0.FILLER_0_10_109.decap_12
flabel metal1 9025 17599 9059 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_121.VGND
flabel metal1 9025 18143 9059 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_121.VPWR
flabel nwell 9025 18143 9059 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_121.VPB
flabel pwell 9025 17599 9059 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_121.VNB
rlabel comment 9088 17616 9088 17616 6 sr_0.FILLER_0_10_121.decap_12
flabel metal1 7921 18143 7955 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_133.VPWR
flabel metal1 7921 17599 7955 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_133.VGND
flabel nwell 7921 18143 7955 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_133.VPB
flabel pwell 7921 17599 7955 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_133.VNB
rlabel comment 7984 17616 7984 17616 6 sr_0.FILLER_0_10_133.decap_6
rlabel metal1 7432 17568 7984 17664 1 sr_0.FILLER_0_10_133.VGND
rlabel metal1 7432 18112 7984 18208 1 sr_0.FILLER_0_10_133.VPWR
flabel metal1 7374 18143 7410 18173 0 FreeSans 250 0 0 0 sr_0.FILLER_0_10_139.VPWR
flabel metal1 7374 17603 7410 17632 0 FreeSans 250 0 0 0 sr_0.FILLER_0_10_139.VGND
flabel nwell 7381 18150 7401 18167 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_139.VPB
flabel pwell 7380 17605 7404 17627 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_139.VNB
rlabel comment 7432 17616 7432 17616 6 sr_0.FILLER_0_10_139.fill_1
rlabel metal1 7340 17568 7432 17664 1 sr_0.FILLER_0_10_139.VGND
rlabel metal1 7340 18112 7432 18208 1 sr_0.FILLER_0_10_139.VPWR
flabel metal1 7185 17599 7219 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_141.VGND
flabel metal1 7185 18143 7219 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_141.VPWR
flabel nwell 7185 18143 7219 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_141.VPB
flabel pwell 7185 17599 7219 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_141.VNB
rlabel comment 7248 17616 7248 17616 6 sr_0.FILLER_0_10_141.decap_12
flabel metal1 7265 18140 7318 18169 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_10_85.VPWR
flabel metal1 7268 17598 7319 17636 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_10_85.VGND
rlabel comment 7340 17616 7340 17616 6 sr_0.TAP_TAPCELL_ROW_10_85.tapvpwrvgnd_1
rlabel metal1 7248 17568 7340 17664 1 sr_0.TAP_TAPCELL_ROW_10_85.VGND
rlabel metal1 7248 18112 7340 18208 1 sr_0.TAP_TAPCELL_ROW_10_85.VPWR
flabel metal1 6081 18143 6115 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_153.VPWR
flabel metal1 6081 17599 6115 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_153.VGND
flabel nwell 6081 18143 6115 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_153.VPB
flabel pwell 6081 17599 6115 17633 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_153.VNB
rlabel comment 6144 17616 6144 17616 6 sr_0.FILLER_0_10_153.decap_8
rlabel metal1 5408 17568 6144 17664 1 sr_0.FILLER_0_10_153.VGND
rlabel metal1 5408 18112 6144 18208 1 sr_0.FILLER_0_10_153.VPWR
flabel metal1 5335 17602 5388 17634 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_161.VGND
flabel metal1 5335 18146 5387 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_161.VPWR
flabel nwell 5346 18151 5380 18169 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_161.VPB
flabel pwell 5345 17606 5377 17628 0 FreeSans 200 0 0 0 sr_0.FILLER_0_10_161.VNB
rlabel comment 5408 17616 5408 17616 6 sr_0.FILLER_0_10_161.fill_2
rlabel metal1 5224 17568 5408 17664 1 sr_0.FILLER_0_10_161.VGND
rlabel metal1 5224 18112 5408 18208 1 sr_0.FILLER_0_10_161.VPWR
flabel metal1 4977 18143 5011 18177 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_10_Right_10.VPWR
flabel metal1 4977 17599 5011 17633 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_10_Right_10.VGND
flabel nwell 4977 18143 5011 18177 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_10_Right_10.VPB
flabel pwell 4977 17599 5011 17633 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_10_Right_10.VNB
rlabel comment 4948 17616 4948 17616 4 sr_0.PHY_EDGE_ROW_10_Right_10.decap_3
rlabel metal1 4948 17568 5224 17664 1 sr_0.PHY_EDGE_ROW_10_Right_10.VGND
rlabel metal1 4948 18112 5224 18208 1 sr_0.PHY_EDGE_ROW_10_Right_10.VPWR
flabel metal1 19881 18687 19915 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_3.VGND
flabel metal1 19881 18143 19915 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_3.VPWR
flabel nwell 19881 18143 19915 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_3.VPB
flabel pwell 19881 18687 19915 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_3.VNB
rlabel comment 19944 18704 19944 18704 8 sr_0.FILLER_0_11_3.decap_12
flabel metal1 18777 18687 18811 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_15.VGND
flabel metal1 18777 18143 18811 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_15.VPWR
flabel nwell 18777 18143 18811 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_15.VPB
flabel pwell 18777 18687 18811 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_15.VNB
rlabel comment 18840 18704 18840 18704 8 sr_0.FILLER_0_11_15.decap_12
flabel metal1 20157 18143 20191 18177 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_11_Left_39.VPWR
flabel metal1 20157 18687 20191 18721 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_11_Left_39.VGND
flabel nwell 20157 18143 20191 18177 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_11_Left_39.VPB
flabel pwell 20157 18687 20191 18721 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_11_Left_39.VNB
rlabel comment 20220 18704 20220 18704 8 sr_0.PHY_EDGE_ROW_11_Left_39.decap_3
rlabel metal1 19944 18656 20220 18752 5 sr_0.PHY_EDGE_ROW_11_Left_39.VGND
rlabel metal1 19944 18112 20220 18208 5 sr_0.PHY_EDGE_ROW_11_Left_39.VPWR
flabel metal1 17673 18687 17707 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_27.VGND
flabel metal1 17673 18143 17707 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_27.VPWR
flabel nwell 17673 18143 17707 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_27.VPB
flabel pwell 17673 18687 17707 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_27.VNB
rlabel comment 17736 18704 17736 18704 8 sr_0.FILLER_0_11_27.decap_12
flabel metal1 16569 18687 16603 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_39.VGND
flabel metal1 16569 18143 16603 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_39.VPWR
flabel nwell 16569 18143 16603 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_39.VPB
flabel pwell 16569 18687 16603 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_39.VNB
rlabel comment 16632 18704 16632 18704 8 sr_0.FILLER_0_11_39.decap_12
flabel metal1 15465 18687 15499 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_51.VGND
flabel metal1 15465 18143 15499 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_51.VPWR
flabel nwell 15465 18143 15499 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_51.VPB
flabel pwell 15465 18687 15499 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_51.VNB
rlabel comment 15528 18704 15528 18704 8 sr_0.FILLER_0_11_51.decap_4
rlabel metal1 15160 18656 15528 18752 5 sr_0.FILLER_0_11_51.VGND
rlabel metal1 15160 18112 15528 18208 5 sr_0.FILLER_0_11_51.VPWR
flabel metal1 15102 18147 15138 18177 0 FreeSans 250 0 0 0 sr_0.FILLER_0_11_55.VPWR
flabel metal1 15102 18688 15138 18717 0 FreeSans 250 0 0 0 sr_0.FILLER_0_11_55.VGND
flabel nwell 15109 18153 15129 18170 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_55.VPB
flabel pwell 15108 18693 15132 18715 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_55.VNB
rlabel comment 15160 18704 15160 18704 8 sr_0.FILLER_0_11_55.fill_1
rlabel metal1 15068 18656 15160 18752 5 sr_0.FILLER_0_11_55.VGND
rlabel metal1 15068 18112 15160 18208 5 sr_0.FILLER_0_11_55.VPWR
flabel metal1 14913 18687 14947 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_57.VGND
flabel metal1 14913 18143 14947 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_57.VPWR
flabel nwell 14913 18143 14947 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_57.VPB
flabel pwell 14913 18687 14947 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_57.VNB
rlabel comment 14976 18704 14976 18704 8 sr_0.FILLER_0_11_57.decap_12
flabel metal1 14993 18151 15046 18180 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_11_86.VPWR
flabel metal1 14996 18684 15047 18722 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_11_86.VGND
rlabel comment 15068 18704 15068 18704 8 sr_0.TAP_TAPCELL_ROW_11_86.tapvpwrvgnd_1
rlabel metal1 14976 18656 15068 18752 5 sr_0.TAP_TAPCELL_ROW_11_86.VGND
rlabel metal1 14976 18112 15068 18208 5 sr_0.TAP_TAPCELL_ROW_11_86.VPWR
flabel metal1 13809 18687 13843 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_69.VGND
flabel metal1 13809 18143 13843 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_69.VPWR
flabel nwell 13809 18143 13843 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_69.VPB
flabel pwell 13809 18687 13843 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_69.VNB
rlabel comment 13872 18704 13872 18704 8 sr_0.FILLER_0_11_69.decap_12
flabel metal1 12705 18687 12739 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_81.VGND
flabel metal1 12705 18143 12739 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_81.VPWR
flabel nwell 12705 18143 12739 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_81.VPB
flabel pwell 12705 18687 12739 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_81.VNB
rlabel comment 12768 18704 12768 18704 8 sr_0.FILLER_0_11_81.decap_12
flabel metal1 11601 18687 11635 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_93.VGND
flabel metal1 11601 18143 11635 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_93.VPWR
flabel nwell 11601 18143 11635 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_93.VPB
flabel pwell 11601 18687 11635 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_93.VNB
rlabel comment 11664 18704 11664 18704 8 sr_0.FILLER_0_11_93.decap_12
flabel metal1 10497 18143 10531 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_105.VPWR
flabel metal1 10497 18687 10531 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_105.VGND
flabel nwell 10497 18143 10531 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_105.VPB
flabel pwell 10497 18687 10531 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_105.VNB
rlabel comment 10560 18704 10560 18704 8 sr_0.FILLER_0_11_105.decap_6
rlabel metal1 10008 18656 10560 18752 5 sr_0.FILLER_0_11_105.VGND
rlabel metal1 10008 18112 10560 18208 5 sr_0.FILLER_0_11_105.VPWR
flabel metal1 9950 18147 9986 18177 0 FreeSans 250 0 0 0 sr_0.FILLER_0_11_111.VPWR
flabel metal1 9950 18688 9986 18717 0 FreeSans 250 0 0 0 sr_0.FILLER_0_11_111.VGND
flabel nwell 9957 18153 9977 18170 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_111.VPB
flabel pwell 9956 18693 9980 18715 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_111.VNB
rlabel comment 10008 18704 10008 18704 8 sr_0.FILLER_0_11_111.fill_1
rlabel metal1 9916 18656 10008 18752 5 sr_0.FILLER_0_11_111.VGND
rlabel metal1 9916 18112 10008 18208 5 sr_0.FILLER_0_11_111.VPWR
flabel metal1 9761 18687 9795 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_113.VGND
flabel metal1 9761 18143 9795 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_113.VPWR
flabel nwell 9761 18143 9795 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_113.VPB
flabel pwell 9761 18687 9795 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_113.VNB
rlabel comment 9824 18704 9824 18704 8 sr_0.FILLER_0_11_113.decap_12
flabel metal1 8657 18687 8691 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_125.VGND
flabel metal1 8657 18143 8691 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_125.VPWR
flabel nwell 8657 18143 8691 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_125.VPB
flabel pwell 8657 18687 8691 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_125.VNB
rlabel comment 8720 18704 8720 18704 8 sr_0.FILLER_0_11_125.decap_12
flabel metal1 9841 18151 9894 18180 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_11_87.VPWR
flabel metal1 9844 18684 9895 18722 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_11_87.VGND
rlabel comment 9916 18704 9916 18704 8 sr_0.TAP_TAPCELL_ROW_11_87.tapvpwrvgnd_1
rlabel metal1 9824 18656 9916 18752 5 sr_0.TAP_TAPCELL_ROW_11_87.VGND
rlabel metal1 9824 18112 9916 18208 5 sr_0.TAP_TAPCELL_ROW_11_87.VPWR
flabel metal1 7553 18687 7587 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_137.VGND
flabel metal1 7553 18143 7587 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_137.VPWR
flabel nwell 7553 18143 7587 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_137.VPB
flabel pwell 7553 18687 7587 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_137.VNB
rlabel comment 7616 18704 7616 18704 8 sr_0.FILLER_0_11_137.decap_12
flabel metal1 6449 18687 6483 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_149.VGND
flabel metal1 6449 18143 6483 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_149.VPWR
flabel nwell 6449 18143 6483 18177 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_149.VPB
flabel pwell 6449 18687 6483 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_149.VNB
rlabel comment 6512 18704 6512 18704 8 sr_0.FILLER_0_11_149.decap_12
flabel metal1 5335 18686 5388 18718 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_161.VGND
flabel metal1 5335 18143 5387 18174 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_161.VPWR
flabel nwell 5346 18151 5380 18169 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_161.VPB
flabel pwell 5345 18692 5377 18714 0 FreeSans 200 0 0 0 sr_0.FILLER_0_11_161.VNB
rlabel comment 5408 18704 5408 18704 8 sr_0.FILLER_0_11_161.fill_2
rlabel metal1 5224 18656 5408 18752 5 sr_0.FILLER_0_11_161.VGND
rlabel metal1 5224 18112 5408 18208 5 sr_0.FILLER_0_11_161.VPWR
flabel metal1 4977 18143 5011 18177 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_11_Right_11.VPWR
flabel metal1 4977 18687 5011 18721 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_11_Right_11.VGND
flabel nwell 4977 18143 5011 18177 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_11_Right_11.VPB
flabel pwell 4977 18687 5011 18721 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_11_Right_11.VNB
rlabel comment 4948 18704 4948 18704 2 sr_0.PHY_EDGE_ROW_11_Right_11.decap_3
rlabel metal1 4948 18656 5224 18752 5 sr_0.PHY_EDGE_ROW_11_Right_11.VGND
rlabel metal1 4948 18112 5224 18208 5 sr_0.PHY_EDGE_ROW_11_Right_11.VPWR
flabel metal1 19881 18687 19915 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_3.VGND
flabel metal1 19881 19231 19915 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_3.VPWR
flabel nwell 19881 19231 19915 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_3.VPB
flabel pwell 19881 18687 19915 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_3.VNB
rlabel comment 19944 18704 19944 18704 6 sr_0.FILLER_0_12_3.decap_12
flabel metal1 18777 18687 18811 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_15.VGND
flabel metal1 18777 19231 18811 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_15.VPWR
flabel nwell 18777 19231 18811 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_15.VPB
flabel pwell 18777 18687 18811 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_15.VNB
rlabel comment 18840 18704 18840 18704 6 sr_0.FILLER_0_12_15.decap_12
flabel metal1 20157 19231 20191 19265 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_12_Left_40.VPWR
flabel metal1 20157 18687 20191 18721 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_12_Left_40.VGND
flabel nwell 20157 19231 20191 19265 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_12_Left_40.VPB
flabel pwell 20157 18687 20191 18721 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_12_Left_40.VNB
rlabel comment 20220 18704 20220 18704 6 sr_0.PHY_EDGE_ROW_12_Left_40.decap_3
rlabel metal1 19944 18656 20220 18752 1 sr_0.PHY_EDGE_ROW_12_Left_40.VGND
rlabel metal1 19944 19200 20220 19296 1 sr_0.PHY_EDGE_ROW_12_Left_40.VPWR
flabel metal1 17678 19231 17714 19261 0 FreeSans 250 0 0 0 sr_0.FILLER_0_12_27.VPWR
flabel metal1 17678 18691 17714 18720 0 FreeSans 250 0 0 0 sr_0.FILLER_0_12_27.VGND
flabel nwell 17685 19238 17705 19255 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_27.VPB
flabel pwell 17684 18693 17708 18715 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_27.VNB
rlabel comment 17736 18704 17736 18704 6 sr_0.FILLER_0_12_27.fill_1
rlabel metal1 17644 18656 17736 18752 1 sr_0.FILLER_0_12_27.VGND
rlabel metal1 17644 19200 17736 19296 1 sr_0.FILLER_0_12_27.VPWR
flabel metal1 17489 18687 17523 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_29.VGND
flabel metal1 17489 19231 17523 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_29.VPWR
flabel nwell 17489 19231 17523 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_29.VPB
flabel pwell 17489 18687 17523 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_29.VNB
rlabel comment 17552 18704 17552 18704 6 sr_0.FILLER_0_12_29.decap_12
flabel metal1 16385 18687 16419 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_41.VGND
flabel metal1 16385 19231 16419 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_41.VPWR
flabel nwell 16385 19231 16419 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_41.VPB
flabel pwell 16385 18687 16419 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_41.VNB
rlabel comment 16448 18704 16448 18704 6 sr_0.FILLER_0_12_41.decap_12
flabel metal1 17569 19228 17622 19257 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_12_88.VPWR
flabel metal1 17572 18686 17623 18724 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_12_88.VGND
rlabel comment 17644 18704 17644 18704 6 sr_0.TAP_TAPCELL_ROW_12_88.tapvpwrvgnd_1
rlabel metal1 17552 18656 17644 18752 1 sr_0.TAP_TAPCELL_ROW_12_88.VGND
rlabel metal1 17552 19200 17644 19296 1 sr_0.TAP_TAPCELL_ROW_12_88.VPWR
flabel metal1 15281 18687 15315 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_53.VGND
flabel metal1 15281 19231 15315 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_53.VPWR
flabel nwell 15281 19231 15315 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_53.VPB
flabel pwell 15281 18687 15315 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_53.VNB
rlabel comment 15344 18704 15344 18704 6 sr_0.FILLER_0_12_53.decap_12
flabel metal1 14177 18687 14211 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_65.VGND
flabel metal1 14177 19231 14211 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_65.VPWR
flabel nwell 14177 19231 14211 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_65.VPB
flabel pwell 14177 18687 14211 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_65.VNB
rlabel comment 14240 18704 14240 18704 6 sr_0.FILLER_0_12_65.decap_12
flabel metal1 13073 19231 13107 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_77.VPWR
flabel metal1 13073 18687 13107 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_77.VGND
flabel nwell 13073 19231 13107 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_77.VPB
flabel pwell 13073 18687 13107 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_77.VNB
rlabel comment 13136 18704 13136 18704 6 sr_0.FILLER_0_12_77.decap_6
rlabel metal1 12584 18656 13136 18752 1 sr_0.FILLER_0_12_77.VGND
rlabel metal1 12584 19200 13136 19296 1 sr_0.FILLER_0_12_77.VPWR
flabel metal1 12526 19231 12562 19261 0 FreeSans 250 0 0 0 sr_0.FILLER_0_12_83.VPWR
flabel metal1 12526 18691 12562 18720 0 FreeSans 250 0 0 0 sr_0.FILLER_0_12_83.VGND
flabel nwell 12533 19238 12553 19255 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_83.VPB
flabel pwell 12532 18693 12556 18715 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_83.VNB
rlabel comment 12584 18704 12584 18704 6 sr_0.FILLER_0_12_83.fill_1
rlabel metal1 12492 18656 12584 18752 1 sr_0.FILLER_0_12_83.VGND
rlabel metal1 12492 19200 12584 19296 1 sr_0.FILLER_0_12_83.VPWR
flabel metal1 12337 18687 12371 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_85.VGND
flabel metal1 12337 19231 12371 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_85.VPWR
flabel nwell 12337 19231 12371 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_85.VPB
flabel pwell 12337 18687 12371 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_85.VNB
rlabel comment 12400 18704 12400 18704 6 sr_0.FILLER_0_12_85.decap_12
flabel metal1 11233 18687 11267 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_97.VGND
flabel metal1 11233 19231 11267 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_97.VPWR
flabel nwell 11233 19231 11267 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_97.VPB
flabel pwell 11233 18687 11267 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_97.VNB
rlabel comment 11296 18704 11296 18704 6 sr_0.FILLER_0_12_97.decap_12
flabel metal1 12417 19228 12470 19257 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_12_89.VPWR
flabel metal1 12420 18686 12471 18724 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_12_89.VGND
rlabel comment 12492 18704 12492 18704 6 sr_0.TAP_TAPCELL_ROW_12_89.tapvpwrvgnd_1
rlabel metal1 12400 18656 12492 18752 1 sr_0.TAP_TAPCELL_ROW_12_89.VGND
rlabel metal1 12400 19200 12492 19296 1 sr_0.TAP_TAPCELL_ROW_12_89.VPWR
flabel metal1 10129 18687 10163 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_109.VGND
flabel metal1 10129 19231 10163 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_109.VPWR
flabel nwell 10129 19231 10163 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_109.VPB
flabel pwell 10129 18687 10163 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_109.VNB
rlabel comment 10192 18704 10192 18704 6 sr_0.FILLER_0_12_109.decap_12
flabel metal1 9025 18687 9059 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_121.VGND
flabel metal1 9025 19231 9059 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_121.VPWR
flabel nwell 9025 19231 9059 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_121.VPB
flabel pwell 9025 18687 9059 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_121.VNB
rlabel comment 9088 18704 9088 18704 6 sr_0.FILLER_0_12_121.decap_12
flabel metal1 7921 19231 7955 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_133.VPWR
flabel metal1 7921 18687 7955 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_133.VGND
flabel nwell 7921 19231 7955 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_133.VPB
flabel pwell 7921 18687 7955 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_133.VNB
rlabel comment 7984 18704 7984 18704 6 sr_0.FILLER_0_12_133.decap_6
rlabel metal1 7432 18656 7984 18752 1 sr_0.FILLER_0_12_133.VGND
rlabel metal1 7432 19200 7984 19296 1 sr_0.FILLER_0_12_133.VPWR
flabel metal1 7374 19231 7410 19261 0 FreeSans 250 0 0 0 sr_0.FILLER_0_12_139.VPWR
flabel metal1 7374 18691 7410 18720 0 FreeSans 250 0 0 0 sr_0.FILLER_0_12_139.VGND
flabel nwell 7381 19238 7401 19255 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_139.VPB
flabel pwell 7380 18693 7404 18715 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_139.VNB
rlabel comment 7432 18704 7432 18704 6 sr_0.FILLER_0_12_139.fill_1
rlabel metal1 7340 18656 7432 18752 1 sr_0.FILLER_0_12_139.VGND
rlabel metal1 7340 19200 7432 19296 1 sr_0.FILLER_0_12_139.VPWR
flabel metal1 7185 18687 7219 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_141.VGND
flabel metal1 7185 19231 7219 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_141.VPWR
flabel nwell 7185 19231 7219 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_141.VPB
flabel pwell 7185 18687 7219 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_141.VNB
rlabel comment 7248 18704 7248 18704 6 sr_0.FILLER_0_12_141.decap_12
flabel metal1 7265 19228 7318 19257 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_12_90.VPWR
flabel metal1 7268 18686 7319 18724 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_12_90.VGND
rlabel comment 7340 18704 7340 18704 6 sr_0.TAP_TAPCELL_ROW_12_90.tapvpwrvgnd_1
rlabel metal1 7248 18656 7340 18752 1 sr_0.TAP_TAPCELL_ROW_12_90.VGND
rlabel metal1 7248 19200 7340 19296 1 sr_0.TAP_TAPCELL_ROW_12_90.VPWR
flabel metal1 6081 19231 6115 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_153.VPWR
flabel metal1 6081 18687 6115 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_153.VGND
flabel nwell 6081 19231 6115 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_153.VPB
flabel pwell 6081 18687 6115 18721 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_153.VNB
rlabel comment 6144 18704 6144 18704 6 sr_0.FILLER_0_12_153.decap_8
rlabel metal1 5408 18656 6144 18752 1 sr_0.FILLER_0_12_153.VGND
rlabel metal1 5408 19200 6144 19296 1 sr_0.FILLER_0_12_153.VPWR
flabel metal1 5335 18690 5388 18722 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_161.VGND
flabel metal1 5335 19234 5387 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_161.VPWR
flabel nwell 5346 19239 5380 19257 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_161.VPB
flabel pwell 5345 18694 5377 18716 0 FreeSans 200 0 0 0 sr_0.FILLER_0_12_161.VNB
rlabel comment 5408 18704 5408 18704 6 sr_0.FILLER_0_12_161.fill_2
rlabel metal1 5224 18656 5408 18752 1 sr_0.FILLER_0_12_161.VGND
rlabel metal1 5224 19200 5408 19296 1 sr_0.FILLER_0_12_161.VPWR
flabel metal1 4977 19231 5011 19265 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_12_Right_12.VPWR
flabel metal1 4977 18687 5011 18721 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_12_Right_12.VGND
flabel nwell 4977 19231 5011 19265 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_12_Right_12.VPB
flabel pwell 4977 18687 5011 18721 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_12_Right_12.VNB
rlabel comment 4948 18704 4948 18704 4 sr_0.PHY_EDGE_ROW_12_Right_12.decap_3
rlabel metal1 4948 18656 5224 18752 1 sr_0.PHY_EDGE_ROW_12_Right_12.VGND
rlabel metal1 4948 19200 5224 19296 1 sr_0.PHY_EDGE_ROW_12_Right_12.VPWR
flabel metal1 19881 19775 19915 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_3.VGND
flabel metal1 19881 19231 19915 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_3.VPWR
flabel nwell 19881 19231 19915 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_3.VPB
flabel pwell 19881 19775 19915 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_3.VNB
rlabel comment 19944 19792 19944 19792 8 sr_0.FILLER_0_13_3.decap_12
flabel metal1 18777 19775 18811 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_15.VGND
flabel metal1 18777 19231 18811 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_15.VPWR
flabel nwell 18777 19231 18811 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_15.VPB
flabel pwell 18777 19775 18811 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_15.VNB
rlabel comment 18840 19792 18840 19792 8 sr_0.FILLER_0_13_15.decap_12
flabel metal1 19881 19775 19915 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_3.VGND
flabel metal1 19881 20319 19915 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_3.VPWR
flabel nwell 19881 20319 19915 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_3.VPB
flabel pwell 19881 19775 19915 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_3.VNB
rlabel comment 19944 19792 19944 19792 6 sr_0.FILLER_0_14_3.decap_12
flabel metal1 18777 19775 18811 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_15.VGND
flabel metal1 18777 20319 18811 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_15.VPWR
flabel nwell 18777 20319 18811 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_15.VPB
flabel pwell 18777 19775 18811 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_15.VNB
rlabel comment 18840 19792 18840 19792 6 sr_0.FILLER_0_14_15.decap_12
flabel metal1 20157 19231 20191 19265 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_13_Left_41.VPWR
flabel metal1 20157 19775 20191 19809 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_13_Left_41.VGND
flabel nwell 20157 19231 20191 19265 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_13_Left_41.VPB
flabel pwell 20157 19775 20191 19809 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_13_Left_41.VNB
rlabel comment 20220 19792 20220 19792 8 sr_0.PHY_EDGE_ROW_13_Left_41.decap_3
rlabel metal1 19944 19744 20220 19840 5 sr_0.PHY_EDGE_ROW_13_Left_41.VGND
rlabel metal1 19944 19200 20220 19296 5 sr_0.PHY_EDGE_ROW_13_Left_41.VPWR
flabel metal1 20157 20319 20191 20353 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_14_Left_42.VPWR
flabel metal1 20157 19775 20191 19809 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_14_Left_42.VGND
flabel nwell 20157 20319 20191 20353 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_14_Left_42.VPB
flabel pwell 20157 19775 20191 19809 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_14_Left_42.VNB
rlabel comment 20220 19792 20220 19792 6 sr_0.PHY_EDGE_ROW_14_Left_42.decap_3
rlabel metal1 19944 19744 20220 19840 1 sr_0.PHY_EDGE_ROW_14_Left_42.VGND
rlabel metal1 19944 20288 20220 20384 1 sr_0.PHY_EDGE_ROW_14_Left_42.VPWR
flabel metal1 17673 19775 17707 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_27.VGND
flabel metal1 17673 19231 17707 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_27.VPWR
flabel nwell 17673 19231 17707 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_27.VPB
flabel pwell 17673 19775 17707 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_27.VNB
rlabel comment 17736 19792 17736 19792 8 sr_0.FILLER_0_13_27.decap_12
flabel metal1 16569 19775 16603 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_39.VGND
flabel metal1 16569 19231 16603 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_39.VPWR
flabel nwell 16569 19231 16603 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_39.VPB
flabel pwell 16569 19775 16603 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_39.VNB
rlabel comment 16632 19792 16632 19792 8 sr_0.FILLER_0_13_39.decap_12
flabel metal1 17678 20319 17714 20349 0 FreeSans 250 0 0 0 sr_0.FILLER_0_14_27.VPWR
flabel metal1 17678 19779 17714 19808 0 FreeSans 250 0 0 0 sr_0.FILLER_0_14_27.VGND
flabel nwell 17685 20326 17705 20343 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_27.VPB
flabel pwell 17684 19781 17708 19803 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_27.VNB
rlabel comment 17736 19792 17736 19792 6 sr_0.FILLER_0_14_27.fill_1
rlabel metal1 17644 19744 17736 19840 1 sr_0.FILLER_0_14_27.VGND
rlabel metal1 17644 20288 17736 20384 1 sr_0.FILLER_0_14_27.VPWR
flabel metal1 17489 19775 17523 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_29.VGND
flabel metal1 17489 20319 17523 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_29.VPWR
flabel nwell 17489 20319 17523 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_29.VPB
flabel pwell 17489 19775 17523 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_29.VNB
rlabel comment 17552 19792 17552 19792 6 sr_0.FILLER_0_14_29.decap_12
flabel metal1 16385 19775 16419 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_41.VGND
flabel metal1 16385 20319 16419 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_41.VPWR
flabel nwell 16385 20319 16419 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_41.VPB
flabel pwell 16385 19775 16419 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_41.VNB
rlabel comment 16448 19792 16448 19792 6 sr_0.FILLER_0_14_41.decap_12
flabel metal1 17569 20316 17622 20345 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_14_93.VPWR
flabel metal1 17572 19774 17623 19812 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_14_93.VGND
rlabel comment 17644 19792 17644 19792 6 sr_0.TAP_TAPCELL_ROW_14_93.tapvpwrvgnd_1
rlabel metal1 17552 19744 17644 19840 1 sr_0.TAP_TAPCELL_ROW_14_93.VGND
rlabel metal1 17552 20288 17644 20384 1 sr_0.TAP_TAPCELL_ROW_14_93.VPWR
flabel metal1 15465 19775 15499 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_51.VGND
flabel metal1 15465 19231 15499 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_51.VPWR
flabel nwell 15465 19231 15499 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_51.VPB
flabel pwell 15465 19775 15499 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_51.VNB
rlabel comment 15528 19792 15528 19792 8 sr_0.FILLER_0_13_51.decap_4
rlabel metal1 15160 19744 15528 19840 5 sr_0.FILLER_0_13_51.VGND
rlabel metal1 15160 19200 15528 19296 5 sr_0.FILLER_0_13_51.VPWR
flabel metal1 15102 19235 15138 19265 0 FreeSans 250 0 0 0 sr_0.FILLER_0_13_55.VPWR
flabel metal1 15102 19776 15138 19805 0 FreeSans 250 0 0 0 sr_0.FILLER_0_13_55.VGND
flabel nwell 15109 19241 15129 19258 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_55.VPB
flabel pwell 15108 19781 15132 19803 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_55.VNB
rlabel comment 15160 19792 15160 19792 8 sr_0.FILLER_0_13_55.fill_1
rlabel metal1 15068 19744 15160 19840 5 sr_0.FILLER_0_13_55.VGND
rlabel metal1 15068 19200 15160 19296 5 sr_0.FILLER_0_13_55.VPWR
flabel metal1 14913 19775 14947 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_57.VGND
flabel metal1 14913 19231 14947 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_57.VPWR
flabel nwell 14913 19231 14947 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_57.VPB
flabel pwell 14913 19775 14947 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_57.VNB
rlabel comment 14976 19792 14976 19792 8 sr_0.FILLER_0_13_57.decap_12
flabel metal1 15281 19775 15315 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_53.VGND
flabel metal1 15281 20319 15315 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_53.VPWR
flabel nwell 15281 20319 15315 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_53.VPB
flabel pwell 15281 19775 15315 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_53.VNB
rlabel comment 15344 19792 15344 19792 6 sr_0.FILLER_0_14_53.decap_12
flabel metal1 14993 19239 15046 19268 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_13_91.VPWR
flabel metal1 14996 19772 15047 19810 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_13_91.VGND
rlabel comment 15068 19792 15068 19792 8 sr_0.TAP_TAPCELL_ROW_13_91.tapvpwrvgnd_1
rlabel metal1 14976 19744 15068 19840 5 sr_0.TAP_TAPCELL_ROW_13_91.VGND
rlabel metal1 14976 19200 15068 19296 5 sr_0.TAP_TAPCELL_ROW_13_91.VPWR
flabel metal1 13809 19775 13843 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_69.VGND
flabel metal1 13809 19231 13843 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_69.VPWR
flabel nwell 13809 19231 13843 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_69.VPB
flabel pwell 13809 19775 13843 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_69.VNB
rlabel comment 13872 19792 13872 19792 8 sr_0.FILLER_0_13_69.decap_12
flabel metal1 12705 19775 12739 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_81.VGND
flabel metal1 12705 19231 12739 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_81.VPWR
flabel nwell 12705 19231 12739 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_81.VPB
flabel pwell 12705 19775 12739 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_81.VNB
rlabel comment 12768 19792 12768 19792 8 sr_0.FILLER_0_13_81.decap_12
flabel metal1 14177 19775 14211 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_65.VGND
flabel metal1 14177 20319 14211 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_65.VPWR
flabel nwell 14177 20319 14211 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_65.VPB
flabel pwell 14177 19775 14211 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_65.VNB
rlabel comment 14240 19792 14240 19792 6 sr_0.FILLER_0_14_65.decap_12
flabel metal1 13073 20319 13107 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_77.VPWR
flabel metal1 13073 19775 13107 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_77.VGND
flabel nwell 13073 20319 13107 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_77.VPB
flabel pwell 13073 19775 13107 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_77.VNB
rlabel comment 13136 19792 13136 19792 6 sr_0.FILLER_0_14_77.decap_6
rlabel metal1 12584 19744 13136 19840 1 sr_0.FILLER_0_14_77.VGND
rlabel metal1 12584 20288 13136 20384 1 sr_0.FILLER_0_14_77.VPWR
flabel metal1 12526 20319 12562 20349 0 FreeSans 250 0 0 0 sr_0.FILLER_0_14_83.VPWR
flabel metal1 12526 19779 12562 19808 0 FreeSans 250 0 0 0 sr_0.FILLER_0_14_83.VGND
flabel nwell 12533 20326 12553 20343 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_83.VPB
flabel pwell 12532 19781 12556 19803 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_83.VNB
rlabel comment 12584 19792 12584 19792 6 sr_0.FILLER_0_14_83.fill_1
rlabel metal1 12492 19744 12584 19840 1 sr_0.FILLER_0_14_83.VGND
rlabel metal1 12492 20288 12584 20384 1 sr_0.FILLER_0_14_83.VPWR
flabel metal1 11601 19775 11635 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_93.VGND
flabel metal1 11601 19231 11635 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_93.VPWR
flabel nwell 11601 19231 11635 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_93.VPB
flabel pwell 11601 19775 11635 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_93.VNB
rlabel comment 11664 19792 11664 19792 8 sr_0.FILLER_0_13_93.decap_12
flabel metal1 12337 19775 12371 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_85.VGND
flabel metal1 12337 20319 12371 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_85.VPWR
flabel nwell 12337 20319 12371 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_85.VPB
flabel pwell 12337 19775 12371 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_85.VNB
rlabel comment 12400 19792 12400 19792 6 sr_0.FILLER_0_14_85.decap_12
flabel metal1 11233 19775 11267 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_97.VGND
flabel metal1 11233 20319 11267 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_97.VPWR
flabel nwell 11233 20319 11267 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_97.VPB
flabel pwell 11233 19775 11267 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_97.VNB
rlabel comment 11296 19792 11296 19792 6 sr_0.FILLER_0_14_97.decap_12
flabel metal1 12417 20316 12470 20345 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_14_94.VPWR
flabel metal1 12420 19774 12471 19812 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_14_94.VGND
rlabel comment 12492 19792 12492 19792 6 sr_0.TAP_TAPCELL_ROW_14_94.tapvpwrvgnd_1
rlabel metal1 12400 19744 12492 19840 1 sr_0.TAP_TAPCELL_ROW_14_94.VGND
rlabel metal1 12400 20288 12492 20384 1 sr_0.TAP_TAPCELL_ROW_14_94.VPWR
flabel metal1 10497 19231 10531 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_105.VPWR
flabel metal1 10497 19775 10531 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_105.VGND
flabel nwell 10497 19231 10531 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_105.VPB
flabel pwell 10497 19775 10531 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_105.VNB
rlabel comment 10560 19792 10560 19792 8 sr_0.FILLER_0_13_105.decap_6
rlabel metal1 10008 19744 10560 19840 5 sr_0.FILLER_0_13_105.VGND
rlabel metal1 10008 19200 10560 19296 5 sr_0.FILLER_0_13_105.VPWR
flabel metal1 9950 19235 9986 19265 0 FreeSans 250 0 0 0 sr_0.FILLER_0_13_111.VPWR
flabel metal1 9950 19776 9986 19805 0 FreeSans 250 0 0 0 sr_0.FILLER_0_13_111.VGND
flabel nwell 9957 19241 9977 19258 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_111.VPB
flabel pwell 9956 19781 9980 19803 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_111.VNB
rlabel comment 10008 19792 10008 19792 8 sr_0.FILLER_0_13_111.fill_1
rlabel metal1 9916 19744 10008 19840 5 sr_0.FILLER_0_13_111.VGND
rlabel metal1 9916 19200 10008 19296 5 sr_0.FILLER_0_13_111.VPWR
flabel metal1 9761 19775 9795 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_113.VGND
flabel metal1 9761 19231 9795 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_113.VPWR
flabel nwell 9761 19231 9795 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_113.VPB
flabel pwell 9761 19775 9795 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_113.VNB
rlabel comment 9824 19792 9824 19792 8 sr_0.FILLER_0_13_113.decap_12
flabel metal1 8657 19775 8691 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_125.VGND
flabel metal1 8657 19231 8691 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_125.VPWR
flabel nwell 8657 19231 8691 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_125.VPB
flabel pwell 8657 19775 8691 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_125.VNB
rlabel comment 8720 19792 8720 19792 8 sr_0.FILLER_0_13_125.decap_12
flabel metal1 10129 19775 10163 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_109.VGND
flabel metal1 10129 20319 10163 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_109.VPWR
flabel nwell 10129 20319 10163 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_109.VPB
flabel pwell 10129 19775 10163 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_109.VNB
rlabel comment 10192 19792 10192 19792 6 sr_0.FILLER_0_14_109.decap_12
flabel metal1 9025 19775 9059 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_121.VGND
flabel metal1 9025 20319 9059 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_121.VPWR
flabel nwell 9025 20319 9059 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_121.VPB
flabel pwell 9025 19775 9059 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_121.VNB
rlabel comment 9088 19792 9088 19792 6 sr_0.FILLER_0_14_121.decap_12
flabel metal1 9841 19239 9894 19268 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_13_92.VPWR
flabel metal1 9844 19772 9895 19810 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_13_92.VGND
rlabel comment 9916 19792 9916 19792 8 sr_0.TAP_TAPCELL_ROW_13_92.tapvpwrvgnd_1
rlabel metal1 9824 19744 9916 19840 5 sr_0.TAP_TAPCELL_ROW_13_92.VGND
rlabel metal1 9824 19200 9916 19296 5 sr_0.TAP_TAPCELL_ROW_13_92.VPWR
flabel metal1 7553 19775 7587 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_137.VGND
flabel metal1 7553 19231 7587 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_137.VPWR
flabel nwell 7553 19231 7587 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_137.VPB
flabel pwell 7553 19775 7587 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_137.VNB
rlabel comment 7616 19792 7616 19792 8 sr_0.FILLER_0_13_137.decap_12
flabel metal1 7921 20319 7955 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_133.VPWR
flabel metal1 7921 19775 7955 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_133.VGND
flabel nwell 7921 20319 7955 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_133.VPB
flabel pwell 7921 19775 7955 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_133.VNB
rlabel comment 7984 19792 7984 19792 6 sr_0.FILLER_0_14_133.decap_6
rlabel metal1 7432 19744 7984 19840 1 sr_0.FILLER_0_14_133.VGND
rlabel metal1 7432 20288 7984 20384 1 sr_0.FILLER_0_14_133.VPWR
flabel metal1 7374 20319 7410 20349 0 FreeSans 250 0 0 0 sr_0.FILLER_0_14_139.VPWR
flabel metal1 7374 19779 7410 19808 0 FreeSans 250 0 0 0 sr_0.FILLER_0_14_139.VGND
flabel nwell 7381 20326 7401 20343 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_139.VPB
flabel pwell 7380 19781 7404 19803 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_139.VNB
rlabel comment 7432 19792 7432 19792 6 sr_0.FILLER_0_14_139.fill_1
rlabel metal1 7340 19744 7432 19840 1 sr_0.FILLER_0_14_139.VGND
rlabel metal1 7340 20288 7432 20384 1 sr_0.FILLER_0_14_139.VPWR
flabel metal1 7185 19775 7219 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_141.VGND
flabel metal1 7185 20319 7219 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_141.VPWR
flabel nwell 7185 20319 7219 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_141.VPB
flabel pwell 7185 19775 7219 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_141.VNB
rlabel comment 7248 19792 7248 19792 6 sr_0.FILLER_0_14_141.decap_12
flabel metal1 7265 20316 7318 20345 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_14_95.VPWR
flabel metal1 7268 19774 7319 19812 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_14_95.VGND
rlabel comment 7340 19792 7340 19792 6 sr_0.TAP_TAPCELL_ROW_14_95.tapvpwrvgnd_1
rlabel metal1 7248 19744 7340 19840 1 sr_0.TAP_TAPCELL_ROW_14_95.VGND
rlabel metal1 7248 20288 7340 20384 1 sr_0.TAP_TAPCELL_ROW_14_95.VPWR
flabel metal1 6449 19775 6483 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_149.VGND
flabel metal1 6449 19231 6483 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_149.VPWR
flabel nwell 6449 19231 6483 19265 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_149.VPB
flabel pwell 6449 19775 6483 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_149.VNB
rlabel comment 6512 19792 6512 19792 8 sr_0.FILLER_0_13_149.decap_12
flabel metal1 5335 19774 5388 19806 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_161.VGND
flabel metal1 5335 19231 5387 19262 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_161.VPWR
flabel nwell 5346 19239 5380 19257 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_161.VPB
flabel pwell 5345 19780 5377 19802 0 FreeSans 200 0 0 0 sr_0.FILLER_0_13_161.VNB
rlabel comment 5408 19792 5408 19792 8 sr_0.FILLER_0_13_161.fill_2
rlabel metal1 5224 19744 5408 19840 5 sr_0.FILLER_0_13_161.VGND
rlabel metal1 5224 19200 5408 19296 5 sr_0.FILLER_0_13_161.VPWR
flabel metal1 6081 20319 6115 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_153.VPWR
flabel metal1 6081 19775 6115 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_153.VGND
flabel nwell 6081 20319 6115 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_153.VPB
flabel pwell 6081 19775 6115 19809 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_153.VNB
rlabel comment 6144 19792 6144 19792 6 sr_0.FILLER_0_14_153.decap_8
rlabel metal1 5408 19744 6144 19840 1 sr_0.FILLER_0_14_153.VGND
rlabel metal1 5408 20288 6144 20384 1 sr_0.FILLER_0_14_153.VPWR
flabel metal1 5335 19778 5388 19810 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_161.VGND
flabel metal1 5335 20322 5387 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_161.VPWR
flabel nwell 5346 20327 5380 20345 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_161.VPB
flabel pwell 5345 19782 5377 19804 0 FreeSans 200 0 0 0 sr_0.FILLER_0_14_161.VNB
rlabel comment 5408 19792 5408 19792 6 sr_0.FILLER_0_14_161.fill_2
rlabel metal1 5224 19744 5408 19840 1 sr_0.FILLER_0_14_161.VGND
rlabel metal1 5224 20288 5408 20384 1 sr_0.FILLER_0_14_161.VPWR
flabel metal1 4977 19231 5011 19265 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_13_Right_13.VPWR
flabel metal1 4977 19775 5011 19809 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_13_Right_13.VGND
flabel nwell 4977 19231 5011 19265 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_13_Right_13.VPB
flabel pwell 4977 19775 5011 19809 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_13_Right_13.VNB
rlabel comment 4948 19792 4948 19792 2 sr_0.PHY_EDGE_ROW_13_Right_13.decap_3
rlabel metal1 4948 19744 5224 19840 5 sr_0.PHY_EDGE_ROW_13_Right_13.VGND
rlabel metal1 4948 19200 5224 19296 5 sr_0.PHY_EDGE_ROW_13_Right_13.VPWR
flabel metal1 4977 20319 5011 20353 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_14_Right_14.VPWR
flabel metal1 4977 19775 5011 19809 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_14_Right_14.VGND
flabel nwell 4977 20319 5011 20353 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_14_Right_14.VPB
flabel pwell 4977 19775 5011 19809 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_14_Right_14.VNB
rlabel comment 4948 19792 4948 19792 4 sr_0.PHY_EDGE_ROW_14_Right_14.decap_3
rlabel metal1 4948 19744 5224 19840 1 sr_0.PHY_EDGE_ROW_14_Right_14.VGND
rlabel metal1 4948 20288 5224 20384 1 sr_0.PHY_EDGE_ROW_14_Right_14.VPWR
flabel metal1 19881 20863 19915 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_3.VGND
flabel metal1 19881 20319 19915 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_3.VPWR
flabel nwell 19881 20319 19915 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_3.VPB
flabel pwell 19881 20863 19915 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_3.VNB
rlabel comment 19944 20880 19944 20880 8 sr_0.FILLER_0_15_3.decap_12
flabel metal1 18777 20863 18811 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_15.VGND
flabel metal1 18777 20319 18811 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_15.VPWR
flabel nwell 18777 20319 18811 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_15.VPB
flabel pwell 18777 20863 18811 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_15.VNB
rlabel comment 18840 20880 18840 20880 8 sr_0.FILLER_0_15_15.decap_12
flabel metal1 20157 20319 20191 20353 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_15_Left_43.VPWR
flabel metal1 20157 20863 20191 20897 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_15_Left_43.VGND
flabel nwell 20157 20319 20191 20353 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_15_Left_43.VPB
flabel pwell 20157 20863 20191 20897 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_15_Left_43.VNB
rlabel comment 20220 20880 20220 20880 8 sr_0.PHY_EDGE_ROW_15_Left_43.decap_3
rlabel metal1 19944 20832 20220 20928 5 sr_0.PHY_EDGE_ROW_15_Left_43.VGND
rlabel metal1 19944 20288 20220 20384 5 sr_0.PHY_EDGE_ROW_15_Left_43.VPWR
flabel metal1 17673 20863 17707 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_27.VGND
flabel metal1 17673 20319 17707 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_27.VPWR
flabel nwell 17673 20319 17707 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_27.VPB
flabel pwell 17673 20863 17707 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_27.VNB
rlabel comment 17736 20880 17736 20880 8 sr_0.FILLER_0_15_27.decap_12
flabel metal1 16569 20863 16603 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_39.VGND
flabel metal1 16569 20319 16603 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_39.VPWR
flabel nwell 16569 20319 16603 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_39.VPB
flabel pwell 16569 20863 16603 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_39.VNB
rlabel comment 16632 20880 16632 20880 8 sr_0.FILLER_0_15_39.decap_12
flabel metal1 15465 20863 15499 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_51.VGND
flabel metal1 15465 20319 15499 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_51.VPWR
flabel nwell 15465 20319 15499 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_51.VPB
flabel pwell 15465 20863 15499 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_51.VNB
rlabel comment 15528 20880 15528 20880 8 sr_0.FILLER_0_15_51.decap_4
rlabel metal1 15160 20832 15528 20928 5 sr_0.FILLER_0_15_51.VGND
rlabel metal1 15160 20288 15528 20384 5 sr_0.FILLER_0_15_51.VPWR
flabel metal1 15102 20323 15138 20353 0 FreeSans 250 0 0 0 sr_0.FILLER_0_15_55.VPWR
flabel metal1 15102 20864 15138 20893 0 FreeSans 250 0 0 0 sr_0.FILLER_0_15_55.VGND
flabel nwell 15109 20329 15129 20346 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_55.VPB
flabel pwell 15108 20869 15132 20891 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_55.VNB
rlabel comment 15160 20880 15160 20880 8 sr_0.FILLER_0_15_55.fill_1
rlabel metal1 15068 20832 15160 20928 5 sr_0.FILLER_0_15_55.VGND
rlabel metal1 15068 20288 15160 20384 5 sr_0.FILLER_0_15_55.VPWR
flabel metal1 14913 20863 14947 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_57.VGND
flabel metal1 14913 20319 14947 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_57.VPWR
flabel nwell 14913 20319 14947 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_57.VPB
flabel pwell 14913 20863 14947 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_57.VNB
rlabel comment 14976 20880 14976 20880 8 sr_0.FILLER_0_15_57.decap_12
flabel metal1 14993 20327 15046 20356 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_15_96.VPWR
flabel metal1 14996 20860 15047 20898 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_15_96.VGND
rlabel comment 15068 20880 15068 20880 8 sr_0.TAP_TAPCELL_ROW_15_96.tapvpwrvgnd_1
rlabel metal1 14976 20832 15068 20928 5 sr_0.TAP_TAPCELL_ROW_15_96.VGND
rlabel metal1 14976 20288 15068 20384 5 sr_0.TAP_TAPCELL_ROW_15_96.VPWR
flabel metal1 13809 20863 13843 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_69.VGND
flabel metal1 13809 20319 13843 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_69.VPWR
flabel nwell 13809 20319 13843 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_69.VPB
flabel pwell 13809 20863 13843 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_69.VNB
rlabel comment 13872 20880 13872 20880 8 sr_0.FILLER_0_15_69.decap_12
flabel metal1 12705 20863 12739 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_81.VGND
flabel metal1 12705 20319 12739 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_81.VPWR
flabel nwell 12705 20319 12739 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_81.VPB
flabel pwell 12705 20863 12739 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_81.VNB
rlabel comment 12768 20880 12768 20880 8 sr_0.FILLER_0_15_81.decap_12
flabel metal1 11601 20863 11635 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_93.VGND
flabel metal1 11601 20319 11635 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_93.VPWR
flabel nwell 11601 20319 11635 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_93.VPB
flabel pwell 11601 20863 11635 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_93.VNB
rlabel comment 11664 20880 11664 20880 8 sr_0.FILLER_0_15_93.decap_12
flabel metal1 10497 20319 10531 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_105.VPWR
flabel metal1 10497 20863 10531 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_105.VGND
flabel nwell 10497 20319 10531 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_105.VPB
flabel pwell 10497 20863 10531 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_105.VNB
rlabel comment 10560 20880 10560 20880 8 sr_0.FILLER_0_15_105.decap_6
rlabel metal1 10008 20832 10560 20928 5 sr_0.FILLER_0_15_105.VGND
rlabel metal1 10008 20288 10560 20384 5 sr_0.FILLER_0_15_105.VPWR
flabel metal1 9950 20323 9986 20353 0 FreeSans 250 0 0 0 sr_0.FILLER_0_15_111.VPWR
flabel metal1 9950 20864 9986 20893 0 FreeSans 250 0 0 0 sr_0.FILLER_0_15_111.VGND
flabel nwell 9957 20329 9977 20346 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_111.VPB
flabel pwell 9956 20869 9980 20891 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_111.VNB
rlabel comment 10008 20880 10008 20880 8 sr_0.FILLER_0_15_111.fill_1
rlabel metal1 9916 20832 10008 20928 5 sr_0.FILLER_0_15_111.VGND
rlabel metal1 9916 20288 10008 20384 5 sr_0.FILLER_0_15_111.VPWR
flabel metal1 9761 20863 9795 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_113.VGND
flabel metal1 9761 20319 9795 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_113.VPWR
flabel nwell 9761 20319 9795 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_113.VPB
flabel pwell 9761 20863 9795 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_113.VNB
rlabel comment 9824 20880 9824 20880 8 sr_0.FILLER_0_15_113.decap_12
flabel metal1 8657 20863 8691 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_125.VGND
flabel metal1 8657 20319 8691 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_125.VPWR
flabel nwell 8657 20319 8691 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_125.VPB
flabel pwell 8657 20863 8691 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_125.VNB
rlabel comment 8720 20880 8720 20880 8 sr_0.FILLER_0_15_125.decap_12
flabel metal1 9841 20327 9894 20356 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_15_97.VPWR
flabel metal1 9844 20860 9895 20898 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_15_97.VGND
rlabel comment 9916 20880 9916 20880 8 sr_0.TAP_TAPCELL_ROW_15_97.tapvpwrvgnd_1
rlabel metal1 9824 20832 9916 20928 5 sr_0.TAP_TAPCELL_ROW_15_97.VGND
rlabel metal1 9824 20288 9916 20384 5 sr_0.TAP_TAPCELL_ROW_15_97.VPWR
flabel metal1 7553 20863 7587 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_137.VGND
flabel metal1 7553 20319 7587 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_137.VPWR
flabel nwell 7553 20319 7587 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_137.VPB
flabel pwell 7553 20863 7587 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_137.VNB
rlabel comment 7616 20880 7616 20880 8 sr_0.FILLER_0_15_137.decap_12
flabel metal1 6449 20863 6483 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_149.VGND
flabel metal1 6449 20319 6483 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_149.VPWR
flabel nwell 6449 20319 6483 20353 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_149.VPB
flabel pwell 6449 20863 6483 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_149.VNB
rlabel comment 6512 20880 6512 20880 8 sr_0.FILLER_0_15_149.decap_12
flabel metal1 5335 20862 5388 20894 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_161.VGND
flabel metal1 5335 20319 5387 20350 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_161.VPWR
flabel nwell 5346 20327 5380 20345 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_161.VPB
flabel pwell 5345 20868 5377 20890 0 FreeSans 200 0 0 0 sr_0.FILLER_0_15_161.VNB
rlabel comment 5408 20880 5408 20880 8 sr_0.FILLER_0_15_161.fill_2
rlabel metal1 5224 20832 5408 20928 5 sr_0.FILLER_0_15_161.VGND
rlabel metal1 5224 20288 5408 20384 5 sr_0.FILLER_0_15_161.VPWR
flabel metal1 4977 20319 5011 20353 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_15_Right_15.VPWR
flabel metal1 4977 20863 5011 20897 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_15_Right_15.VGND
flabel nwell 4977 20319 5011 20353 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_15_Right_15.VPB
flabel pwell 4977 20863 5011 20897 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_15_Right_15.VNB
rlabel comment 4948 20880 4948 20880 2 sr_0.PHY_EDGE_ROW_15_Right_15.decap_3
rlabel metal1 4948 20832 5224 20928 5 sr_0.PHY_EDGE_ROW_15_Right_15.VGND
rlabel metal1 4948 20288 5224 20384 5 sr_0.PHY_EDGE_ROW_15_Right_15.VPWR
flabel metal1 19881 20863 19915 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_3.VGND
flabel metal1 19881 21407 19915 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_3.VPWR
flabel nwell 19881 21407 19915 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_3.VPB
flabel pwell 19881 20863 19915 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_3.VNB
rlabel comment 19944 20880 19944 20880 6 sr_0.FILLER_0_16_3.decap_12
flabel metal1 18777 20863 18811 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_15.VGND
flabel metal1 18777 21407 18811 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_15.VPWR
flabel nwell 18777 21407 18811 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_15.VPB
flabel pwell 18777 20863 18811 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_15.VNB
rlabel comment 18840 20880 18840 20880 6 sr_0.FILLER_0_16_15.decap_12
flabel metal1 20157 21407 20191 21441 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_16_Left_44.VPWR
flabel metal1 20157 20863 20191 20897 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_16_Left_44.VGND
flabel nwell 20157 21407 20191 21441 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_16_Left_44.VPB
flabel pwell 20157 20863 20191 20897 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_16_Left_44.VNB
rlabel comment 20220 20880 20220 20880 6 sr_0.PHY_EDGE_ROW_16_Left_44.decap_3
rlabel metal1 19944 20832 20220 20928 1 sr_0.PHY_EDGE_ROW_16_Left_44.VGND
rlabel metal1 19944 21376 20220 21472 1 sr_0.PHY_EDGE_ROW_16_Left_44.VPWR
flabel metal1 17678 21407 17714 21437 0 FreeSans 250 0 0 0 sr_0.FILLER_0_16_27.VPWR
flabel metal1 17678 20867 17714 20896 0 FreeSans 250 0 0 0 sr_0.FILLER_0_16_27.VGND
flabel nwell 17685 21414 17705 21431 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_27.VPB
flabel pwell 17684 20869 17708 20891 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_27.VNB
rlabel comment 17736 20880 17736 20880 6 sr_0.FILLER_0_16_27.fill_1
rlabel metal1 17644 20832 17736 20928 1 sr_0.FILLER_0_16_27.VGND
rlabel metal1 17644 21376 17736 21472 1 sr_0.FILLER_0_16_27.VPWR
flabel metal1 17489 20863 17523 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_29.VGND
flabel metal1 17489 21407 17523 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_29.VPWR
flabel nwell 17489 21407 17523 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_29.VPB
flabel pwell 17489 20863 17523 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_29.VNB
rlabel comment 17552 20880 17552 20880 6 sr_0.FILLER_0_16_29.decap_12
flabel metal1 16385 20863 16419 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_41.VGND
flabel metal1 16385 21407 16419 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_41.VPWR
flabel nwell 16385 21407 16419 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_41.VPB
flabel pwell 16385 20863 16419 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_41.VNB
rlabel comment 16448 20880 16448 20880 6 sr_0.FILLER_0_16_41.decap_12
flabel metal1 17569 21404 17622 21433 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_16_98.VPWR
flabel metal1 17572 20862 17623 20900 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_16_98.VGND
rlabel comment 17644 20880 17644 20880 6 sr_0.TAP_TAPCELL_ROW_16_98.tapvpwrvgnd_1
rlabel metal1 17552 20832 17644 20928 1 sr_0.TAP_TAPCELL_ROW_16_98.VGND
rlabel metal1 17552 21376 17644 21472 1 sr_0.TAP_TAPCELL_ROW_16_98.VPWR
flabel metal1 15281 20863 15315 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_53.VGND
flabel metal1 15281 21407 15315 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_53.VPWR
flabel nwell 15281 21407 15315 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_53.VPB
flabel pwell 15281 20863 15315 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_53.VNB
rlabel comment 15344 20880 15344 20880 6 sr_0.FILLER_0_16_53.decap_12
flabel metal1 14177 20863 14211 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_65.VGND
flabel metal1 14177 21407 14211 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_65.VPWR
flabel nwell 14177 21407 14211 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_65.VPB
flabel pwell 14177 20863 14211 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_65.VNB
rlabel comment 14240 20880 14240 20880 6 sr_0.FILLER_0_16_65.decap_12
flabel metal1 13073 21407 13107 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_77.VPWR
flabel metal1 13073 20863 13107 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_77.VGND
flabel nwell 13073 21407 13107 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_77.VPB
flabel pwell 13073 20863 13107 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_77.VNB
rlabel comment 13136 20880 13136 20880 6 sr_0.FILLER_0_16_77.decap_6
rlabel metal1 12584 20832 13136 20928 1 sr_0.FILLER_0_16_77.VGND
rlabel metal1 12584 21376 13136 21472 1 sr_0.FILLER_0_16_77.VPWR
flabel metal1 12526 21407 12562 21437 0 FreeSans 250 0 0 0 sr_0.FILLER_0_16_83.VPWR
flabel metal1 12526 20867 12562 20896 0 FreeSans 250 0 0 0 sr_0.FILLER_0_16_83.VGND
flabel nwell 12533 21414 12553 21431 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_83.VPB
flabel pwell 12532 20869 12556 20891 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_83.VNB
rlabel comment 12584 20880 12584 20880 6 sr_0.FILLER_0_16_83.fill_1
rlabel metal1 12492 20832 12584 20928 1 sr_0.FILLER_0_16_83.VGND
rlabel metal1 12492 21376 12584 21472 1 sr_0.FILLER_0_16_83.VPWR
flabel metal1 12337 20863 12371 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_85.VGND
flabel metal1 12337 21407 12371 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_85.VPWR
flabel nwell 12337 21407 12371 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_85.VPB
flabel pwell 12337 20863 12371 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_85.VNB
rlabel comment 12400 20880 12400 20880 6 sr_0.FILLER_0_16_85.decap_12
flabel metal1 11233 20863 11267 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_97.VGND
flabel metal1 11233 21407 11267 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_97.VPWR
flabel nwell 11233 21407 11267 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_97.VPB
flabel pwell 11233 20863 11267 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_97.VNB
rlabel comment 11296 20880 11296 20880 6 sr_0.FILLER_0_16_97.decap_12
flabel metal1 12417 21404 12470 21433 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_16_99.VPWR
flabel metal1 12420 20862 12471 20900 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_16_99.VGND
rlabel comment 12492 20880 12492 20880 6 sr_0.TAP_TAPCELL_ROW_16_99.tapvpwrvgnd_1
rlabel metal1 12400 20832 12492 20928 1 sr_0.TAP_TAPCELL_ROW_16_99.VGND
rlabel metal1 12400 21376 12492 21472 1 sr_0.TAP_TAPCELL_ROW_16_99.VPWR
flabel metal1 10129 20863 10163 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_109.VGND
flabel metal1 10129 21407 10163 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_109.VPWR
flabel nwell 10129 21407 10163 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_109.VPB
flabel pwell 10129 20863 10163 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_109.VNB
rlabel comment 10192 20880 10192 20880 6 sr_0.FILLER_0_16_109.decap_12
flabel metal1 9025 20863 9059 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_121.VGND
flabel metal1 9025 21407 9059 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_121.VPWR
flabel nwell 9025 21407 9059 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_121.VPB
flabel pwell 9025 20863 9059 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_121.VNB
rlabel comment 9088 20880 9088 20880 6 sr_0.FILLER_0_16_121.decap_12
flabel metal1 7921 21407 7955 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_133.VPWR
flabel metal1 7921 20863 7955 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_133.VGND
flabel nwell 7921 21407 7955 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_133.VPB
flabel pwell 7921 20863 7955 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_133.VNB
rlabel comment 7984 20880 7984 20880 6 sr_0.FILLER_0_16_133.decap_6
rlabel metal1 7432 20832 7984 20928 1 sr_0.FILLER_0_16_133.VGND
rlabel metal1 7432 21376 7984 21472 1 sr_0.FILLER_0_16_133.VPWR
flabel metal1 7374 21407 7410 21437 0 FreeSans 250 0 0 0 sr_0.FILLER_0_16_139.VPWR
flabel metal1 7374 20867 7410 20896 0 FreeSans 250 0 0 0 sr_0.FILLER_0_16_139.VGND
flabel nwell 7381 21414 7401 21431 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_139.VPB
flabel pwell 7380 20869 7404 20891 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_139.VNB
rlabel comment 7432 20880 7432 20880 6 sr_0.FILLER_0_16_139.fill_1
rlabel metal1 7340 20832 7432 20928 1 sr_0.FILLER_0_16_139.VGND
rlabel metal1 7340 21376 7432 21472 1 sr_0.FILLER_0_16_139.VPWR
flabel metal1 7185 20863 7219 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_141.VGND
flabel metal1 7185 21407 7219 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_141.VPWR
flabel nwell 7185 21407 7219 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_141.VPB
flabel pwell 7185 20863 7219 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_141.VNB
rlabel comment 7248 20880 7248 20880 6 sr_0.FILLER_0_16_141.decap_12
flabel metal1 7265 21404 7318 21433 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_16_100.VPWR
flabel metal1 7268 20862 7319 20900 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_16_100.VGND
rlabel comment 7340 20880 7340 20880 6 sr_0.TAP_TAPCELL_ROW_16_100.tapvpwrvgnd_1
rlabel metal1 7248 20832 7340 20928 1 sr_0.TAP_TAPCELL_ROW_16_100.VGND
rlabel metal1 7248 21376 7340 21472 1 sr_0.TAP_TAPCELL_ROW_16_100.VPWR
flabel metal1 6081 21407 6115 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_153.VPWR
flabel metal1 6081 20863 6115 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_153.VGND
flabel nwell 6081 21407 6115 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_153.VPB
flabel pwell 6081 20863 6115 20897 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_153.VNB
rlabel comment 6144 20880 6144 20880 6 sr_0.FILLER_0_16_153.decap_8
rlabel metal1 5408 20832 6144 20928 1 sr_0.FILLER_0_16_153.VGND
rlabel metal1 5408 21376 6144 21472 1 sr_0.FILLER_0_16_153.VPWR
flabel metal1 5335 20866 5388 20898 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_161.VGND
flabel metal1 5335 21410 5387 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_161.VPWR
flabel nwell 5346 21415 5380 21433 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_161.VPB
flabel pwell 5345 20870 5377 20892 0 FreeSans 200 0 0 0 sr_0.FILLER_0_16_161.VNB
rlabel comment 5408 20880 5408 20880 6 sr_0.FILLER_0_16_161.fill_2
rlabel metal1 5224 20832 5408 20928 1 sr_0.FILLER_0_16_161.VGND
rlabel metal1 5224 21376 5408 21472 1 sr_0.FILLER_0_16_161.VPWR
flabel metal1 4977 21407 5011 21441 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_16_Right_16.VPWR
flabel metal1 4977 20863 5011 20897 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_16_Right_16.VGND
flabel nwell 4977 21407 5011 21441 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_16_Right_16.VPB
flabel pwell 4977 20863 5011 20897 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_16_Right_16.VNB
rlabel comment 4948 20880 4948 20880 4 sr_0.PHY_EDGE_ROW_16_Right_16.decap_3
rlabel metal1 4948 20832 5224 20928 1 sr_0.PHY_EDGE_ROW_16_Right_16.VGND
rlabel metal1 4948 21376 5224 21472 1 sr_0.PHY_EDGE_ROW_16_Right_16.VPWR
flabel metal1 19881 21951 19915 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_3.VGND
flabel metal1 19881 21407 19915 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_3.VPWR
flabel nwell 19881 21407 19915 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_3.VPB
flabel pwell 19881 21951 19915 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_3.VNB
rlabel comment 19944 21968 19944 21968 8 sr_0.FILLER_0_17_3.decap_12
flabel metal1 18777 21951 18811 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_15.VGND
flabel metal1 18777 21407 18811 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_15.VPWR
flabel nwell 18777 21407 18811 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_15.VPB
flabel pwell 18777 21951 18811 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_15.VNB
rlabel comment 18840 21968 18840 21968 8 sr_0.FILLER_0_17_15.decap_12
flabel metal1 20157 21407 20191 21441 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_17_Left_45.VPWR
flabel metal1 20157 21951 20191 21985 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_17_Left_45.VGND
flabel nwell 20157 21407 20191 21441 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_17_Left_45.VPB
flabel pwell 20157 21951 20191 21985 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_17_Left_45.VNB
rlabel comment 20220 21968 20220 21968 8 sr_0.PHY_EDGE_ROW_17_Left_45.decap_3
rlabel metal1 19944 21920 20220 22016 5 sr_0.PHY_EDGE_ROW_17_Left_45.VGND
rlabel metal1 19944 21376 20220 21472 5 sr_0.PHY_EDGE_ROW_17_Left_45.VPWR
flabel metal1 17673 21951 17707 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_27.VGND
flabel metal1 17673 21407 17707 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_27.VPWR
flabel nwell 17673 21407 17707 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_27.VPB
flabel pwell 17673 21951 17707 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_27.VNB
rlabel comment 17736 21968 17736 21968 8 sr_0.FILLER_0_17_27.decap_12
flabel metal1 16569 21951 16603 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_39.VGND
flabel metal1 16569 21407 16603 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_39.VPWR
flabel nwell 16569 21407 16603 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_39.VPB
flabel pwell 16569 21951 16603 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_39.VNB
rlabel comment 16632 21968 16632 21968 8 sr_0.FILLER_0_17_39.decap_12
flabel metal1 15465 21951 15499 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_51.VGND
flabel metal1 15465 21407 15499 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_51.VPWR
flabel nwell 15465 21407 15499 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_51.VPB
flabel pwell 15465 21951 15499 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_51.VNB
rlabel comment 15528 21968 15528 21968 8 sr_0.FILLER_0_17_51.decap_4
rlabel metal1 15160 21920 15528 22016 5 sr_0.FILLER_0_17_51.VGND
rlabel metal1 15160 21376 15528 21472 5 sr_0.FILLER_0_17_51.VPWR
flabel metal1 15102 21411 15138 21441 0 FreeSans 250 0 0 0 sr_0.FILLER_0_17_55.VPWR
flabel metal1 15102 21952 15138 21981 0 FreeSans 250 0 0 0 sr_0.FILLER_0_17_55.VGND
flabel nwell 15109 21417 15129 21434 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_55.VPB
flabel pwell 15108 21957 15132 21979 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_55.VNB
rlabel comment 15160 21968 15160 21968 8 sr_0.FILLER_0_17_55.fill_1
rlabel metal1 15068 21920 15160 22016 5 sr_0.FILLER_0_17_55.VGND
rlabel metal1 15068 21376 15160 21472 5 sr_0.FILLER_0_17_55.VPWR
flabel metal1 14913 21951 14947 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_57.VGND
flabel metal1 14913 21407 14947 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_57.VPWR
flabel nwell 14913 21407 14947 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_57.VPB
flabel pwell 14913 21951 14947 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_57.VNB
rlabel comment 14976 21968 14976 21968 8 sr_0.FILLER_0_17_57.decap_12
flabel metal1 14993 21415 15046 21444 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_17_101.VPWR
flabel metal1 14996 21948 15047 21986 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_17_101.VGND
rlabel comment 15068 21968 15068 21968 8 sr_0.TAP_TAPCELL_ROW_17_101.tapvpwrvgnd_1
rlabel metal1 14976 21920 15068 22016 5 sr_0.TAP_TAPCELL_ROW_17_101.VGND
rlabel metal1 14976 21376 15068 21472 5 sr_0.TAP_TAPCELL_ROW_17_101.VPWR
flabel metal1 13809 21951 13843 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_69.VGND
flabel metal1 13809 21407 13843 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_69.VPWR
flabel nwell 13809 21407 13843 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_69.VPB
flabel pwell 13809 21951 13843 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_69.VNB
rlabel comment 13872 21968 13872 21968 8 sr_0.FILLER_0_17_69.decap_12
flabel metal1 12705 21951 12739 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_81.VGND
flabel metal1 12705 21407 12739 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_81.VPWR
flabel nwell 12705 21407 12739 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_81.VPB
flabel pwell 12705 21951 12739 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_81.VNB
rlabel comment 12768 21968 12768 21968 8 sr_0.FILLER_0_17_81.decap_12
flabel metal1 11601 21951 11635 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_93.VGND
flabel metal1 11601 21407 11635 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_93.VPWR
flabel nwell 11601 21407 11635 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_93.VPB
flabel pwell 11601 21951 11635 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_93.VNB
rlabel comment 11664 21968 11664 21968 8 sr_0.FILLER_0_17_93.decap_12
flabel metal1 10497 21407 10531 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_105.VPWR
flabel metal1 10497 21951 10531 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_105.VGND
flabel nwell 10497 21407 10531 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_105.VPB
flabel pwell 10497 21951 10531 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_105.VNB
rlabel comment 10560 21968 10560 21968 8 sr_0.FILLER_0_17_105.decap_6
rlabel metal1 10008 21920 10560 22016 5 sr_0.FILLER_0_17_105.VGND
rlabel metal1 10008 21376 10560 21472 5 sr_0.FILLER_0_17_105.VPWR
flabel metal1 9950 21411 9986 21441 0 FreeSans 250 0 0 0 sr_0.FILLER_0_17_111.VPWR
flabel metal1 9950 21952 9986 21981 0 FreeSans 250 0 0 0 sr_0.FILLER_0_17_111.VGND
flabel nwell 9957 21417 9977 21434 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_111.VPB
flabel pwell 9956 21957 9980 21979 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_111.VNB
rlabel comment 10008 21968 10008 21968 8 sr_0.FILLER_0_17_111.fill_1
rlabel metal1 9916 21920 10008 22016 5 sr_0.FILLER_0_17_111.VGND
rlabel metal1 9916 21376 10008 21472 5 sr_0.FILLER_0_17_111.VPWR
flabel metal1 9761 21951 9795 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_113.VGND
flabel metal1 9761 21407 9795 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_113.VPWR
flabel nwell 9761 21407 9795 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_113.VPB
flabel pwell 9761 21951 9795 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_113.VNB
rlabel comment 9824 21968 9824 21968 8 sr_0.FILLER_0_17_113.decap_12
flabel metal1 8657 21951 8691 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_125.VGND
flabel metal1 8657 21407 8691 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_125.VPWR
flabel nwell 8657 21407 8691 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_125.VPB
flabel pwell 8657 21951 8691 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_125.VNB
rlabel comment 8720 21968 8720 21968 8 sr_0.FILLER_0_17_125.decap_12
flabel metal1 9841 21415 9894 21444 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_17_102.VPWR
flabel metal1 9844 21948 9895 21986 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_17_102.VGND
rlabel comment 9916 21968 9916 21968 8 sr_0.TAP_TAPCELL_ROW_17_102.tapvpwrvgnd_1
rlabel metal1 9824 21920 9916 22016 5 sr_0.TAP_TAPCELL_ROW_17_102.VGND
rlabel metal1 9824 21376 9916 21472 5 sr_0.TAP_TAPCELL_ROW_17_102.VPWR
flabel metal1 7553 21951 7587 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_137.VGND
flabel metal1 7553 21407 7587 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_137.VPWR
flabel nwell 7553 21407 7587 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_137.VPB
flabel pwell 7553 21951 7587 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_137.VNB
rlabel comment 7616 21968 7616 21968 8 sr_0.FILLER_0_17_137.decap_12
flabel metal1 6449 21951 6483 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_149.VGND
flabel metal1 6449 21407 6483 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_149.VPWR
flabel nwell 6449 21407 6483 21441 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_149.VPB
flabel pwell 6449 21951 6483 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_149.VNB
rlabel comment 6512 21968 6512 21968 8 sr_0.FILLER_0_17_149.decap_12
flabel metal1 5335 21950 5388 21982 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_161.VGND
flabel metal1 5335 21407 5387 21438 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_161.VPWR
flabel nwell 5346 21415 5380 21433 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_161.VPB
flabel pwell 5345 21956 5377 21978 0 FreeSans 200 0 0 0 sr_0.FILLER_0_17_161.VNB
rlabel comment 5408 21968 5408 21968 8 sr_0.FILLER_0_17_161.fill_2
rlabel metal1 5224 21920 5408 22016 5 sr_0.FILLER_0_17_161.VGND
rlabel metal1 5224 21376 5408 21472 5 sr_0.FILLER_0_17_161.VPWR
flabel metal1 4977 21407 5011 21441 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_17_Right_17.VPWR
flabel metal1 4977 21951 5011 21985 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_17_Right_17.VGND
flabel nwell 4977 21407 5011 21441 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_17_Right_17.VPB
flabel pwell 4977 21951 5011 21985 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_17_Right_17.VNB
rlabel comment 4948 21968 4948 21968 2 sr_0.PHY_EDGE_ROW_17_Right_17.decap_3
rlabel metal1 4948 21920 5224 22016 5 sr_0.PHY_EDGE_ROW_17_Right_17.VGND
rlabel metal1 4948 21376 5224 21472 5 sr_0.PHY_EDGE_ROW_17_Right_17.VPWR
flabel metal1 19881 21951 19915 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_3.VGND
flabel metal1 19881 22495 19915 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_3.VPWR
flabel nwell 19881 22495 19915 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_3.VPB
flabel pwell 19881 21951 19915 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_3.VNB
rlabel comment 19944 21968 19944 21968 6 sr_0.FILLER_0_18_3.decap_12
flabel metal1 18777 21951 18811 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_15.VGND
flabel metal1 18777 22495 18811 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_15.VPWR
flabel nwell 18777 22495 18811 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_15.VPB
flabel pwell 18777 21951 18811 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_15.VNB
rlabel comment 18840 21968 18840 21968 6 sr_0.FILLER_0_18_15.decap_12
flabel metal1 20157 22495 20191 22529 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_18_Left_46.VPWR
flabel metal1 20157 21951 20191 21985 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_18_Left_46.VGND
flabel nwell 20157 22495 20191 22529 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_18_Left_46.VPB
flabel pwell 20157 21951 20191 21985 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_18_Left_46.VNB
rlabel comment 20220 21968 20220 21968 6 sr_0.PHY_EDGE_ROW_18_Left_46.decap_3
rlabel metal1 19944 21920 20220 22016 1 sr_0.PHY_EDGE_ROW_18_Left_46.VGND
rlabel metal1 19944 22464 20220 22560 1 sr_0.PHY_EDGE_ROW_18_Left_46.VPWR
flabel metal1 17678 22495 17714 22525 0 FreeSans 250 0 0 0 sr_0.FILLER_0_18_27.VPWR
flabel metal1 17678 21955 17714 21984 0 FreeSans 250 0 0 0 sr_0.FILLER_0_18_27.VGND
flabel nwell 17685 22502 17705 22519 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_27.VPB
flabel pwell 17684 21957 17708 21979 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_27.VNB
rlabel comment 17736 21968 17736 21968 6 sr_0.FILLER_0_18_27.fill_1
rlabel metal1 17644 21920 17736 22016 1 sr_0.FILLER_0_18_27.VGND
rlabel metal1 17644 22464 17736 22560 1 sr_0.FILLER_0_18_27.VPWR
flabel metal1 17489 21951 17523 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_29.VGND
flabel metal1 17489 22495 17523 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_29.VPWR
flabel nwell 17489 22495 17523 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_29.VPB
flabel pwell 17489 21951 17523 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_29.VNB
rlabel comment 17552 21968 17552 21968 6 sr_0.FILLER_0_18_29.decap_12
flabel metal1 16385 21951 16419 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_41.VGND
flabel metal1 16385 22495 16419 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_41.VPWR
flabel nwell 16385 22495 16419 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_41.VPB
flabel pwell 16385 21951 16419 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_41.VNB
rlabel comment 16448 21968 16448 21968 6 sr_0.FILLER_0_18_41.decap_12
flabel metal1 17569 22492 17622 22521 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_18_103.VPWR
flabel metal1 17572 21950 17623 21988 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_18_103.VGND
rlabel comment 17644 21968 17644 21968 6 sr_0.TAP_TAPCELL_ROW_18_103.tapvpwrvgnd_1
rlabel metal1 17552 21920 17644 22016 1 sr_0.TAP_TAPCELL_ROW_18_103.VGND
rlabel metal1 17552 22464 17644 22560 1 sr_0.TAP_TAPCELL_ROW_18_103.VPWR
flabel metal1 15281 21951 15315 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_53.VGND
flabel metal1 15281 22495 15315 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_53.VPWR
flabel nwell 15281 22495 15315 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_53.VPB
flabel pwell 15281 21951 15315 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_53.VNB
rlabel comment 15344 21968 15344 21968 6 sr_0.FILLER_0_18_53.decap_12
flabel metal1 14177 21951 14211 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_65.VGND
flabel metal1 14177 22495 14211 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_65.VPWR
flabel nwell 14177 22495 14211 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_65.VPB
flabel pwell 14177 21951 14211 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_65.VNB
rlabel comment 14240 21968 14240 21968 6 sr_0.FILLER_0_18_65.decap_12
flabel metal1 13073 22495 13107 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_77.VPWR
flabel metal1 13073 21951 13107 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_77.VGND
flabel nwell 13073 22495 13107 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_77.VPB
flabel pwell 13073 21951 13107 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_77.VNB
rlabel comment 13136 21968 13136 21968 6 sr_0.FILLER_0_18_77.decap_6
rlabel metal1 12584 21920 13136 22016 1 sr_0.FILLER_0_18_77.VGND
rlabel metal1 12584 22464 13136 22560 1 sr_0.FILLER_0_18_77.VPWR
flabel metal1 12526 22495 12562 22525 0 FreeSans 250 0 0 0 sr_0.FILLER_0_18_83.VPWR
flabel metal1 12526 21955 12562 21984 0 FreeSans 250 0 0 0 sr_0.FILLER_0_18_83.VGND
flabel nwell 12533 22502 12553 22519 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_83.VPB
flabel pwell 12532 21957 12556 21979 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_83.VNB
rlabel comment 12584 21968 12584 21968 6 sr_0.FILLER_0_18_83.fill_1
rlabel metal1 12492 21920 12584 22016 1 sr_0.FILLER_0_18_83.VGND
rlabel metal1 12492 22464 12584 22560 1 sr_0.FILLER_0_18_83.VPWR
flabel metal1 12337 21951 12371 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_85.VGND
flabel metal1 12337 22495 12371 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_85.VPWR
flabel nwell 12337 22495 12371 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_85.VPB
flabel pwell 12337 21951 12371 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_85.VNB
rlabel comment 12400 21968 12400 21968 6 sr_0.FILLER_0_18_85.decap_12
flabel metal1 11233 21951 11267 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_97.VGND
flabel metal1 11233 22495 11267 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_97.VPWR
flabel nwell 11233 22495 11267 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_97.VPB
flabel pwell 11233 21951 11267 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_97.VNB
rlabel comment 11296 21968 11296 21968 6 sr_0.FILLER_0_18_97.decap_12
flabel metal1 12417 22492 12470 22521 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_18_104.VPWR
flabel metal1 12420 21950 12471 21988 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_18_104.VGND
rlabel comment 12492 21968 12492 21968 6 sr_0.TAP_TAPCELL_ROW_18_104.tapvpwrvgnd_1
rlabel metal1 12400 21920 12492 22016 1 sr_0.TAP_TAPCELL_ROW_18_104.VGND
rlabel metal1 12400 22464 12492 22560 1 sr_0.TAP_TAPCELL_ROW_18_104.VPWR
flabel metal1 10129 21951 10163 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_109.VGND
flabel metal1 10129 22495 10163 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_109.VPWR
flabel nwell 10129 22495 10163 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_109.VPB
flabel pwell 10129 21951 10163 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_109.VNB
rlabel comment 10192 21968 10192 21968 6 sr_0.FILLER_0_18_109.decap_12
flabel metal1 9025 21951 9059 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_121.VGND
flabel metal1 9025 22495 9059 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_121.VPWR
flabel nwell 9025 22495 9059 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_121.VPB
flabel pwell 9025 21951 9059 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_121.VNB
rlabel comment 9088 21968 9088 21968 6 sr_0.FILLER_0_18_121.decap_12
flabel metal1 7921 22495 7955 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_133.VPWR
flabel metal1 7921 21951 7955 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_133.VGND
flabel nwell 7921 22495 7955 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_133.VPB
flabel pwell 7921 21951 7955 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_133.VNB
rlabel comment 7984 21968 7984 21968 6 sr_0.FILLER_0_18_133.decap_6
rlabel metal1 7432 21920 7984 22016 1 sr_0.FILLER_0_18_133.VGND
rlabel metal1 7432 22464 7984 22560 1 sr_0.FILLER_0_18_133.VPWR
flabel metal1 7374 22495 7410 22525 0 FreeSans 250 0 0 0 sr_0.FILLER_0_18_139.VPWR
flabel metal1 7374 21955 7410 21984 0 FreeSans 250 0 0 0 sr_0.FILLER_0_18_139.VGND
flabel nwell 7381 22502 7401 22519 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_139.VPB
flabel pwell 7380 21957 7404 21979 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_139.VNB
rlabel comment 7432 21968 7432 21968 6 sr_0.FILLER_0_18_139.fill_1
rlabel metal1 7340 21920 7432 22016 1 sr_0.FILLER_0_18_139.VGND
rlabel metal1 7340 22464 7432 22560 1 sr_0.FILLER_0_18_139.VPWR
flabel metal1 7185 21951 7219 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_141.VGND
flabel metal1 7185 22495 7219 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_141.VPWR
flabel nwell 7185 22495 7219 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_141.VPB
flabel pwell 7185 21951 7219 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_141.VNB
rlabel comment 7248 21968 7248 21968 6 sr_0.FILLER_0_18_141.decap_12
flabel metal1 7265 22492 7318 22521 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_18_105.VPWR
flabel metal1 7268 21950 7319 21988 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_18_105.VGND
rlabel comment 7340 21968 7340 21968 6 sr_0.TAP_TAPCELL_ROW_18_105.tapvpwrvgnd_1
rlabel metal1 7248 21920 7340 22016 1 sr_0.TAP_TAPCELL_ROW_18_105.VGND
rlabel metal1 7248 22464 7340 22560 1 sr_0.TAP_TAPCELL_ROW_18_105.VPWR
flabel metal1 6081 22495 6115 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_153.VPWR
flabel metal1 6081 21951 6115 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_153.VGND
flabel nwell 6081 22495 6115 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_153.VPB
flabel pwell 6081 21951 6115 21985 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_153.VNB
rlabel comment 6144 21968 6144 21968 6 sr_0.FILLER_0_18_153.decap_8
rlabel metal1 5408 21920 6144 22016 1 sr_0.FILLER_0_18_153.VGND
rlabel metal1 5408 22464 6144 22560 1 sr_0.FILLER_0_18_153.VPWR
flabel metal1 5335 21954 5388 21986 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_161.VGND
flabel metal1 5335 22498 5387 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_161.VPWR
flabel nwell 5346 22503 5380 22521 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_161.VPB
flabel pwell 5345 21958 5377 21980 0 FreeSans 200 0 0 0 sr_0.FILLER_0_18_161.VNB
rlabel comment 5408 21968 5408 21968 6 sr_0.FILLER_0_18_161.fill_2
rlabel metal1 5224 21920 5408 22016 1 sr_0.FILLER_0_18_161.VGND
rlabel metal1 5224 22464 5408 22560 1 sr_0.FILLER_0_18_161.VPWR
flabel metal1 4977 22495 5011 22529 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_18_Right_18.VPWR
flabel metal1 4977 21951 5011 21985 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_18_Right_18.VGND
flabel nwell 4977 22495 5011 22529 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_18_Right_18.VPB
flabel pwell 4977 21951 5011 21985 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_18_Right_18.VNB
rlabel comment 4948 21968 4948 21968 4 sr_0.PHY_EDGE_ROW_18_Right_18.decap_3
rlabel metal1 4948 21920 5224 22016 1 sr_0.PHY_EDGE_ROW_18_Right_18.VGND
rlabel metal1 4948 22464 5224 22560 1 sr_0.PHY_EDGE_ROW_18_Right_18.VPWR
flabel metal1 19881 23039 19915 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_3.VGND
flabel metal1 19881 22495 19915 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_3.VPWR
flabel nwell 19881 22495 19915 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_3.VPB
flabel pwell 19881 23039 19915 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_3.VNB
rlabel comment 19944 23056 19944 23056 8 sr_0.FILLER_0_19_3.decap_12
flabel metal1 18777 23039 18811 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_15.VGND
flabel metal1 18777 22495 18811 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_15.VPWR
flabel nwell 18777 22495 18811 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_15.VPB
flabel pwell 18777 23039 18811 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_15.VNB
rlabel comment 18840 23056 18840 23056 8 sr_0.FILLER_0_19_15.decap_12
flabel metal1 19881 23039 19915 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_3.VGND
flabel metal1 19881 23583 19915 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_3.VPWR
flabel nwell 19881 23583 19915 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_3.VPB
flabel pwell 19881 23039 19915 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_3.VNB
rlabel comment 19944 23056 19944 23056 6 sr_0.FILLER_0_20_3.decap_12
flabel metal1 18777 23039 18811 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_15.VGND
flabel metal1 18777 23583 18811 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_15.VPWR
flabel nwell 18777 23583 18811 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_15.VPB
flabel pwell 18777 23039 18811 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_15.VNB
rlabel comment 18840 23056 18840 23056 6 sr_0.FILLER_0_20_15.decap_12
flabel metal1 20157 22495 20191 22529 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_19_Left_47.VPWR
flabel metal1 20157 23039 20191 23073 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_19_Left_47.VGND
flabel nwell 20157 22495 20191 22529 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_19_Left_47.VPB
flabel pwell 20157 23039 20191 23073 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_19_Left_47.VNB
rlabel comment 20220 23056 20220 23056 8 sr_0.PHY_EDGE_ROW_19_Left_47.decap_3
rlabel metal1 19944 23008 20220 23104 5 sr_0.PHY_EDGE_ROW_19_Left_47.VGND
rlabel metal1 19944 22464 20220 22560 5 sr_0.PHY_EDGE_ROW_19_Left_47.VPWR
flabel metal1 20157 23583 20191 23617 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_20_Left_48.VPWR
flabel metal1 20157 23039 20191 23073 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_20_Left_48.VGND
flabel nwell 20157 23583 20191 23617 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_20_Left_48.VPB
flabel pwell 20157 23039 20191 23073 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_20_Left_48.VNB
rlabel comment 20220 23056 20220 23056 6 sr_0.PHY_EDGE_ROW_20_Left_48.decap_3
rlabel metal1 19944 23008 20220 23104 1 sr_0.PHY_EDGE_ROW_20_Left_48.VGND
rlabel metal1 19944 23552 20220 23648 1 sr_0.PHY_EDGE_ROW_20_Left_48.VPWR
flabel metal1 17673 23039 17707 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_27.VGND
flabel metal1 17673 22495 17707 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_27.VPWR
flabel nwell 17673 22495 17707 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_27.VPB
flabel pwell 17673 23039 17707 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_27.VNB
rlabel comment 17736 23056 17736 23056 8 sr_0.FILLER_0_19_27.decap_12
flabel metal1 16569 23039 16603 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_39.VGND
flabel metal1 16569 22495 16603 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_39.VPWR
flabel nwell 16569 22495 16603 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_39.VPB
flabel pwell 16569 23039 16603 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_39.VNB
rlabel comment 16632 23056 16632 23056 8 sr_0.FILLER_0_19_39.decap_12
flabel metal1 17678 23583 17714 23613 0 FreeSans 250 0 0 0 sr_0.FILLER_0_20_27.VPWR
flabel metal1 17678 23043 17714 23072 0 FreeSans 250 0 0 0 sr_0.FILLER_0_20_27.VGND
flabel nwell 17685 23590 17705 23607 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_27.VPB
flabel pwell 17684 23045 17708 23067 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_27.VNB
rlabel comment 17736 23056 17736 23056 6 sr_0.FILLER_0_20_27.fill_1
rlabel metal1 17644 23008 17736 23104 1 sr_0.FILLER_0_20_27.VGND
rlabel metal1 17644 23552 17736 23648 1 sr_0.FILLER_0_20_27.VPWR
flabel metal1 17489 23039 17523 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_29.VGND
flabel metal1 17489 23583 17523 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_29.VPWR
flabel nwell 17489 23583 17523 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_29.VPB
flabel pwell 17489 23039 17523 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_29.VNB
rlabel comment 17552 23056 17552 23056 6 sr_0.FILLER_0_20_29.decap_12
flabel metal1 16385 23039 16419 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_41.VGND
flabel metal1 16385 23583 16419 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_41.VPWR
flabel nwell 16385 23583 16419 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_41.VPB
flabel pwell 16385 23039 16419 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_41.VNB
rlabel comment 16448 23056 16448 23056 6 sr_0.FILLER_0_20_41.decap_12
flabel metal1 17569 23580 17622 23609 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_20_108.VPWR
flabel metal1 17572 23038 17623 23076 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_20_108.VGND
rlabel comment 17644 23056 17644 23056 6 sr_0.TAP_TAPCELL_ROW_20_108.tapvpwrvgnd_1
rlabel metal1 17552 23008 17644 23104 1 sr_0.TAP_TAPCELL_ROW_20_108.VGND
rlabel metal1 17552 23552 17644 23648 1 sr_0.TAP_TAPCELL_ROW_20_108.VPWR
flabel metal1 15465 23039 15499 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_51.VGND
flabel metal1 15465 22495 15499 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_51.VPWR
flabel nwell 15465 22495 15499 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_51.VPB
flabel pwell 15465 23039 15499 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_51.VNB
rlabel comment 15528 23056 15528 23056 8 sr_0.FILLER_0_19_51.decap_4
rlabel metal1 15160 23008 15528 23104 5 sr_0.FILLER_0_19_51.VGND
rlabel metal1 15160 22464 15528 22560 5 sr_0.FILLER_0_19_51.VPWR
flabel metal1 15102 22499 15138 22529 0 FreeSans 250 0 0 0 sr_0.FILLER_0_19_55.VPWR
flabel metal1 15102 23040 15138 23069 0 FreeSans 250 0 0 0 sr_0.FILLER_0_19_55.VGND
flabel nwell 15109 22505 15129 22522 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_55.VPB
flabel pwell 15108 23045 15132 23067 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_55.VNB
rlabel comment 15160 23056 15160 23056 8 sr_0.FILLER_0_19_55.fill_1
rlabel metal1 15068 23008 15160 23104 5 sr_0.FILLER_0_19_55.VGND
rlabel metal1 15068 22464 15160 22560 5 sr_0.FILLER_0_19_55.VPWR
flabel metal1 14913 23039 14947 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_57.VGND
flabel metal1 14913 22495 14947 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_57.VPWR
flabel nwell 14913 22495 14947 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_57.VPB
flabel pwell 14913 23039 14947 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_57.VNB
rlabel comment 14976 23056 14976 23056 8 sr_0.FILLER_0_19_57.decap_12
flabel metal1 15281 23039 15315 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_53.VGND
flabel metal1 15281 23583 15315 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_53.VPWR
flabel nwell 15281 23583 15315 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_53.VPB
flabel pwell 15281 23039 15315 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_53.VNB
rlabel comment 15344 23056 15344 23056 6 sr_0.FILLER_0_20_53.decap_12
flabel metal1 14993 22503 15046 22532 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_19_106.VPWR
flabel metal1 14996 23036 15047 23074 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_19_106.VGND
rlabel comment 15068 23056 15068 23056 8 sr_0.TAP_TAPCELL_ROW_19_106.tapvpwrvgnd_1
rlabel metal1 14976 23008 15068 23104 5 sr_0.TAP_TAPCELL_ROW_19_106.VGND
rlabel metal1 14976 22464 15068 22560 5 sr_0.TAP_TAPCELL_ROW_19_106.VPWR
flabel metal1 13809 23039 13843 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_69.VGND
flabel metal1 13809 22495 13843 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_69.VPWR
flabel nwell 13809 22495 13843 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_69.VPB
flabel pwell 13809 23039 13843 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_69.VNB
rlabel comment 13872 23056 13872 23056 8 sr_0.FILLER_0_19_69.decap_12
flabel metal1 12705 23039 12739 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_81.VGND
flabel metal1 12705 22495 12739 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_81.VPWR
flabel nwell 12705 22495 12739 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_81.VPB
flabel pwell 12705 23039 12739 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_81.VNB
rlabel comment 12768 23056 12768 23056 8 sr_0.FILLER_0_19_81.decap_12
flabel metal1 14177 23039 14211 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_65.VGND
flabel metal1 14177 23583 14211 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_65.VPWR
flabel nwell 14177 23583 14211 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_65.VPB
flabel pwell 14177 23039 14211 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_65.VNB
rlabel comment 14240 23056 14240 23056 6 sr_0.FILLER_0_20_65.decap_12
flabel metal1 13073 23583 13107 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_77.VPWR
flabel metal1 13073 23039 13107 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_77.VGND
flabel nwell 13073 23583 13107 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_77.VPB
flabel pwell 13073 23039 13107 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_77.VNB
rlabel comment 13136 23056 13136 23056 6 sr_0.FILLER_0_20_77.decap_6
rlabel metal1 12584 23008 13136 23104 1 sr_0.FILLER_0_20_77.VGND
rlabel metal1 12584 23552 13136 23648 1 sr_0.FILLER_0_20_77.VPWR
flabel metal1 12526 23583 12562 23613 0 FreeSans 250 0 0 0 sr_0.FILLER_0_20_83.VPWR
flabel metal1 12526 23043 12562 23072 0 FreeSans 250 0 0 0 sr_0.FILLER_0_20_83.VGND
flabel nwell 12533 23590 12553 23607 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_83.VPB
flabel pwell 12532 23045 12556 23067 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_83.VNB
rlabel comment 12584 23056 12584 23056 6 sr_0.FILLER_0_20_83.fill_1
rlabel metal1 12492 23008 12584 23104 1 sr_0.FILLER_0_20_83.VGND
rlabel metal1 12492 23552 12584 23648 1 sr_0.FILLER_0_20_83.VPWR
flabel metal1 11601 23039 11635 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_93.VGND
flabel metal1 11601 22495 11635 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_93.VPWR
flabel nwell 11601 22495 11635 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_93.VPB
flabel pwell 11601 23039 11635 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_93.VNB
rlabel comment 11664 23056 11664 23056 8 sr_0.FILLER_0_19_93.decap_12
flabel metal1 12337 23039 12371 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_85.VGND
flabel metal1 12337 23583 12371 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_85.VPWR
flabel nwell 12337 23583 12371 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_85.VPB
flabel pwell 12337 23039 12371 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_85.VNB
rlabel comment 12400 23056 12400 23056 6 sr_0.FILLER_0_20_85.decap_12
flabel metal1 11233 23039 11267 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_97.VGND
flabel metal1 11233 23583 11267 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_97.VPWR
flabel nwell 11233 23583 11267 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_97.VPB
flabel pwell 11233 23039 11267 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_97.VNB
rlabel comment 11296 23056 11296 23056 6 sr_0.FILLER_0_20_97.decap_12
flabel metal1 12417 23580 12470 23609 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_20_109.VPWR
flabel metal1 12420 23038 12471 23076 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_20_109.VGND
rlabel comment 12492 23056 12492 23056 6 sr_0.TAP_TAPCELL_ROW_20_109.tapvpwrvgnd_1
rlabel metal1 12400 23008 12492 23104 1 sr_0.TAP_TAPCELL_ROW_20_109.VGND
rlabel metal1 12400 23552 12492 23648 1 sr_0.TAP_TAPCELL_ROW_20_109.VPWR
flabel metal1 10497 22495 10531 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_105.VPWR
flabel metal1 10497 23039 10531 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_105.VGND
flabel nwell 10497 22495 10531 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_105.VPB
flabel pwell 10497 23039 10531 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_105.VNB
rlabel comment 10560 23056 10560 23056 8 sr_0.FILLER_0_19_105.decap_6
rlabel metal1 10008 23008 10560 23104 5 sr_0.FILLER_0_19_105.VGND
rlabel metal1 10008 22464 10560 22560 5 sr_0.FILLER_0_19_105.VPWR
flabel metal1 9950 22499 9986 22529 0 FreeSans 250 0 0 0 sr_0.FILLER_0_19_111.VPWR
flabel metal1 9950 23040 9986 23069 0 FreeSans 250 0 0 0 sr_0.FILLER_0_19_111.VGND
flabel nwell 9957 22505 9977 22522 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_111.VPB
flabel pwell 9956 23045 9980 23067 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_111.VNB
rlabel comment 10008 23056 10008 23056 8 sr_0.FILLER_0_19_111.fill_1
rlabel metal1 9916 23008 10008 23104 5 sr_0.FILLER_0_19_111.VGND
rlabel metal1 9916 22464 10008 22560 5 sr_0.FILLER_0_19_111.VPWR
flabel metal1 9761 23039 9795 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_113.VGND
flabel metal1 9761 22495 9795 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_113.VPWR
flabel nwell 9761 22495 9795 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_113.VPB
flabel pwell 9761 23039 9795 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_113.VNB
rlabel comment 9824 23056 9824 23056 8 sr_0.FILLER_0_19_113.decap_12
flabel metal1 8657 23039 8691 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_125.VGND
flabel metal1 8657 22495 8691 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_125.VPWR
flabel nwell 8657 22495 8691 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_125.VPB
flabel pwell 8657 23039 8691 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_125.VNB
rlabel comment 8720 23056 8720 23056 8 sr_0.FILLER_0_19_125.decap_12
flabel metal1 10129 23039 10163 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_109.VGND
flabel metal1 10129 23583 10163 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_109.VPWR
flabel nwell 10129 23583 10163 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_109.VPB
flabel pwell 10129 23039 10163 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_109.VNB
rlabel comment 10192 23056 10192 23056 6 sr_0.FILLER_0_20_109.decap_12
flabel metal1 9025 23039 9059 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_121.VGND
flabel metal1 9025 23583 9059 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_121.VPWR
flabel nwell 9025 23583 9059 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_121.VPB
flabel pwell 9025 23039 9059 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_121.VNB
rlabel comment 9088 23056 9088 23056 6 sr_0.FILLER_0_20_121.decap_12
flabel metal1 9841 22503 9894 22532 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_19_107.VPWR
flabel metal1 9844 23036 9895 23074 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_19_107.VGND
rlabel comment 9916 23056 9916 23056 8 sr_0.TAP_TAPCELL_ROW_19_107.tapvpwrvgnd_1
rlabel metal1 9824 23008 9916 23104 5 sr_0.TAP_TAPCELL_ROW_19_107.VGND
rlabel metal1 9824 22464 9916 22560 5 sr_0.TAP_TAPCELL_ROW_19_107.VPWR
flabel metal1 7553 23039 7587 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_137.VGND
flabel metal1 7553 22495 7587 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_137.VPWR
flabel nwell 7553 22495 7587 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_137.VPB
flabel pwell 7553 23039 7587 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_137.VNB
rlabel comment 7616 23056 7616 23056 8 sr_0.FILLER_0_19_137.decap_12
flabel metal1 7921 23583 7955 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_133.VPWR
flabel metal1 7921 23039 7955 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_133.VGND
flabel nwell 7921 23583 7955 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_133.VPB
flabel pwell 7921 23039 7955 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_133.VNB
rlabel comment 7984 23056 7984 23056 6 sr_0.FILLER_0_20_133.decap_6
rlabel metal1 7432 23008 7984 23104 1 sr_0.FILLER_0_20_133.VGND
rlabel metal1 7432 23552 7984 23648 1 sr_0.FILLER_0_20_133.VPWR
flabel metal1 7374 23583 7410 23613 0 FreeSans 250 0 0 0 sr_0.FILLER_0_20_139.VPWR
flabel metal1 7374 23043 7410 23072 0 FreeSans 250 0 0 0 sr_0.FILLER_0_20_139.VGND
flabel nwell 7381 23590 7401 23607 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_139.VPB
flabel pwell 7380 23045 7404 23067 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_139.VNB
rlabel comment 7432 23056 7432 23056 6 sr_0.FILLER_0_20_139.fill_1
rlabel metal1 7340 23008 7432 23104 1 sr_0.FILLER_0_20_139.VGND
rlabel metal1 7340 23552 7432 23648 1 sr_0.FILLER_0_20_139.VPWR
flabel metal1 7185 23039 7219 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_141.VGND
flabel metal1 7185 23583 7219 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_141.VPWR
flabel nwell 7185 23583 7219 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_141.VPB
flabel pwell 7185 23039 7219 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_141.VNB
rlabel comment 7248 23056 7248 23056 6 sr_0.FILLER_0_20_141.decap_12
flabel metal1 7265 23580 7318 23609 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_20_110.VPWR
flabel metal1 7268 23038 7319 23076 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_20_110.VGND
rlabel comment 7340 23056 7340 23056 6 sr_0.TAP_TAPCELL_ROW_20_110.tapvpwrvgnd_1
rlabel metal1 7248 23008 7340 23104 1 sr_0.TAP_TAPCELL_ROW_20_110.VGND
rlabel metal1 7248 23552 7340 23648 1 sr_0.TAP_TAPCELL_ROW_20_110.VPWR
flabel metal1 6449 23039 6483 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_149.VGND
flabel metal1 6449 22495 6483 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_149.VPWR
flabel nwell 6449 22495 6483 22529 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_149.VPB
flabel pwell 6449 23039 6483 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_149.VNB
rlabel comment 6512 23056 6512 23056 8 sr_0.FILLER_0_19_149.decap_12
flabel metal1 5335 23038 5388 23070 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_161.VGND
flabel metal1 5335 22495 5387 22526 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_161.VPWR
flabel nwell 5346 22503 5380 22521 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_161.VPB
flabel pwell 5345 23044 5377 23066 0 FreeSans 200 0 0 0 sr_0.FILLER_0_19_161.VNB
rlabel comment 5408 23056 5408 23056 8 sr_0.FILLER_0_19_161.fill_2
rlabel metal1 5224 23008 5408 23104 5 sr_0.FILLER_0_19_161.VGND
rlabel metal1 5224 22464 5408 22560 5 sr_0.FILLER_0_19_161.VPWR
flabel metal1 6081 23583 6115 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_153.VPWR
flabel metal1 6081 23039 6115 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_153.VGND
flabel nwell 6081 23583 6115 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_153.VPB
flabel pwell 6081 23039 6115 23073 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_153.VNB
rlabel comment 6144 23056 6144 23056 6 sr_0.FILLER_0_20_153.decap_8
rlabel metal1 5408 23008 6144 23104 1 sr_0.FILLER_0_20_153.VGND
rlabel metal1 5408 23552 6144 23648 1 sr_0.FILLER_0_20_153.VPWR
flabel metal1 5335 23042 5388 23074 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_161.VGND
flabel metal1 5335 23586 5387 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_161.VPWR
flabel nwell 5346 23591 5380 23609 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_161.VPB
flabel pwell 5345 23046 5377 23068 0 FreeSans 200 0 0 0 sr_0.FILLER_0_20_161.VNB
rlabel comment 5408 23056 5408 23056 6 sr_0.FILLER_0_20_161.fill_2
rlabel metal1 5224 23008 5408 23104 1 sr_0.FILLER_0_20_161.VGND
rlabel metal1 5224 23552 5408 23648 1 sr_0.FILLER_0_20_161.VPWR
flabel metal1 4977 22495 5011 22529 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_19_Right_19.VPWR
flabel metal1 4977 23039 5011 23073 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_19_Right_19.VGND
flabel nwell 4977 22495 5011 22529 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_19_Right_19.VPB
flabel pwell 4977 23039 5011 23073 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_19_Right_19.VNB
rlabel comment 4948 23056 4948 23056 2 sr_0.PHY_EDGE_ROW_19_Right_19.decap_3
rlabel metal1 4948 23008 5224 23104 5 sr_0.PHY_EDGE_ROW_19_Right_19.VGND
rlabel metal1 4948 22464 5224 22560 5 sr_0.PHY_EDGE_ROW_19_Right_19.VPWR
flabel metal1 4977 23583 5011 23617 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_20_Right_20.VPWR
flabel metal1 4977 23039 5011 23073 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_20_Right_20.VGND
flabel nwell 4977 23583 5011 23617 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_20_Right_20.VPB
flabel pwell 4977 23039 5011 23073 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_20_Right_20.VNB
rlabel comment 4948 23056 4948 23056 4 sr_0.PHY_EDGE_ROW_20_Right_20.decap_3
rlabel metal1 4948 23008 5224 23104 1 sr_0.PHY_EDGE_ROW_20_Right_20.VGND
rlabel metal1 4948 23552 5224 23648 1 sr_0.PHY_EDGE_ROW_20_Right_20.VPWR
flabel metal1 19881 24127 19915 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_3.VGND
flabel metal1 19881 23583 19915 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_3.VPWR
flabel nwell 19881 23583 19915 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_3.VPB
flabel pwell 19881 24127 19915 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_3.VNB
rlabel comment 19944 24144 19944 24144 8 sr_0.FILLER_0_21_3.decap_12
flabel metal1 18777 24127 18811 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_15.VGND
flabel metal1 18777 23583 18811 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_15.VPWR
flabel nwell 18777 23583 18811 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_15.VPB
flabel pwell 18777 24127 18811 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_15.VNB
rlabel comment 18840 24144 18840 24144 8 sr_0.FILLER_0_21_15.decap_12
flabel metal1 20157 23583 20191 23617 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_21_Left_49.VPWR
flabel metal1 20157 24127 20191 24161 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_21_Left_49.VGND
flabel nwell 20157 23583 20191 23617 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_21_Left_49.VPB
flabel pwell 20157 24127 20191 24161 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_21_Left_49.VNB
rlabel comment 20220 24144 20220 24144 8 sr_0.PHY_EDGE_ROW_21_Left_49.decap_3
rlabel metal1 19944 24096 20220 24192 5 sr_0.PHY_EDGE_ROW_21_Left_49.VGND
rlabel metal1 19944 23552 20220 23648 5 sr_0.PHY_EDGE_ROW_21_Left_49.VPWR
flabel metal1 17673 24127 17707 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_27.VGND
flabel metal1 17673 23583 17707 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_27.VPWR
flabel nwell 17673 23583 17707 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_27.VPB
flabel pwell 17673 24127 17707 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_27.VNB
rlabel comment 17736 24144 17736 24144 8 sr_0.FILLER_0_21_27.decap_12
flabel metal1 16569 24127 16603 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_39.VGND
flabel metal1 16569 23583 16603 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_39.VPWR
flabel nwell 16569 23583 16603 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_39.VPB
flabel pwell 16569 24127 16603 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_39.VNB
rlabel comment 16632 24144 16632 24144 8 sr_0.FILLER_0_21_39.decap_12
flabel metal1 15465 24127 15499 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_51.VGND
flabel metal1 15465 23583 15499 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_51.VPWR
flabel nwell 15465 23583 15499 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_51.VPB
flabel pwell 15465 24127 15499 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_51.VNB
rlabel comment 15528 24144 15528 24144 8 sr_0.FILLER_0_21_51.decap_4
rlabel metal1 15160 24096 15528 24192 5 sr_0.FILLER_0_21_51.VGND
rlabel metal1 15160 23552 15528 23648 5 sr_0.FILLER_0_21_51.VPWR
flabel metal1 15102 23587 15138 23617 0 FreeSans 250 0 0 0 sr_0.FILLER_0_21_55.VPWR
flabel metal1 15102 24128 15138 24157 0 FreeSans 250 0 0 0 sr_0.FILLER_0_21_55.VGND
flabel nwell 15109 23593 15129 23610 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_55.VPB
flabel pwell 15108 24133 15132 24155 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_55.VNB
rlabel comment 15160 24144 15160 24144 8 sr_0.FILLER_0_21_55.fill_1
rlabel metal1 15068 24096 15160 24192 5 sr_0.FILLER_0_21_55.VGND
rlabel metal1 15068 23552 15160 23648 5 sr_0.FILLER_0_21_55.VPWR
flabel metal1 14913 24127 14947 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_57.VGND
flabel metal1 14913 23583 14947 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_57.VPWR
flabel nwell 14913 23583 14947 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_57.VPB
flabel pwell 14913 24127 14947 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_57.VNB
rlabel comment 14976 24144 14976 24144 8 sr_0.FILLER_0_21_57.decap_12
flabel metal1 14993 23591 15046 23620 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_21_111.VPWR
flabel metal1 14996 24124 15047 24162 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_21_111.VGND
rlabel comment 15068 24144 15068 24144 8 sr_0.TAP_TAPCELL_ROW_21_111.tapvpwrvgnd_1
rlabel metal1 14976 24096 15068 24192 5 sr_0.TAP_TAPCELL_ROW_21_111.VGND
rlabel metal1 14976 23552 15068 23648 5 sr_0.TAP_TAPCELL_ROW_21_111.VPWR
flabel metal1 13809 24127 13843 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_69.VGND
flabel metal1 13809 23583 13843 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_69.VPWR
flabel nwell 13809 23583 13843 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_69.VPB
flabel pwell 13809 24127 13843 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_69.VNB
rlabel comment 13872 24144 13872 24144 8 sr_0.FILLER_0_21_69.decap_12
flabel metal1 12705 24127 12739 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_81.VGND
flabel metal1 12705 23583 12739 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_81.VPWR
flabel nwell 12705 23583 12739 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_81.VPB
flabel pwell 12705 24127 12739 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_81.VNB
rlabel comment 12768 24144 12768 24144 8 sr_0.FILLER_0_21_81.decap_12
flabel metal1 11601 24127 11635 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_93.VGND
flabel metal1 11601 23583 11635 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_93.VPWR
flabel nwell 11601 23583 11635 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_93.VPB
flabel pwell 11601 24127 11635 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_93.VNB
rlabel comment 11664 24144 11664 24144 8 sr_0.FILLER_0_21_93.decap_12
flabel metal1 10497 23583 10531 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_105.VPWR
flabel metal1 10497 24127 10531 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_105.VGND
flabel nwell 10497 23583 10531 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_105.VPB
flabel pwell 10497 24127 10531 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_105.VNB
rlabel comment 10560 24144 10560 24144 8 sr_0.FILLER_0_21_105.decap_6
rlabel metal1 10008 24096 10560 24192 5 sr_0.FILLER_0_21_105.VGND
rlabel metal1 10008 23552 10560 23648 5 sr_0.FILLER_0_21_105.VPWR
flabel metal1 9950 23587 9986 23617 0 FreeSans 250 0 0 0 sr_0.FILLER_0_21_111.VPWR
flabel metal1 9950 24128 9986 24157 0 FreeSans 250 0 0 0 sr_0.FILLER_0_21_111.VGND
flabel nwell 9957 23593 9977 23610 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_111.VPB
flabel pwell 9956 24133 9980 24155 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_111.VNB
rlabel comment 10008 24144 10008 24144 8 sr_0.FILLER_0_21_111.fill_1
rlabel metal1 9916 24096 10008 24192 5 sr_0.FILLER_0_21_111.VGND
rlabel metal1 9916 23552 10008 23648 5 sr_0.FILLER_0_21_111.VPWR
flabel metal1 9761 24127 9795 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_113.VGND
flabel metal1 9761 23583 9795 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_113.VPWR
flabel nwell 9761 23583 9795 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_113.VPB
flabel pwell 9761 24127 9795 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_113.VNB
rlabel comment 9824 24144 9824 24144 8 sr_0.FILLER_0_21_113.decap_12
flabel metal1 8657 24127 8691 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_125.VGND
flabel metal1 8657 23583 8691 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_125.VPWR
flabel nwell 8657 23583 8691 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_125.VPB
flabel pwell 8657 24127 8691 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_125.VNB
rlabel comment 8720 24144 8720 24144 8 sr_0.FILLER_0_21_125.decap_12
flabel metal1 9841 23591 9894 23620 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_21_112.VPWR
flabel metal1 9844 24124 9895 24162 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_21_112.VGND
rlabel comment 9916 24144 9916 24144 8 sr_0.TAP_TAPCELL_ROW_21_112.tapvpwrvgnd_1
rlabel metal1 9824 24096 9916 24192 5 sr_0.TAP_TAPCELL_ROW_21_112.VGND
rlabel metal1 9824 23552 9916 23648 5 sr_0.TAP_TAPCELL_ROW_21_112.VPWR
flabel metal1 7553 24127 7587 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_137.VGND
flabel metal1 7553 23583 7587 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_137.VPWR
flabel nwell 7553 23583 7587 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_137.VPB
flabel pwell 7553 24127 7587 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_137.VNB
rlabel comment 7616 24144 7616 24144 8 sr_0.FILLER_0_21_137.decap_12
flabel metal1 6449 24127 6483 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_149.VGND
flabel metal1 6449 23583 6483 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_149.VPWR
flabel nwell 6449 23583 6483 23617 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_149.VPB
flabel pwell 6449 24127 6483 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_149.VNB
rlabel comment 6512 24144 6512 24144 8 sr_0.FILLER_0_21_149.decap_12
flabel metal1 5335 24126 5388 24158 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_161.VGND
flabel metal1 5335 23583 5387 23614 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_161.VPWR
flabel nwell 5346 23591 5380 23609 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_161.VPB
flabel pwell 5345 24132 5377 24154 0 FreeSans 200 0 0 0 sr_0.FILLER_0_21_161.VNB
rlabel comment 5408 24144 5408 24144 8 sr_0.FILLER_0_21_161.fill_2
rlabel metal1 5224 24096 5408 24192 5 sr_0.FILLER_0_21_161.VGND
rlabel metal1 5224 23552 5408 23648 5 sr_0.FILLER_0_21_161.VPWR
flabel metal1 4977 23583 5011 23617 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_21_Right_21.VPWR
flabel metal1 4977 24127 5011 24161 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_21_Right_21.VGND
flabel nwell 4977 23583 5011 23617 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_21_Right_21.VPB
flabel pwell 4977 24127 5011 24161 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_21_Right_21.VNB
rlabel comment 4948 24144 4948 24144 2 sr_0.PHY_EDGE_ROW_21_Right_21.decap_3
rlabel metal1 4948 24096 5224 24192 5 sr_0.PHY_EDGE_ROW_21_Right_21.VGND
rlabel metal1 4948 23552 5224 23648 5 sr_0.PHY_EDGE_ROW_21_Right_21.VPWR
flabel metal1 19881 24127 19915 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_3.VGND
flabel metal1 19881 24671 19915 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_3.VPWR
flabel nwell 19881 24671 19915 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_3.VPB
flabel pwell 19881 24127 19915 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_3.VNB
rlabel comment 19944 24144 19944 24144 6 sr_0.FILLER_0_22_3.decap_12
flabel metal1 18777 24127 18811 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_15.VGND
flabel metal1 18777 24671 18811 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_15.VPWR
flabel nwell 18777 24671 18811 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_15.VPB
flabel pwell 18777 24127 18811 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_15.VNB
rlabel comment 18840 24144 18840 24144 6 sr_0.FILLER_0_22_15.decap_12
flabel metal1 20157 24671 20191 24705 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_22_Left_50.VPWR
flabel metal1 20157 24127 20191 24161 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_22_Left_50.VGND
flabel nwell 20157 24671 20191 24705 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_22_Left_50.VPB
flabel pwell 20157 24127 20191 24161 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_22_Left_50.VNB
rlabel comment 20220 24144 20220 24144 6 sr_0.PHY_EDGE_ROW_22_Left_50.decap_3
rlabel metal1 19944 24096 20220 24192 1 sr_0.PHY_EDGE_ROW_22_Left_50.VGND
rlabel metal1 19944 24640 20220 24736 1 sr_0.PHY_EDGE_ROW_22_Left_50.VPWR
flabel metal1 17678 24671 17714 24701 0 FreeSans 250 0 0 0 sr_0.FILLER_0_22_27.VPWR
flabel metal1 17678 24131 17714 24160 0 FreeSans 250 0 0 0 sr_0.FILLER_0_22_27.VGND
flabel nwell 17685 24678 17705 24695 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_27.VPB
flabel pwell 17684 24133 17708 24155 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_27.VNB
rlabel comment 17736 24144 17736 24144 6 sr_0.FILLER_0_22_27.fill_1
rlabel metal1 17644 24096 17736 24192 1 sr_0.FILLER_0_22_27.VGND
rlabel metal1 17644 24640 17736 24736 1 sr_0.FILLER_0_22_27.VPWR
flabel metal1 17489 24127 17523 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_29.VGND
flabel metal1 17489 24671 17523 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_29.VPWR
flabel nwell 17489 24671 17523 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_29.VPB
flabel pwell 17489 24127 17523 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_29.VNB
rlabel comment 17552 24144 17552 24144 6 sr_0.FILLER_0_22_29.decap_12
flabel metal1 16385 24127 16419 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_41.VGND
flabel metal1 16385 24671 16419 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_41.VPWR
flabel nwell 16385 24671 16419 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_41.VPB
flabel pwell 16385 24127 16419 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_41.VNB
rlabel comment 16448 24144 16448 24144 6 sr_0.FILLER_0_22_41.decap_12
flabel metal1 17569 24668 17622 24697 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_22_113.VPWR
flabel metal1 17572 24126 17623 24164 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_22_113.VGND
rlabel comment 17644 24144 17644 24144 6 sr_0.TAP_TAPCELL_ROW_22_113.tapvpwrvgnd_1
rlabel metal1 17552 24096 17644 24192 1 sr_0.TAP_TAPCELL_ROW_22_113.VGND
rlabel metal1 17552 24640 17644 24736 1 sr_0.TAP_TAPCELL_ROW_22_113.VPWR
flabel metal1 15281 24127 15315 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_53.VGND
flabel metal1 15281 24671 15315 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_53.VPWR
flabel nwell 15281 24671 15315 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_53.VPB
flabel pwell 15281 24127 15315 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_53.VNB
rlabel comment 15344 24144 15344 24144 6 sr_0.FILLER_0_22_53.decap_12
flabel metal1 14177 24127 14211 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_65.VGND
flabel metal1 14177 24671 14211 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_65.VPWR
flabel nwell 14177 24671 14211 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_65.VPB
flabel pwell 14177 24127 14211 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_65.VNB
rlabel comment 14240 24144 14240 24144 6 sr_0.FILLER_0_22_65.decap_12
flabel metal1 13073 24671 13107 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_77.VPWR
flabel metal1 13073 24127 13107 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_77.VGND
flabel nwell 13073 24671 13107 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_77.VPB
flabel pwell 13073 24127 13107 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_77.VNB
rlabel comment 13136 24144 13136 24144 6 sr_0.FILLER_0_22_77.decap_6
rlabel metal1 12584 24096 13136 24192 1 sr_0.FILLER_0_22_77.VGND
rlabel metal1 12584 24640 13136 24736 1 sr_0.FILLER_0_22_77.VPWR
flabel metal1 12526 24671 12562 24701 0 FreeSans 250 0 0 0 sr_0.FILLER_0_22_83.VPWR
flabel metal1 12526 24131 12562 24160 0 FreeSans 250 0 0 0 sr_0.FILLER_0_22_83.VGND
flabel nwell 12533 24678 12553 24695 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_83.VPB
flabel pwell 12532 24133 12556 24155 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_83.VNB
rlabel comment 12584 24144 12584 24144 6 sr_0.FILLER_0_22_83.fill_1
rlabel metal1 12492 24096 12584 24192 1 sr_0.FILLER_0_22_83.VGND
rlabel metal1 12492 24640 12584 24736 1 sr_0.FILLER_0_22_83.VPWR
flabel metal1 12337 24127 12371 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_85.VGND
flabel metal1 12337 24671 12371 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_85.VPWR
flabel nwell 12337 24671 12371 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_85.VPB
flabel pwell 12337 24127 12371 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_85.VNB
rlabel comment 12400 24144 12400 24144 6 sr_0.FILLER_0_22_85.decap_12
flabel metal1 11233 24127 11267 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_97.VGND
flabel metal1 11233 24671 11267 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_97.VPWR
flabel nwell 11233 24671 11267 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_97.VPB
flabel pwell 11233 24127 11267 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_97.VNB
rlabel comment 11296 24144 11296 24144 6 sr_0.FILLER_0_22_97.decap_12
flabel metal1 12417 24668 12470 24697 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_22_114.VPWR
flabel metal1 12420 24126 12471 24164 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_22_114.VGND
rlabel comment 12492 24144 12492 24144 6 sr_0.TAP_TAPCELL_ROW_22_114.tapvpwrvgnd_1
rlabel metal1 12400 24096 12492 24192 1 sr_0.TAP_TAPCELL_ROW_22_114.VGND
rlabel metal1 12400 24640 12492 24736 1 sr_0.TAP_TAPCELL_ROW_22_114.VPWR
flabel metal1 10129 24127 10163 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_109.VGND
flabel metal1 10129 24671 10163 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_109.VPWR
flabel nwell 10129 24671 10163 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_109.VPB
flabel pwell 10129 24127 10163 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_109.VNB
rlabel comment 10192 24144 10192 24144 6 sr_0.FILLER_0_22_109.decap_12
flabel metal1 9025 24127 9059 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_121.VGND
flabel metal1 9025 24671 9059 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_121.VPWR
flabel nwell 9025 24671 9059 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_121.VPB
flabel pwell 9025 24127 9059 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_121.VNB
rlabel comment 9088 24144 9088 24144 6 sr_0.FILLER_0_22_121.decap_12
flabel metal1 7921 24671 7955 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_133.VPWR
flabel metal1 7921 24127 7955 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_133.VGND
flabel nwell 7921 24671 7955 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_133.VPB
flabel pwell 7921 24127 7955 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_133.VNB
rlabel comment 7984 24144 7984 24144 6 sr_0.FILLER_0_22_133.decap_6
rlabel metal1 7432 24096 7984 24192 1 sr_0.FILLER_0_22_133.VGND
rlabel metal1 7432 24640 7984 24736 1 sr_0.FILLER_0_22_133.VPWR
flabel metal1 7374 24671 7410 24701 0 FreeSans 250 0 0 0 sr_0.FILLER_0_22_139.VPWR
flabel metal1 7374 24131 7410 24160 0 FreeSans 250 0 0 0 sr_0.FILLER_0_22_139.VGND
flabel nwell 7381 24678 7401 24695 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_139.VPB
flabel pwell 7380 24133 7404 24155 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_139.VNB
rlabel comment 7432 24144 7432 24144 6 sr_0.FILLER_0_22_139.fill_1
rlabel metal1 7340 24096 7432 24192 1 sr_0.FILLER_0_22_139.VGND
rlabel metal1 7340 24640 7432 24736 1 sr_0.FILLER_0_22_139.VPWR
flabel metal1 7185 24127 7219 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_141.VGND
flabel metal1 7185 24671 7219 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_141.VPWR
flabel nwell 7185 24671 7219 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_141.VPB
flabel pwell 7185 24127 7219 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_141.VNB
rlabel comment 7248 24144 7248 24144 6 sr_0.FILLER_0_22_141.decap_12
flabel metal1 7265 24668 7318 24697 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_22_115.VPWR
flabel metal1 7268 24126 7319 24164 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_22_115.VGND
rlabel comment 7340 24144 7340 24144 6 sr_0.TAP_TAPCELL_ROW_22_115.tapvpwrvgnd_1
rlabel metal1 7248 24096 7340 24192 1 sr_0.TAP_TAPCELL_ROW_22_115.VGND
rlabel metal1 7248 24640 7340 24736 1 sr_0.TAP_TAPCELL_ROW_22_115.VPWR
flabel metal1 6081 24671 6115 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_153.VPWR
flabel metal1 6081 24127 6115 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_153.VGND
flabel nwell 6081 24671 6115 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_153.VPB
flabel pwell 6081 24127 6115 24161 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_153.VNB
rlabel comment 6144 24144 6144 24144 6 sr_0.FILLER_0_22_153.decap_8
rlabel metal1 5408 24096 6144 24192 1 sr_0.FILLER_0_22_153.VGND
rlabel metal1 5408 24640 6144 24736 1 sr_0.FILLER_0_22_153.VPWR
flabel metal1 5335 24130 5388 24162 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_161.VGND
flabel metal1 5335 24674 5387 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_161.VPWR
flabel nwell 5346 24679 5380 24697 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_161.VPB
flabel pwell 5345 24134 5377 24156 0 FreeSans 200 0 0 0 sr_0.FILLER_0_22_161.VNB
rlabel comment 5408 24144 5408 24144 6 sr_0.FILLER_0_22_161.fill_2
rlabel metal1 5224 24096 5408 24192 1 sr_0.FILLER_0_22_161.VGND
rlabel metal1 5224 24640 5408 24736 1 sr_0.FILLER_0_22_161.VPWR
flabel metal1 4977 24671 5011 24705 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_22_Right_22.VPWR
flabel metal1 4977 24127 5011 24161 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_22_Right_22.VGND
flabel nwell 4977 24671 5011 24705 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_22_Right_22.VPB
flabel pwell 4977 24127 5011 24161 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_22_Right_22.VNB
rlabel comment 4948 24144 4948 24144 4 sr_0.PHY_EDGE_ROW_22_Right_22.decap_3
rlabel metal1 4948 24096 5224 24192 1 sr_0.PHY_EDGE_ROW_22_Right_22.VGND
rlabel metal1 4948 24640 5224 24736 1 sr_0.PHY_EDGE_ROW_22_Right_22.VPWR
flabel metal1 19881 25215 19915 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_3.VGND
flabel metal1 19881 24671 19915 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_3.VPWR
flabel nwell 19881 24671 19915 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_3.VPB
flabel pwell 19881 25215 19915 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_3.VNB
rlabel comment 19944 25232 19944 25232 8 sr_0.FILLER_0_23_3.decap_12
flabel metal1 18777 25215 18811 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_15.VGND
flabel metal1 18777 24671 18811 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_15.VPWR
flabel nwell 18777 24671 18811 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_15.VPB
flabel pwell 18777 25215 18811 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_15.VNB
rlabel comment 18840 25232 18840 25232 8 sr_0.FILLER_0_23_15.decap_12
flabel metal1 20157 24671 20191 24705 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_23_Left_51.VPWR
flabel metal1 20157 25215 20191 25249 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_23_Left_51.VGND
flabel nwell 20157 24671 20191 24705 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_23_Left_51.VPB
flabel pwell 20157 25215 20191 25249 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_23_Left_51.VNB
rlabel comment 20220 25232 20220 25232 8 sr_0.PHY_EDGE_ROW_23_Left_51.decap_3
rlabel metal1 19944 25184 20220 25280 5 sr_0.PHY_EDGE_ROW_23_Left_51.VGND
rlabel metal1 19944 24640 20220 24736 5 sr_0.PHY_EDGE_ROW_23_Left_51.VPWR
flabel metal1 17673 25215 17707 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_27.VGND
flabel metal1 17673 24671 17707 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_27.VPWR
flabel nwell 17673 24671 17707 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_27.VPB
flabel pwell 17673 25215 17707 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_27.VNB
rlabel comment 17736 25232 17736 25232 8 sr_0.FILLER_0_23_27.decap_12
flabel metal1 16569 25215 16603 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_39.VGND
flabel metal1 16569 24671 16603 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_39.VPWR
flabel nwell 16569 24671 16603 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_39.VPB
flabel pwell 16569 25215 16603 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_39.VNB
rlabel comment 16632 25232 16632 25232 8 sr_0.FILLER_0_23_39.decap_12
flabel metal1 15465 25215 15499 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_51.VGND
flabel metal1 15465 24671 15499 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_51.VPWR
flabel nwell 15465 24671 15499 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_51.VPB
flabel pwell 15465 25215 15499 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_51.VNB
rlabel comment 15528 25232 15528 25232 8 sr_0.FILLER_0_23_51.decap_4
rlabel metal1 15160 25184 15528 25280 5 sr_0.FILLER_0_23_51.VGND
rlabel metal1 15160 24640 15528 24736 5 sr_0.FILLER_0_23_51.VPWR
flabel metal1 15102 24675 15138 24705 0 FreeSans 250 0 0 0 sr_0.FILLER_0_23_55.VPWR
flabel metal1 15102 25216 15138 25245 0 FreeSans 250 0 0 0 sr_0.FILLER_0_23_55.VGND
flabel nwell 15109 24681 15129 24698 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_55.VPB
flabel pwell 15108 25221 15132 25243 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_55.VNB
rlabel comment 15160 25232 15160 25232 8 sr_0.FILLER_0_23_55.fill_1
rlabel metal1 15068 25184 15160 25280 5 sr_0.FILLER_0_23_55.VGND
rlabel metal1 15068 24640 15160 24736 5 sr_0.FILLER_0_23_55.VPWR
flabel metal1 14913 25215 14947 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_57.VGND
flabel metal1 14913 24671 14947 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_57.VPWR
flabel nwell 14913 24671 14947 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_57.VPB
flabel pwell 14913 25215 14947 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_57.VNB
rlabel comment 14976 25232 14976 25232 8 sr_0.FILLER_0_23_57.decap_12
flabel metal1 14993 24679 15046 24708 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_23_116.VPWR
flabel metal1 14996 25212 15047 25250 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_23_116.VGND
rlabel comment 15068 25232 15068 25232 8 sr_0.TAP_TAPCELL_ROW_23_116.tapvpwrvgnd_1
rlabel metal1 14976 25184 15068 25280 5 sr_0.TAP_TAPCELL_ROW_23_116.VGND
rlabel metal1 14976 24640 15068 24736 5 sr_0.TAP_TAPCELL_ROW_23_116.VPWR
flabel metal1 13809 25215 13843 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_69.VGND
flabel metal1 13809 24671 13843 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_69.VPWR
flabel nwell 13809 24671 13843 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_69.VPB
flabel pwell 13809 25215 13843 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_69.VNB
rlabel comment 13872 25232 13872 25232 8 sr_0.FILLER_0_23_69.decap_12
flabel metal1 12705 25215 12739 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_81.VGND
flabel metal1 12705 24671 12739 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_81.VPWR
flabel nwell 12705 24671 12739 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_81.VPB
flabel pwell 12705 25215 12739 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_81.VNB
rlabel comment 12768 25232 12768 25232 8 sr_0.FILLER_0_23_81.decap_12
flabel metal1 11601 25215 11635 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_93.VGND
flabel metal1 11601 24671 11635 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_93.VPWR
flabel nwell 11601 24671 11635 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_93.VPB
flabel pwell 11601 25215 11635 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_93.VNB
rlabel comment 11664 25232 11664 25232 8 sr_0.FILLER_0_23_93.decap_12
flabel metal1 10497 24671 10531 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_105.VPWR
flabel metal1 10497 25215 10531 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_105.VGND
flabel nwell 10497 24671 10531 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_105.VPB
flabel pwell 10497 25215 10531 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_105.VNB
rlabel comment 10560 25232 10560 25232 8 sr_0.FILLER_0_23_105.decap_6
rlabel metal1 10008 25184 10560 25280 5 sr_0.FILLER_0_23_105.VGND
rlabel metal1 10008 24640 10560 24736 5 sr_0.FILLER_0_23_105.VPWR
flabel metal1 9950 24675 9986 24705 0 FreeSans 250 0 0 0 sr_0.FILLER_0_23_111.VPWR
flabel metal1 9950 25216 9986 25245 0 FreeSans 250 0 0 0 sr_0.FILLER_0_23_111.VGND
flabel nwell 9957 24681 9977 24698 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_111.VPB
flabel pwell 9956 25221 9980 25243 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_111.VNB
rlabel comment 10008 25232 10008 25232 8 sr_0.FILLER_0_23_111.fill_1
rlabel metal1 9916 25184 10008 25280 5 sr_0.FILLER_0_23_111.VGND
rlabel metal1 9916 24640 10008 24736 5 sr_0.FILLER_0_23_111.VPWR
flabel metal1 9761 25215 9795 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_113.VGND
flabel metal1 9761 24671 9795 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_113.VPWR
flabel nwell 9761 24671 9795 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_113.VPB
flabel pwell 9761 25215 9795 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_113.VNB
rlabel comment 9824 25232 9824 25232 8 sr_0.FILLER_0_23_113.decap_12
flabel metal1 8657 25215 8691 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_125.VGND
flabel metal1 8657 24671 8691 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_125.VPWR
flabel nwell 8657 24671 8691 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_125.VPB
flabel pwell 8657 25215 8691 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_125.VNB
rlabel comment 8720 25232 8720 25232 8 sr_0.FILLER_0_23_125.decap_12
flabel metal1 9841 24679 9894 24708 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_23_117.VPWR
flabel metal1 9844 25212 9895 25250 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_23_117.VGND
rlabel comment 9916 25232 9916 25232 8 sr_0.TAP_TAPCELL_ROW_23_117.tapvpwrvgnd_1
rlabel metal1 9824 25184 9916 25280 5 sr_0.TAP_TAPCELL_ROW_23_117.VGND
rlabel metal1 9824 24640 9916 24736 5 sr_0.TAP_TAPCELL_ROW_23_117.VPWR
flabel metal1 7553 25215 7587 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_137.VGND
flabel metal1 7553 24671 7587 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_137.VPWR
flabel nwell 7553 24671 7587 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_137.VPB
flabel pwell 7553 25215 7587 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_137.VNB
rlabel comment 7616 25232 7616 25232 8 sr_0.FILLER_0_23_137.decap_12
flabel metal1 6449 25215 6483 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_149.VGND
flabel metal1 6449 24671 6483 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_149.VPWR
flabel nwell 6449 24671 6483 24705 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_149.VPB
flabel pwell 6449 25215 6483 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_149.VNB
rlabel comment 6512 25232 6512 25232 8 sr_0.FILLER_0_23_149.decap_12
flabel metal1 5335 25214 5388 25246 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_161.VGND
flabel metal1 5335 24671 5387 24702 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_161.VPWR
flabel nwell 5346 24679 5380 24697 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_161.VPB
flabel pwell 5345 25220 5377 25242 0 FreeSans 200 0 0 0 sr_0.FILLER_0_23_161.VNB
rlabel comment 5408 25232 5408 25232 8 sr_0.FILLER_0_23_161.fill_2
rlabel metal1 5224 25184 5408 25280 5 sr_0.FILLER_0_23_161.VGND
rlabel metal1 5224 24640 5408 24736 5 sr_0.FILLER_0_23_161.VPWR
flabel metal1 4977 24671 5011 24705 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_23_Right_23.VPWR
flabel metal1 4977 25215 5011 25249 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_23_Right_23.VGND
flabel nwell 4977 24671 5011 24705 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_23_Right_23.VPB
flabel pwell 4977 25215 5011 25249 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_23_Right_23.VNB
rlabel comment 4948 25232 4948 25232 2 sr_0.PHY_EDGE_ROW_23_Right_23.decap_3
rlabel metal1 4948 25184 5224 25280 5 sr_0.PHY_EDGE_ROW_23_Right_23.VGND
rlabel metal1 4948 24640 5224 24736 5 sr_0.PHY_EDGE_ROW_23_Right_23.VPWR
flabel metal1 19881 25215 19915 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_3.VGND
flabel metal1 19881 25759 19915 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_3.VPWR
flabel nwell 19881 25759 19915 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_3.VPB
flabel pwell 19881 25215 19915 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_3.VNB
rlabel comment 19944 25232 19944 25232 6 sr_0.FILLER_0_24_3.decap_12
flabel metal1 18777 25215 18811 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_15.VGND
flabel metal1 18777 25759 18811 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_15.VPWR
flabel nwell 18777 25759 18811 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_15.VPB
flabel pwell 18777 25215 18811 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_15.VNB
rlabel comment 18840 25232 18840 25232 6 sr_0.FILLER_0_24_15.decap_12
flabel metal1 20157 25759 20191 25793 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_24_Left_52.VPWR
flabel metal1 20157 25215 20191 25249 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_24_Left_52.VGND
flabel nwell 20157 25759 20191 25793 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_24_Left_52.VPB
flabel pwell 20157 25215 20191 25249 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_24_Left_52.VNB
rlabel comment 20220 25232 20220 25232 6 sr_0.PHY_EDGE_ROW_24_Left_52.decap_3
rlabel metal1 19944 25184 20220 25280 1 sr_0.PHY_EDGE_ROW_24_Left_52.VGND
rlabel metal1 19944 25728 20220 25824 1 sr_0.PHY_EDGE_ROW_24_Left_52.VPWR
flabel metal1 17678 25759 17714 25789 0 FreeSans 250 0 0 0 sr_0.FILLER_0_24_27.VPWR
flabel metal1 17678 25219 17714 25248 0 FreeSans 250 0 0 0 sr_0.FILLER_0_24_27.VGND
flabel nwell 17685 25766 17705 25783 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_27.VPB
flabel pwell 17684 25221 17708 25243 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_27.VNB
rlabel comment 17736 25232 17736 25232 6 sr_0.FILLER_0_24_27.fill_1
rlabel metal1 17644 25184 17736 25280 1 sr_0.FILLER_0_24_27.VGND
rlabel metal1 17644 25728 17736 25824 1 sr_0.FILLER_0_24_27.VPWR
flabel metal1 17489 25215 17523 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_29.VGND
flabel metal1 17489 25759 17523 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_29.VPWR
flabel nwell 17489 25759 17523 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_29.VPB
flabel pwell 17489 25215 17523 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_29.VNB
rlabel comment 17552 25232 17552 25232 6 sr_0.FILLER_0_24_29.decap_12
flabel metal1 16385 25215 16419 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_41.VGND
flabel metal1 16385 25759 16419 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_41.VPWR
flabel nwell 16385 25759 16419 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_41.VPB
flabel pwell 16385 25215 16419 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_41.VNB
rlabel comment 16448 25232 16448 25232 6 sr_0.FILLER_0_24_41.decap_12
flabel metal1 17569 25756 17622 25785 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_24_118.VPWR
flabel metal1 17572 25214 17623 25252 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_24_118.VGND
rlabel comment 17644 25232 17644 25232 6 sr_0.TAP_TAPCELL_ROW_24_118.tapvpwrvgnd_1
rlabel metal1 17552 25184 17644 25280 1 sr_0.TAP_TAPCELL_ROW_24_118.VGND
rlabel metal1 17552 25728 17644 25824 1 sr_0.TAP_TAPCELL_ROW_24_118.VPWR
flabel metal1 15281 25215 15315 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_53.VGND
flabel metal1 15281 25759 15315 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_53.VPWR
flabel nwell 15281 25759 15315 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_53.VPB
flabel pwell 15281 25215 15315 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_53.VNB
rlabel comment 15344 25232 15344 25232 6 sr_0.FILLER_0_24_53.decap_12
flabel metal1 14177 25215 14211 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_65.VGND
flabel metal1 14177 25759 14211 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_65.VPWR
flabel nwell 14177 25759 14211 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_65.VPB
flabel pwell 14177 25215 14211 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_65.VNB
rlabel comment 14240 25232 14240 25232 6 sr_0.FILLER_0_24_65.decap_12
flabel metal1 13073 25759 13107 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_77.VPWR
flabel metal1 13073 25215 13107 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_77.VGND
flabel nwell 13073 25759 13107 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_77.VPB
flabel pwell 13073 25215 13107 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_77.VNB
rlabel comment 13136 25232 13136 25232 6 sr_0.FILLER_0_24_77.decap_6
rlabel metal1 12584 25184 13136 25280 1 sr_0.FILLER_0_24_77.VGND
rlabel metal1 12584 25728 13136 25824 1 sr_0.FILLER_0_24_77.VPWR
flabel metal1 12526 25759 12562 25789 0 FreeSans 250 0 0 0 sr_0.FILLER_0_24_83.VPWR
flabel metal1 12526 25219 12562 25248 0 FreeSans 250 0 0 0 sr_0.FILLER_0_24_83.VGND
flabel nwell 12533 25766 12553 25783 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_83.VPB
flabel pwell 12532 25221 12556 25243 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_83.VNB
rlabel comment 12584 25232 12584 25232 6 sr_0.FILLER_0_24_83.fill_1
rlabel metal1 12492 25184 12584 25280 1 sr_0.FILLER_0_24_83.VGND
rlabel metal1 12492 25728 12584 25824 1 sr_0.FILLER_0_24_83.VPWR
flabel metal1 12337 25215 12371 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_85.VGND
flabel metal1 12337 25759 12371 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_85.VPWR
flabel nwell 12337 25759 12371 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_85.VPB
flabel pwell 12337 25215 12371 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_85.VNB
rlabel comment 12400 25232 12400 25232 6 sr_0.FILLER_0_24_85.decap_12
flabel metal1 11233 25215 11267 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_97.VGND
flabel metal1 11233 25759 11267 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_97.VPWR
flabel nwell 11233 25759 11267 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_97.VPB
flabel pwell 11233 25215 11267 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_97.VNB
rlabel comment 11296 25232 11296 25232 6 sr_0.FILLER_0_24_97.decap_12
flabel metal1 12417 25756 12470 25785 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_24_119.VPWR
flabel metal1 12420 25214 12471 25252 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_24_119.VGND
rlabel comment 12492 25232 12492 25232 6 sr_0.TAP_TAPCELL_ROW_24_119.tapvpwrvgnd_1
rlabel metal1 12400 25184 12492 25280 1 sr_0.TAP_TAPCELL_ROW_24_119.VGND
rlabel metal1 12400 25728 12492 25824 1 sr_0.TAP_TAPCELL_ROW_24_119.VPWR
flabel metal1 10129 25215 10163 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_109.VGND
flabel metal1 10129 25759 10163 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_109.VPWR
flabel nwell 10129 25759 10163 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_109.VPB
flabel pwell 10129 25215 10163 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_109.VNB
rlabel comment 10192 25232 10192 25232 6 sr_0.FILLER_0_24_109.decap_12
flabel metal1 9025 25215 9059 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_121.VGND
flabel metal1 9025 25759 9059 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_121.VPWR
flabel nwell 9025 25759 9059 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_121.VPB
flabel pwell 9025 25215 9059 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_121.VNB
rlabel comment 9088 25232 9088 25232 6 sr_0.FILLER_0_24_121.decap_12
flabel metal1 7921 25759 7955 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_133.VPWR
flabel metal1 7921 25215 7955 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_133.VGND
flabel nwell 7921 25759 7955 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_133.VPB
flabel pwell 7921 25215 7955 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_133.VNB
rlabel comment 7984 25232 7984 25232 6 sr_0.FILLER_0_24_133.decap_6
rlabel metal1 7432 25184 7984 25280 1 sr_0.FILLER_0_24_133.VGND
rlabel metal1 7432 25728 7984 25824 1 sr_0.FILLER_0_24_133.VPWR
flabel metal1 7374 25759 7410 25789 0 FreeSans 250 0 0 0 sr_0.FILLER_0_24_139.VPWR
flabel metal1 7374 25219 7410 25248 0 FreeSans 250 0 0 0 sr_0.FILLER_0_24_139.VGND
flabel nwell 7381 25766 7401 25783 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_139.VPB
flabel pwell 7380 25221 7404 25243 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_139.VNB
rlabel comment 7432 25232 7432 25232 6 sr_0.FILLER_0_24_139.fill_1
rlabel metal1 7340 25184 7432 25280 1 sr_0.FILLER_0_24_139.VGND
rlabel metal1 7340 25728 7432 25824 1 sr_0.FILLER_0_24_139.VPWR
flabel metal1 7185 25215 7219 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_141.VGND
flabel metal1 7185 25759 7219 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_141.VPWR
flabel nwell 7185 25759 7219 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_141.VPB
flabel pwell 7185 25215 7219 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_141.VNB
rlabel comment 7248 25232 7248 25232 6 sr_0.FILLER_0_24_141.decap_12
flabel metal1 7265 25756 7318 25785 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_24_120.VPWR
flabel metal1 7268 25214 7319 25252 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_24_120.VGND
rlabel comment 7340 25232 7340 25232 6 sr_0.TAP_TAPCELL_ROW_24_120.tapvpwrvgnd_1
rlabel metal1 7248 25184 7340 25280 1 sr_0.TAP_TAPCELL_ROW_24_120.VGND
rlabel metal1 7248 25728 7340 25824 1 sr_0.TAP_TAPCELL_ROW_24_120.VPWR
flabel metal1 6081 25759 6115 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_153.VPWR
flabel metal1 6081 25215 6115 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_153.VGND
flabel nwell 6081 25759 6115 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_153.VPB
flabel pwell 6081 25215 6115 25249 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_153.VNB
rlabel comment 6144 25232 6144 25232 6 sr_0.FILLER_0_24_153.decap_8
rlabel metal1 5408 25184 6144 25280 1 sr_0.FILLER_0_24_153.VGND
rlabel metal1 5408 25728 6144 25824 1 sr_0.FILLER_0_24_153.VPWR
flabel metal1 5335 25218 5388 25250 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_161.VGND
flabel metal1 5335 25762 5387 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_161.VPWR
flabel nwell 5346 25767 5380 25785 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_161.VPB
flabel pwell 5345 25222 5377 25244 0 FreeSans 200 0 0 0 sr_0.FILLER_0_24_161.VNB
rlabel comment 5408 25232 5408 25232 6 sr_0.FILLER_0_24_161.fill_2
rlabel metal1 5224 25184 5408 25280 1 sr_0.FILLER_0_24_161.VGND
rlabel metal1 5224 25728 5408 25824 1 sr_0.FILLER_0_24_161.VPWR
flabel metal1 4977 25759 5011 25793 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_24_Right_24.VPWR
flabel metal1 4977 25215 5011 25249 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_24_Right_24.VGND
flabel nwell 4977 25759 5011 25793 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_24_Right_24.VPB
flabel pwell 4977 25215 5011 25249 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_24_Right_24.VNB
rlabel comment 4948 25232 4948 25232 4 sr_0.PHY_EDGE_ROW_24_Right_24.decap_3
rlabel metal1 4948 25184 5224 25280 1 sr_0.PHY_EDGE_ROW_24_Right_24.VGND
rlabel metal1 4948 25728 5224 25824 1 sr_0.PHY_EDGE_ROW_24_Right_24.VPWR
flabel metal1 19881 26303 19915 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_3.VGND
flabel metal1 19881 25759 19915 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_3.VPWR
flabel nwell 19881 25759 19915 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_3.VPB
flabel pwell 19881 26303 19915 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_3.VNB
rlabel comment 19944 26320 19944 26320 8 sr_0.FILLER_0_25_3.decap_12
flabel metal1 18777 26303 18811 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_15.VGND
flabel metal1 18777 25759 18811 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_15.VPWR
flabel nwell 18777 25759 18811 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_15.VPB
flabel pwell 18777 26303 18811 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_15.VNB
rlabel comment 18840 26320 18840 26320 8 sr_0.FILLER_0_25_15.decap_12
flabel metal1 20157 25759 20191 25793 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_25_Left_53.VPWR
flabel metal1 20157 26303 20191 26337 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_25_Left_53.VGND
flabel nwell 20157 25759 20191 25793 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_25_Left_53.VPB
flabel pwell 20157 26303 20191 26337 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_25_Left_53.VNB
rlabel comment 20220 26320 20220 26320 8 sr_0.PHY_EDGE_ROW_25_Left_53.decap_3
rlabel metal1 19944 26272 20220 26368 5 sr_0.PHY_EDGE_ROW_25_Left_53.VGND
rlabel metal1 19944 25728 20220 25824 5 sr_0.PHY_EDGE_ROW_25_Left_53.VPWR
flabel metal1 17673 26303 17707 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_27.VGND
flabel metal1 17673 25759 17707 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_27.VPWR
flabel nwell 17673 25759 17707 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_27.VPB
flabel pwell 17673 26303 17707 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_27.VNB
rlabel comment 17736 26320 17736 26320 8 sr_0.FILLER_0_25_27.decap_12
flabel metal1 16569 26303 16603 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_39.VGND
flabel metal1 16569 25759 16603 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_39.VPWR
flabel nwell 16569 25759 16603 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_39.VPB
flabel pwell 16569 26303 16603 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_39.VNB
rlabel comment 16632 26320 16632 26320 8 sr_0.FILLER_0_25_39.decap_12
flabel metal1 15465 26303 15499 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_51.VGND
flabel metal1 15465 25759 15499 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_51.VPWR
flabel nwell 15465 25759 15499 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_51.VPB
flabel pwell 15465 26303 15499 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_51.VNB
rlabel comment 15528 26320 15528 26320 8 sr_0.FILLER_0_25_51.decap_4
rlabel metal1 15160 26272 15528 26368 5 sr_0.FILLER_0_25_51.VGND
rlabel metal1 15160 25728 15528 25824 5 sr_0.FILLER_0_25_51.VPWR
flabel metal1 15102 25763 15138 25793 0 FreeSans 250 0 0 0 sr_0.FILLER_0_25_55.VPWR
flabel metal1 15102 26304 15138 26333 0 FreeSans 250 0 0 0 sr_0.FILLER_0_25_55.VGND
flabel nwell 15109 25769 15129 25786 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_55.VPB
flabel pwell 15108 26309 15132 26331 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_55.VNB
rlabel comment 15160 26320 15160 26320 8 sr_0.FILLER_0_25_55.fill_1
rlabel metal1 15068 26272 15160 26368 5 sr_0.FILLER_0_25_55.VGND
rlabel metal1 15068 25728 15160 25824 5 sr_0.FILLER_0_25_55.VPWR
flabel metal1 14913 26303 14947 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_57.VGND
flabel metal1 14913 25759 14947 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_57.VPWR
flabel nwell 14913 25759 14947 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_57.VPB
flabel pwell 14913 26303 14947 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_57.VNB
rlabel comment 14976 26320 14976 26320 8 sr_0.FILLER_0_25_57.decap_12
flabel metal1 14993 25767 15046 25796 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_25_121.VPWR
flabel metal1 14996 26300 15047 26338 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_25_121.VGND
rlabel comment 15068 26320 15068 26320 8 sr_0.TAP_TAPCELL_ROW_25_121.tapvpwrvgnd_1
rlabel metal1 14976 26272 15068 26368 5 sr_0.TAP_TAPCELL_ROW_25_121.VGND
rlabel metal1 14976 25728 15068 25824 5 sr_0.TAP_TAPCELL_ROW_25_121.VPWR
flabel metal1 13809 26303 13843 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_69.VGND
flabel metal1 13809 25759 13843 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_69.VPWR
flabel nwell 13809 25759 13843 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_69.VPB
flabel pwell 13809 26303 13843 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_69.VNB
rlabel comment 13872 26320 13872 26320 8 sr_0.FILLER_0_25_69.decap_12
flabel metal1 12705 26303 12739 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_81.VGND
flabel metal1 12705 25759 12739 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_81.VPWR
flabel nwell 12705 25759 12739 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_81.VPB
flabel pwell 12705 26303 12739 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_81.VNB
rlabel comment 12768 26320 12768 26320 8 sr_0.FILLER_0_25_81.decap_12
flabel metal1 11601 26303 11635 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_93.VGND
flabel metal1 11601 25759 11635 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_93.VPWR
flabel nwell 11601 25759 11635 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_93.VPB
flabel pwell 11601 26303 11635 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_93.VNB
rlabel comment 11664 26320 11664 26320 8 sr_0.FILLER_0_25_93.decap_12
flabel metal1 10497 25759 10531 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_105.VPWR
flabel metal1 10497 26303 10531 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_105.VGND
flabel nwell 10497 25759 10531 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_105.VPB
flabel pwell 10497 26303 10531 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_105.VNB
rlabel comment 10560 26320 10560 26320 8 sr_0.FILLER_0_25_105.decap_6
rlabel metal1 10008 26272 10560 26368 5 sr_0.FILLER_0_25_105.VGND
rlabel metal1 10008 25728 10560 25824 5 sr_0.FILLER_0_25_105.VPWR
flabel metal1 9950 25763 9986 25793 0 FreeSans 250 0 0 0 sr_0.FILLER_0_25_111.VPWR
flabel metal1 9950 26304 9986 26333 0 FreeSans 250 0 0 0 sr_0.FILLER_0_25_111.VGND
flabel nwell 9957 25769 9977 25786 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_111.VPB
flabel pwell 9956 26309 9980 26331 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_111.VNB
rlabel comment 10008 26320 10008 26320 8 sr_0.FILLER_0_25_111.fill_1
rlabel metal1 9916 26272 10008 26368 5 sr_0.FILLER_0_25_111.VGND
rlabel metal1 9916 25728 10008 25824 5 sr_0.FILLER_0_25_111.VPWR
flabel metal1 9761 26303 9795 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_113.VGND
flabel metal1 9761 25759 9795 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_113.VPWR
flabel nwell 9761 25759 9795 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_113.VPB
flabel pwell 9761 26303 9795 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_113.VNB
rlabel comment 9824 26320 9824 26320 8 sr_0.FILLER_0_25_113.decap_12
flabel metal1 8657 26303 8691 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_125.VGND
flabel metal1 8657 25759 8691 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_125.VPWR
flabel nwell 8657 25759 8691 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_125.VPB
flabel pwell 8657 26303 8691 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_125.VNB
rlabel comment 8720 26320 8720 26320 8 sr_0.FILLER_0_25_125.decap_12
flabel metal1 9841 25767 9894 25796 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_25_122.VPWR
flabel metal1 9844 26300 9895 26338 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_25_122.VGND
rlabel comment 9916 26320 9916 26320 8 sr_0.TAP_TAPCELL_ROW_25_122.tapvpwrvgnd_1
rlabel metal1 9824 26272 9916 26368 5 sr_0.TAP_TAPCELL_ROW_25_122.VGND
rlabel metal1 9824 25728 9916 25824 5 sr_0.TAP_TAPCELL_ROW_25_122.VPWR
flabel metal1 7553 26303 7587 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_137.VGND
flabel metal1 7553 25759 7587 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_137.VPWR
flabel nwell 7553 25759 7587 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_137.VPB
flabel pwell 7553 26303 7587 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_137.VNB
rlabel comment 7616 26320 7616 26320 8 sr_0.FILLER_0_25_137.decap_12
flabel metal1 6449 26303 6483 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_149.VGND
flabel metal1 6449 25759 6483 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_149.VPWR
flabel nwell 6449 25759 6483 25793 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_149.VPB
flabel pwell 6449 26303 6483 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_149.VNB
rlabel comment 6512 26320 6512 26320 8 sr_0.FILLER_0_25_149.decap_12
flabel metal1 5335 26302 5388 26334 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_161.VGND
flabel metal1 5335 25759 5387 25790 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_161.VPWR
flabel nwell 5346 25767 5380 25785 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_161.VPB
flabel pwell 5345 26308 5377 26330 0 FreeSans 200 0 0 0 sr_0.FILLER_0_25_161.VNB
rlabel comment 5408 26320 5408 26320 8 sr_0.FILLER_0_25_161.fill_2
rlabel metal1 5224 26272 5408 26368 5 sr_0.FILLER_0_25_161.VGND
rlabel metal1 5224 25728 5408 25824 5 sr_0.FILLER_0_25_161.VPWR
flabel metal1 4977 25759 5011 25793 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_25_Right_25.VPWR
flabel metal1 4977 26303 5011 26337 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_25_Right_25.VGND
flabel nwell 4977 25759 5011 25793 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_25_Right_25.VPB
flabel pwell 4977 26303 5011 26337 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_25_Right_25.VNB
rlabel comment 4948 26320 4948 26320 2 sr_0.PHY_EDGE_ROW_25_Right_25.decap_3
rlabel metal1 4948 26272 5224 26368 5 sr_0.PHY_EDGE_ROW_25_Right_25.VGND
rlabel metal1 4948 25728 5224 25824 5 sr_0.PHY_EDGE_ROW_25_Right_25.VPWR
flabel metal1 19881 26303 19915 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_3.VGND
flabel metal1 19881 26847 19915 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_3.VPWR
flabel nwell 19881 26847 19915 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_3.VPB
flabel pwell 19881 26303 19915 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_3.VNB
rlabel comment 19944 26320 19944 26320 6 sr_0.FILLER_0_26_3.decap_12
flabel metal1 18777 26303 18811 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_15.VGND
flabel metal1 18777 26847 18811 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_15.VPWR
flabel nwell 18777 26847 18811 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_15.VPB
flabel pwell 18777 26303 18811 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_15.VNB
rlabel comment 18840 26320 18840 26320 6 sr_0.FILLER_0_26_15.decap_12
flabel metal1 19881 26847 19915 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_3.VPWR
flabel metal1 19881 27391 19915 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_3.VGND
flabel nwell 19881 26847 19915 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_3.VPB
flabel pwell 19881 27391 19915 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_3.VNB
rlabel comment 19944 27408 19944 27408 8 sr_0.FILLER_0_27_3.decap_8
rlabel metal1 19208 27360 19944 27456 5 sr_0.FILLER_0_27_3.VGND
rlabel metal1 19208 26816 19944 26912 5 sr_0.FILLER_0_27_3.VPWR
flabel metal1 19135 27390 19188 27422 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_11.VGND
flabel metal1 19135 26847 19187 26878 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_11.VPWR
flabel nwell 19146 26855 19180 26873 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_11.VPB
flabel pwell 19145 27396 19177 27418 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_11.VNB
rlabel comment 19208 27408 19208 27408 8 sr_0.FILLER_0_27_11.fill_2
rlabel metal1 19024 27360 19208 27456 5 sr_0.FILLER_0_27_11.VGND
rlabel metal1 19024 26816 19208 26912 5 sr_0.FILLER_0_27_11.VPWR
flabel metal1 18409 26847 18443 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_19.VPWR
flabel metal1 18409 27391 18443 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_19.VGND
flabel nwell 18409 26847 18443 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_19.VPB
flabel pwell 18409 27391 18443 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_19.VNB
rlabel comment 18472 27408 18472 27408 8 sr_0.FILLER_0_27_19.decap_8
rlabel metal1 17736 27360 18472 27456 5 sr_0.FILLER_0_27_19.VGND
rlabel metal1 17736 26816 18472 26912 5 sr_0.FILLER_0_27_19.VPWR
flabel metal1 20157 26847 20191 26881 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_26_Left_54.VPWR
flabel metal1 20157 26303 20191 26337 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_26_Left_54.VGND
flabel nwell 20157 26847 20191 26881 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_26_Left_54.VPB
flabel pwell 20157 26303 20191 26337 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_26_Left_54.VNB
rlabel comment 20220 26320 20220 26320 6 sr_0.PHY_EDGE_ROW_26_Left_54.decap_3
rlabel metal1 19944 26272 20220 26368 1 sr_0.PHY_EDGE_ROW_26_Left_54.VGND
rlabel metal1 19944 26816 20220 26912 1 sr_0.PHY_EDGE_ROW_26_Left_54.VPWR
flabel metal1 20157 26847 20191 26881 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_27_Left_55.VPWR
flabel metal1 20157 27391 20191 27425 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_27_Left_55.VGND
flabel nwell 20157 26847 20191 26881 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_27_Left_55.VPB
flabel pwell 20157 27391 20191 27425 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_27_Left_55.VNB
rlabel comment 20220 27408 20220 27408 8 sr_0.PHY_EDGE_ROW_27_Left_55.decap_3
rlabel metal1 19944 27360 20220 27456 5 sr_0.PHY_EDGE_ROW_27_Left_55.VGND
rlabel metal1 19944 26816 20220 26912 5 sr_0.PHY_EDGE_ROW_27_Left_55.VPWR
flabel locali 18593 27085 18627 27119 0 FreeSans 200 0 0 0 sr_0.input3.X
flabel locali 18869 27221 18903 27255 0 FreeSans 200 0 0 0 sr_0.input3.A
flabel locali 18501 27221 18535 27255 0 FreeSans 200 0 0 0 sr_0.input3.X
flabel locali 18869 27153 18903 27187 0 FreeSans 200 0 0 0 sr_0.input3.A
flabel locali 18501 27153 18535 27187 0 FreeSans 200 0 0 0 sr_0.input3.X
flabel metal1 18961 27391 18995 27425 0 FreeSans 200 0 0 0 sr_0.input3.VGND
flabel metal1 18961 26847 18995 26881 0 FreeSans 200 0 0 0 sr_0.input3.VPWR
flabel nwell 18961 26847 18995 26881 0 FreeSans 200 0 0 0 sr_0.input3.VPB
flabel pwell 18961 27391 18995 27425 0 FreeSans 200 0 0 0 sr_0.input3.VNB
rlabel comment 19024 27408 19024 27408 8 sr_0.input3.clkbuf_4
rlabel metal1 18472 27360 19024 27456 5 sr_0.input3.VGND
rlabel metal1 18472 26816 19024 26912 5 sr_0.input3.VPWR
flabel metal1 17678 26847 17714 26877 0 FreeSans 250 0 0 0 sr_0.FILLER_0_26_27.VPWR
flabel metal1 17678 26307 17714 26336 0 FreeSans 250 0 0 0 sr_0.FILLER_0_26_27.VGND
flabel nwell 17685 26854 17705 26871 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_27.VPB
flabel pwell 17684 26309 17708 26331 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_27.VNB
rlabel comment 17736 26320 17736 26320 6 sr_0.FILLER_0_26_27.fill_1
rlabel metal1 17644 26272 17736 26368 1 sr_0.FILLER_0_26_27.VGND
rlabel metal1 17644 26816 17736 26912 1 sr_0.FILLER_0_26_27.VPWR
flabel metal1 17489 26303 17523 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_29.VGND
flabel metal1 17489 26847 17523 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_29.VPWR
flabel nwell 17489 26847 17523 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_29.VPB
flabel pwell 17489 26303 17523 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_29.VNB
rlabel comment 17552 26320 17552 26320 6 sr_0.FILLER_0_26_29.decap_12
flabel metal1 16385 26303 16419 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_41.VGND
flabel metal1 16385 26847 16419 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_41.VPWR
flabel nwell 16385 26847 16419 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_41.VPB
flabel pwell 16385 26303 16419 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_41.VNB
rlabel comment 16448 26320 16448 26320 6 sr_0.FILLER_0_26_41.decap_12
flabel metal1 17678 26851 17714 26881 0 FreeSans 250 0 0 0 sr_0.FILLER_0_27_27.VPWR
flabel metal1 17678 27392 17714 27421 0 FreeSans 250 0 0 0 sr_0.FILLER_0_27_27.VGND
flabel nwell 17685 26857 17705 26874 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_27.VPB
flabel pwell 17684 27397 17708 27419 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_27.VNB
rlabel comment 17736 27408 17736 27408 8 sr_0.FILLER_0_27_27.fill_1
rlabel metal1 17644 27360 17736 27456 5 sr_0.FILLER_0_27_27.VGND
rlabel metal1 17644 26816 17736 26912 5 sr_0.FILLER_0_27_27.VPWR
flabel metal1 17489 27391 17523 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_29.VGND
flabel metal1 17489 26847 17523 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_29.VPWR
flabel nwell 17489 26847 17523 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_29.VPB
flabel pwell 17489 27391 17523 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_29.VNB
rlabel comment 17552 27408 17552 27408 8 sr_0.FILLER_0_27_29.decap_12
flabel metal1 16385 27391 16419 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_41.VGND
flabel metal1 16385 26847 16419 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_41.VPWR
flabel nwell 16385 26847 16419 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_41.VPB
flabel pwell 16385 27391 16419 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_41.VNB
rlabel comment 16448 27408 16448 27408 8 sr_0.FILLER_0_27_41.decap_12
flabel metal1 17569 26844 17622 26873 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_26_123.VPWR
flabel metal1 17572 26302 17623 26340 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_26_123.VGND
rlabel comment 17644 26320 17644 26320 6 sr_0.TAP_TAPCELL_ROW_26_123.tapvpwrvgnd_1
rlabel metal1 17552 26272 17644 26368 1 sr_0.TAP_TAPCELL_ROW_26_123.VGND
rlabel metal1 17552 26816 17644 26912 1 sr_0.TAP_TAPCELL_ROW_26_123.VPWR
flabel metal1 17569 26855 17622 26884 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_27_126.VPWR
flabel metal1 17572 27388 17623 27426 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_27_126.VGND
rlabel comment 17644 27408 17644 27408 8 sr_0.TAP_TAPCELL_ROW_27_126.tapvpwrvgnd_1
rlabel metal1 17552 27360 17644 27456 5 sr_0.TAP_TAPCELL_ROW_27_126.VGND
rlabel metal1 17552 26816 17644 26912 5 sr_0.TAP_TAPCELL_ROW_27_126.VPWR
flabel metal1 15281 26303 15315 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_53.VGND
flabel metal1 15281 26847 15315 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_53.VPWR
flabel nwell 15281 26847 15315 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_53.VPB
flabel pwell 15281 26303 15315 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_53.VNB
rlabel comment 15344 26320 15344 26320 6 sr_0.FILLER_0_26_53.decap_12
flabel metal1 15281 26847 15315 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_53.VPWR
flabel metal1 15281 27391 15315 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_53.VGND
flabel nwell 15281 26847 15315 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_53.VPB
flabel pwell 15281 27391 15315 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_53.VNB
rlabel comment 15344 27408 15344 27408 8 sr_0.FILLER_0_27_53.decap_3
rlabel metal1 15068 27360 15344 27456 5 sr_0.FILLER_0_27_53.VGND
rlabel metal1 15068 26816 15344 26912 5 sr_0.FILLER_0_27_53.VPWR
flabel metal1 14913 27391 14947 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_57.VGND
flabel metal1 14913 26847 14947 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_57.VPWR
flabel nwell 14913 26847 14947 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_57.VPB
flabel pwell 14913 27391 14947 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_57.VNB
rlabel comment 14976 27408 14976 27408 8 sr_0.FILLER_0_27_57.decap_12
flabel metal1 14993 26855 15046 26884 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_27_127.VPWR
flabel metal1 14996 27388 15047 27426 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_27_127.VGND
rlabel comment 15068 27408 15068 27408 8 sr_0.TAP_TAPCELL_ROW_27_127.tapvpwrvgnd_1
rlabel metal1 14976 27360 15068 27456 5 sr_0.TAP_TAPCELL_ROW_27_127.VGND
rlabel metal1 14976 26816 15068 26912 5 sr_0.TAP_TAPCELL_ROW_27_127.VPWR
flabel metal1 14177 26303 14211 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_65.VGND
flabel metal1 14177 26847 14211 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_65.VPWR
flabel nwell 14177 26847 14211 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_65.VPB
flabel pwell 14177 26303 14211 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_65.VNB
rlabel comment 14240 26320 14240 26320 6 sr_0.FILLER_0_26_65.decap_12
flabel metal1 13073 26847 13107 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_77.VPWR
flabel metal1 13073 26303 13107 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_77.VGND
flabel nwell 13073 26847 13107 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_77.VPB
flabel pwell 13073 26303 13107 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_77.VNB
rlabel comment 13136 26320 13136 26320 6 sr_0.FILLER_0_26_77.decap_6
rlabel metal1 12584 26272 13136 26368 1 sr_0.FILLER_0_26_77.VGND
rlabel metal1 12584 26816 13136 26912 1 sr_0.FILLER_0_26_77.VPWR
flabel metal1 12526 26847 12562 26877 0 FreeSans 250 0 0 0 sr_0.FILLER_0_26_83.VPWR
flabel metal1 12526 26307 12562 26336 0 FreeSans 250 0 0 0 sr_0.FILLER_0_26_83.VGND
flabel nwell 12533 26854 12553 26871 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_83.VPB
flabel pwell 12532 26309 12556 26331 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_83.VNB
rlabel comment 12584 26320 12584 26320 6 sr_0.FILLER_0_26_83.fill_1
rlabel metal1 12492 26272 12584 26368 1 sr_0.FILLER_0_26_83.VGND
rlabel metal1 12492 26816 12584 26912 1 sr_0.FILLER_0_26_83.VPWR
flabel metal1 13809 27391 13843 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_69.VGND
flabel metal1 13809 26847 13843 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_69.VPWR
flabel nwell 13809 26847 13843 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_69.VPB
flabel pwell 13809 27391 13843 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_69.VNB
rlabel comment 13872 27408 13872 27408 8 sr_0.FILLER_0_27_69.decap_12
flabel metal1 12705 26847 12739 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_81.VPWR
flabel metal1 12705 27391 12739 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_81.VGND
flabel nwell 12705 26847 12739 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_81.VPB
flabel pwell 12705 27391 12739 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_81.VNB
rlabel comment 12768 27408 12768 27408 8 sr_0.FILLER_0_27_81.decap_3
rlabel metal1 12492 27360 12768 27456 5 sr_0.FILLER_0_27_81.VGND
rlabel metal1 12492 26816 12768 26912 5 sr_0.FILLER_0_27_81.VPWR
flabel metal1 12337 26303 12371 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_85.VGND
flabel metal1 12337 26847 12371 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_85.VPWR
flabel nwell 12337 26847 12371 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_85.VPB
flabel pwell 12337 26303 12371 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_85.VNB
rlabel comment 12400 26320 12400 26320 6 sr_0.FILLER_0_26_85.decap_12
flabel metal1 11233 26303 11267 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_97.VGND
flabel metal1 11233 26847 11267 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_97.VPWR
flabel nwell 11233 26847 11267 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_97.VPB
flabel pwell 11233 26303 11267 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_97.VNB
rlabel comment 11296 26320 11296 26320 6 sr_0.FILLER_0_26_97.decap_12
flabel metal1 12337 27391 12371 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_85.VGND
flabel metal1 12337 26847 12371 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_85.VPWR
flabel nwell 12337 26847 12371 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_85.VPB
flabel pwell 12337 27391 12371 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_85.VNB
rlabel comment 12400 27408 12400 27408 8 sr_0.FILLER_0_27_85.decap_12
flabel metal1 11233 26847 11267 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_97.VPWR
flabel metal1 11233 27391 11267 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_97.VGND
flabel nwell 11233 26847 11267 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_97.VPB
flabel pwell 11233 27391 11267 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_97.VNB
rlabel comment 11296 27408 11296 27408 8 sr_0.FILLER_0_27_97.decap_8
rlabel metal1 10560 27360 11296 27456 5 sr_0.FILLER_0_27_97.VGND
rlabel metal1 10560 26816 11296 26912 5 sr_0.FILLER_0_27_97.VPWR
flabel metal1 12417 26844 12470 26873 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_26_124.VPWR
flabel metal1 12420 26302 12471 26340 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_26_124.VGND
rlabel comment 12492 26320 12492 26320 6 sr_0.TAP_TAPCELL_ROW_26_124.tapvpwrvgnd_1
rlabel metal1 12400 26272 12492 26368 1 sr_0.TAP_TAPCELL_ROW_26_124.VGND
rlabel metal1 12400 26816 12492 26912 1 sr_0.TAP_TAPCELL_ROW_26_124.VPWR
flabel metal1 12417 26855 12470 26884 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_27_128.VPWR
flabel metal1 12420 27388 12471 27426 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_27_128.VGND
rlabel comment 12492 27408 12492 27408 8 sr_0.TAP_TAPCELL_ROW_27_128.tapvpwrvgnd_1
rlabel metal1 12400 27360 12492 27456 5 sr_0.TAP_TAPCELL_ROW_27_128.VGND
rlabel metal1 12400 26816 12492 26912 5 sr_0.TAP_TAPCELL_ROW_27_128.VPWR
flabel metal1 10129 26303 10163 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_109.VGND
flabel metal1 10129 26847 10163 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_109.VPWR
flabel nwell 10129 26847 10163 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_109.VPB
flabel pwell 10129 26303 10163 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_109.VNB
rlabel comment 10192 26320 10192 26320 6 sr_0.FILLER_0_26_109.decap_12
flabel metal1 9025 26303 9059 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_121.VGND
flabel metal1 9025 26847 9059 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_121.VPWR
flabel nwell 9025 26847 9059 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_121.VPB
flabel pwell 9025 26303 9059 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_121.VNB
rlabel comment 9088 26320 9088 26320 6 sr_0.FILLER_0_26_121.decap_12
flabel metal1 10487 27390 10540 27422 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_105.VGND
flabel metal1 10487 26847 10539 26878 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_105.VPWR
flabel nwell 10498 26855 10532 26873 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_105.VPB
flabel pwell 10497 27396 10529 27418 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_105.VNB
rlabel comment 10560 27408 10560 27408 8 sr_0.FILLER_0_27_105.fill_2
rlabel metal1 10376 27360 10560 27456 5 sr_0.FILLER_0_27_105.VGND
rlabel metal1 10376 26816 10560 26912 5 sr_0.FILLER_0_27_105.VPWR
flabel metal1 10027 27390 10080 27422 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_110.VGND
flabel metal1 10027 26847 10079 26878 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_110.VPWR
flabel nwell 10038 26855 10072 26873 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_110.VPB
flabel pwell 10037 27396 10069 27418 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_110.VNB
rlabel comment 10100 27408 10100 27408 8 sr_0.FILLER_0_27_110.fill_2
rlabel metal1 9916 27360 10100 27456 5 sr_0.FILLER_0_27_110.VGND
rlabel metal1 9916 26816 10100 26912 5 sr_0.FILLER_0_27_110.VPWR
flabel metal1 9761 27391 9795 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_113.VGND
flabel metal1 9761 26847 9795 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_113.VPWR
flabel nwell 9761 26847 9795 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_113.VPB
flabel pwell 9761 27391 9795 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_113.VNB
rlabel comment 9824 27408 9824 27408 8 sr_0.FILLER_0_27_113.decap_12
flabel metal1 8657 27391 8691 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_125.VGND
flabel metal1 8657 26847 8691 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_125.VPWR
flabel nwell 8657 26847 8691 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_125.VPB
flabel pwell 8657 27391 8691 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_125.VNB
rlabel comment 8720 27408 8720 27408 8 sr_0.FILLER_0_27_125.decap_12
flabel metal1 9841 26855 9894 26884 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_27_129.VPWR
flabel metal1 9844 27388 9895 27426 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_27_129.VGND
rlabel comment 9916 27408 9916 27408 8 sr_0.TAP_TAPCELL_ROW_27_129.tapvpwrvgnd_1
rlabel metal1 9824 27360 9916 27456 5 sr_0.TAP_TAPCELL_ROW_27_129.VGND
rlabel metal1 9824 26816 9916 26912 5 sr_0.TAP_TAPCELL_ROW_27_129.VPWR
flabel metal1 10131 27391 10165 27425 0 FreeSans 200 0 0 0 sr_0.input2.VGND
flabel metal1 10129 26847 10163 26881 0 FreeSans 200 0 0 0 sr_0.input2.VPWR
flabel locali 10129 26847 10163 26881 0 FreeSans 200 0 0 0 sr_0.input2.VPWR
flabel locali 10131 27391 10165 27425 0 FreeSans 200 0 0 0 sr_0.input2.VGND
flabel locali 10311 27289 10345 27323 0 FreeSans 200 0 0 0 sr_0.input2.X
flabel locali 10311 27017 10345 27051 0 FreeSans 200 0 0 0 sr_0.input2.X
flabel locali 10311 26949 10345 26983 0 FreeSans 200 0 0 0 sr_0.input2.X
flabel locali 10129 27153 10163 27187 0 FreeSans 200 0 0 0 sr_0.input2.A
flabel nwell 10129 26847 10163 26881 0 FreeSans 200 0 0 0 sr_0.input2.VPB
flabel pwell 10131 27391 10165 27425 0 FreeSans 200 0 0 0 sr_0.input2.VNB
rlabel comment 10100 27408 10100 27408 2 sr_0.input2.buf_1
rlabel metal1 10100 27360 10376 27456 5 sr_0.input2.VGND
rlabel metal1 10100 26816 10376 26912 5 sr_0.input2.VPWR
flabel metal1 7921 26847 7955 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_133.VPWR
flabel metal1 7921 26303 7955 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_133.VGND
flabel nwell 7921 26847 7955 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_133.VPB
flabel pwell 7921 26303 7955 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_133.VNB
rlabel comment 7984 26320 7984 26320 6 sr_0.FILLER_0_26_133.decap_6
rlabel metal1 7432 26272 7984 26368 1 sr_0.FILLER_0_26_133.VGND
rlabel metal1 7432 26816 7984 26912 1 sr_0.FILLER_0_26_133.VPWR
flabel metal1 7374 26847 7410 26877 0 FreeSans 250 0 0 0 sr_0.FILLER_0_26_139.VPWR
flabel metal1 7374 26307 7410 26336 0 FreeSans 250 0 0 0 sr_0.FILLER_0_26_139.VGND
flabel nwell 7381 26854 7401 26871 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_139.VPB
flabel pwell 7380 26309 7404 26331 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_139.VNB
rlabel comment 7432 26320 7432 26320 6 sr_0.FILLER_0_26_139.fill_1
rlabel metal1 7340 26272 7432 26368 1 sr_0.FILLER_0_26_139.VGND
rlabel metal1 7340 26816 7432 26912 1 sr_0.FILLER_0_26_139.VPWR
flabel metal1 7185 26303 7219 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_141.VGND
flabel metal1 7185 26847 7219 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_141.VPWR
flabel nwell 7185 26847 7219 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_141.VPB
flabel pwell 7185 26303 7219 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_141.VNB
rlabel comment 7248 26320 7248 26320 6 sr_0.FILLER_0_26_141.decap_12
flabel metal1 7553 26847 7587 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_137.VPWR
flabel metal1 7553 27391 7587 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_137.VGND
flabel nwell 7553 26847 7587 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_137.VPB
flabel pwell 7553 27391 7587 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_137.VNB
rlabel comment 7616 27408 7616 27408 8 sr_0.FILLER_0_27_137.decap_3
rlabel metal1 7340 27360 7616 27456 5 sr_0.FILLER_0_27_137.VGND
rlabel metal1 7340 26816 7616 26912 5 sr_0.FILLER_0_27_137.VPWR
flabel metal1 7185 27391 7219 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_141.VGND
flabel metal1 7185 26847 7219 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_141.VPWR
flabel nwell 7185 26847 7219 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_141.VPB
flabel pwell 7185 27391 7219 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_141.VNB
rlabel comment 7248 27408 7248 27408 8 sr_0.FILLER_0_27_141.decap_12
flabel metal1 7265 26844 7318 26873 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_26_125.VPWR
flabel metal1 7268 26302 7319 26340 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_26_125.VGND
rlabel comment 7340 26320 7340 26320 6 sr_0.TAP_TAPCELL_ROW_26_125.tapvpwrvgnd_1
rlabel metal1 7248 26272 7340 26368 1 sr_0.TAP_TAPCELL_ROW_26_125.VGND
rlabel metal1 7248 26816 7340 26912 1 sr_0.TAP_TAPCELL_ROW_26_125.VPWR
flabel metal1 7265 26855 7318 26884 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_27_130.VPWR
flabel metal1 7268 27388 7319 27426 0 FreeSans 200 0 0 0 sr_0.TAP_TAPCELL_ROW_27_130.VGND
rlabel comment 7340 27408 7340 27408 8 sr_0.TAP_TAPCELL_ROW_27_130.tapvpwrvgnd_1
rlabel metal1 7248 27360 7340 27456 5 sr_0.TAP_TAPCELL_ROW_27_130.VGND
rlabel metal1 7248 26816 7340 26912 5 sr_0.TAP_TAPCELL_ROW_27_130.VPWR
flabel metal1 6081 26847 6115 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_153.VPWR
flabel metal1 6081 26303 6115 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_153.VGND
flabel nwell 6081 26847 6115 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_153.VPB
flabel pwell 6081 26303 6115 26337 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_153.VNB
rlabel comment 6144 26320 6144 26320 6 sr_0.FILLER_0_26_153.decap_8
rlabel metal1 5408 26272 6144 26368 1 sr_0.FILLER_0_26_153.VGND
rlabel metal1 5408 26816 6144 26912 1 sr_0.FILLER_0_26_153.VPWR
flabel metal1 5335 26306 5388 26338 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_161.VGND
flabel metal1 5335 26850 5387 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_161.VPWR
flabel nwell 5346 26855 5380 26873 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_161.VPB
flabel pwell 5345 26310 5377 26332 0 FreeSans 200 0 0 0 sr_0.FILLER_0_26_161.VNB
rlabel comment 5408 26320 5408 26320 6 sr_0.FILLER_0_26_161.fill_2
rlabel metal1 5224 26272 5408 26368 1 sr_0.FILLER_0_26_161.VGND
rlabel metal1 5224 26816 5408 26912 1 sr_0.FILLER_0_26_161.VPWR
flabel metal1 6086 26851 6122 26881 0 FreeSans 250 0 0 0 sr_0.FILLER_0_27_153.VPWR
flabel metal1 6086 27392 6122 27421 0 FreeSans 250 0 0 0 sr_0.FILLER_0_27_153.VGND
flabel nwell 6093 26857 6113 26874 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_153.VPB
flabel pwell 6092 27397 6116 27419 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_153.VNB
rlabel comment 6144 27408 6144 27408 8 sr_0.FILLER_0_27_153.fill_1
rlabel metal1 6052 27360 6144 27456 5 sr_0.FILLER_0_27_153.VGND
rlabel metal1 6052 26816 6144 26912 5 sr_0.FILLER_0_27_153.VPWR
flabel metal1 5437 26847 5471 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_160.VPWR
flabel metal1 5437 27391 5471 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_160.VGND
flabel nwell 5437 26847 5471 26881 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_160.VPB
flabel pwell 5437 27391 5471 27425 0 FreeSans 200 0 0 0 sr_0.FILLER_0_27_160.VNB
rlabel comment 5500 27408 5500 27408 8 sr_0.FILLER_0_27_160.decap_3
rlabel metal1 5224 27360 5500 27456 5 sr_0.FILLER_0_27_160.VGND
rlabel metal1 5224 26816 5500 26912 5 sr_0.FILLER_0_27_160.VPWR
flabel metal1 4977 26847 5011 26881 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_26_Right_26.VPWR
flabel metal1 4977 26303 5011 26337 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_26_Right_26.VGND
flabel nwell 4977 26847 5011 26881 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_26_Right_26.VPB
flabel pwell 4977 26303 5011 26337 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_26_Right_26.VNB
rlabel comment 4948 26320 4948 26320 4 sr_0.PHY_EDGE_ROW_26_Right_26.decap_3
rlabel metal1 4948 26272 5224 26368 1 sr_0.PHY_EDGE_ROW_26_Right_26.VGND
rlabel metal1 4948 26816 5224 26912 1 sr_0.PHY_EDGE_ROW_26_Right_26.VPWR
flabel metal1 4977 26847 5011 26881 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_27_Right_27.VPWR
flabel metal1 4977 27391 5011 27425 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_27_Right_27.VGND
flabel nwell 4977 26847 5011 26881 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_27_Right_27.VPB
flabel pwell 4977 27391 5011 27425 0 FreeSans 200 0 0 0 sr_0.PHY_EDGE_ROW_27_Right_27.VNB
rlabel comment 4948 27408 4948 27408 2 sr_0.PHY_EDGE_ROW_27_Right_27.decap_3
rlabel metal1 4948 27360 5224 27456 5 sr_0.PHY_EDGE_ROW_27_Right_27.VGND
rlabel metal1 4948 26816 5224 26912 5 sr_0.PHY_EDGE_ROW_27_Right_27.VPWR
flabel locali 5621 27085 5655 27119 0 FreeSans 200 0 0 0 sr_0.input1.X
flabel locali 5897 27221 5931 27255 0 FreeSans 200 0 0 0 sr_0.input1.A
flabel locali 5529 27221 5563 27255 0 FreeSans 200 0 0 0 sr_0.input1.X
flabel locali 5897 27153 5931 27187 0 FreeSans 200 0 0 0 sr_0.input1.A
flabel locali 5529 27153 5563 27187 0 FreeSans 200 0 0 0 sr_0.input1.X
flabel metal1 5989 27391 6023 27425 0 FreeSans 200 0 0 0 sr_0.input1.VGND
flabel metal1 5989 26847 6023 26881 0 FreeSans 200 0 0 0 sr_0.input1.VPWR
flabel nwell 5989 26847 6023 26881 0 FreeSans 200 0 0 0 sr_0.input1.VPB
flabel pwell 5989 27391 6023 27425 0 FreeSans 200 0 0 0 sr_0.input1.VNB
rlabel comment 6052 27408 6052 27408 8 sr_0.input1.clkbuf_4
rlabel metal1 5500 27360 6052 27456 5 sr_0.input1.VGND
rlabel metal1 5500 26816 6052 26912 5 sr_0.input1.VPWR
flabel metal1 35230 5800 35430 5990 0 FreeSans 1600 0 0 0 ota_digpot_0.out
flabel metal1 0 2500 200 2690 0 FreeSans 1600 0 0 0 ota_digpot_0.gnd
flabel metal1 0 3440 200 3640 0 FreeSans 1600 0 0 0 ota_digpot_0.vd
flabel metal1 28700 0 28900 190 0 FreeSans 1600 0 0 0 ota_digpot_0.inp
flabel metal1 14050 40 14250 230 0 FreeSans 1600 0 0 0 ota_digpot_0.inn
flabel metal1 29200 9250 29400 9440 0 FreeSans 1600 0 0 0 ota_digpot_0.ib
flabel metal1 24710 9250 24910 9450 0 FreeSans 1600 0 0 0 ota_digpot_0.c0
flabel metal1 21180 9250 21380 9450 0 FreeSans 1600 0 0 0 ota_digpot_0.c1
flabel metal1 17550 9250 17750 9450 0 FreeSans 1600 0 0 0 ota_digpot_0.c2
flabel metal1 14010 9250 14210 9450 0 FreeSans 1600 0 0 0 ota_digpot_0.c3
flabel metal1 10500 9250 10700 9450 0 FreeSans 1600 0 0 0 ota_digpot_0.c4
flabel metal1 7260 9250 7460 9450 0 FreeSans 1600 0 0 0 ota_digpot_0.c5
flabel metal1 4030 9250 4230 9450 0 FreeSans 1600 0 0 0 ota_digpot_0.c6
flabel metal1 750 9250 950 9450 0 FreeSans 1600 0 0 0 ota_digpot_0.c7
flabel metal1 29200 3880 29400 4080 0 FreeSans 256 0 0 0 ota_digpot_0.ota_0.vs
flabel metal1 29210 5560 29410 5760 0 FreeSans 256 0 0 0 ota_digpot_0.ota_0.inn
flabel metal1 29210 4720 29410 4920 0 FreeSans 256 0 0 0 ota_digpot_0.ota_0.inp
flabel metal1 29200 5990 29400 6190 0 FreeSans 256 0 0 0 ota_digpot_0.ota_0.ib
flabel metal1 32050 7170 32250 7370 0 FreeSans 256 0 0 0 ota_digpot_0.ota_0.vd
flabel metal1 35030 5800 35230 6000 0 FreeSans 256 0 0 0 ota_digpot_0.ota_0.out
flabel metal1 30940 4690 30980 4710 0 FreeSans 1600 0 0 0 ota_digpot_0.ota_0.d
flabel metal1 30240 4690 30240 4710 0 FreeSans 1600 0 0 0 ota_digpot_0.ota_0.c
flabel metal2 30760 5910 30780 5930 0 FreeSans 1600 0 0 0 ota_digpot_0.ota_0.b
flabel metal1 24710 7340 24910 7540 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.c0
flabel metal1 21180 7340 21380 7540 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.c1
flabel metal1 17550 7340 17750 7540 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.c2
flabel metal1 14010 7340 14210 7540 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.c3
flabel metal1 10500 7340 10700 7540 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.c4
flabel metal1 7260 7340 7460 7540 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.c5
flabel metal1 4030 7340 4230 7540 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.c6
flabel metal1 750 7340 950 7540 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.c7
flabel metal1 14050 490 14250 690 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.n0
flabel metal1 28700 6550 28900 6750 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.n8
flabel metal1 200 2500 400 2700 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.gnd
flabel metal1 200 3440 400 3640 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.vd
flabel metal1 21750 3440 21950 3640 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_7.vd
flabel metal1 24150 3000 24350 3200 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_7.b
flabel metal1 21750 2500 21950 2700 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_7.vgnd
flabel metal1 21750 1860 21950 2060 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_7.ctrl
flabel metal1 24150 1720 24350 1920 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_7.a
flabel metal1 22470 4260 22490 4270 0 FreeSans 1600 0 0 0 ota_digpot_0.digpotp_0.tg_7.nctrl
flabel metal1 18050 3440 18250 3640 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_6.vd
flabel metal1 20450 3000 20650 3200 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_6.b
flabel metal1 18050 2500 18250 2700 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_6.vgnd
flabel metal1 18050 1860 18250 2060 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_6.ctrl
flabel metal1 20450 1720 20650 1920 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_6.a
flabel metal1 18770 4260 18790 4270 0 FreeSans 1600 0 0 0 ota_digpot_0.digpotp_0.tg_6.nctrl
flabel metal1 14550 3440 14750 3640 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_5.vd
flabel metal1 16950 3000 17150 3200 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_5.b
flabel metal1 14550 2500 14750 2700 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_5.vgnd
flabel metal1 14550 1860 14750 2060 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_5.ctrl
flabel metal1 16950 1720 17150 1920 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_5.a
flabel metal1 15270 4260 15290 4270 0 FreeSans 1600 0 0 0 ota_digpot_0.digpotp_0.tg_5.nctrl
flabel metal1 25550 3440 25750 3640 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_4.vd
flabel metal1 27950 3000 28150 3200 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_4.b
flabel metal1 25550 2500 25750 2700 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_4.vgnd
flabel metal1 25550 1860 25750 2060 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_4.ctrl
flabel metal1 27950 1720 28150 1920 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_4.a
flabel metal1 26270 4260 26290 4270 0 FreeSans 1600 0 0 0 ota_digpot_0.digpotp_0.tg_4.nctrl
flabel metal1 10950 3440 11150 3640 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_3.vd
flabel metal1 13350 3000 13550 3200 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_3.b
flabel metal1 10950 2500 11150 2700 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_3.vgnd
flabel metal1 10950 1860 11150 2060 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_3.ctrl
flabel metal1 13350 1720 13550 1920 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_3.a
flabel metal1 11670 4260 11690 4270 0 FreeSans 1600 0 0 0 ota_digpot_0.digpotp_0.tg_3.nctrl
flabel metal1 7650 3440 7850 3640 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_2.vd
flabel metal1 10050 3000 10250 3200 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_2.b
flabel metal1 7650 2500 7850 2700 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_2.vgnd
flabel metal1 7650 1860 7850 2060 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_2.ctrl
flabel metal1 10050 1720 10250 1920 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_2.a
flabel metal1 8370 4260 8390 4270 0 FreeSans 1600 0 0 0 ota_digpot_0.digpotp_0.tg_2.nctrl
flabel metal1 1050 3440 1250 3640 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_1.vd
flabel metal1 3450 3000 3650 3200 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_1.b
flabel metal1 1050 2500 1250 2700 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_1.vgnd
flabel metal1 1050 1860 1250 2060 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_1.ctrl
flabel metal1 3450 1720 3650 1920 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_1.a
flabel metal1 1770 4260 1790 4270 0 FreeSans 1600 0 0 0 ota_digpot_0.digpotp_0.tg_1.nctrl
flabel metal1 4350 3440 4550 3640 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_0.vd
flabel metal1 6750 3000 6950 3200 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_0.b
flabel metal1 4350 2500 4550 2700 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_0.vgnd
flabel metal1 4350 1860 4550 2060 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_0.ctrl
flabel metal1 6750 1720 6950 1920 0 FreeSans 256 0 0 0 ota_digpot_0.digpotp_0.tg_0.a
flabel metal1 5070 4260 5090 4270 0 FreeSans 1600 0 0 0 ota_digpot_0.digpotp_0.tg_0.nctrl
<< end >>
