magic
tech sky130A
magscale 1 2
timestamp 1698522569
<< psubdiff >>
rect 9590 3750 9770 3774
rect 9590 3546 9770 3570
<< psubdiffcont >>
rect 9590 3570 9770 3750
<< locali >>
rect 9590 3750 9770 3766
rect 9590 3554 9770 3570
<< viali >>
rect 9590 3570 9770 3750
<< metal1 >>
rect 9350 4690 9770 4700
rect 9350 4510 9580 4690
rect 9760 4510 9770 4690
rect 9350 4500 9770 4510
rect 9350 3750 9830 3760
rect 9350 3570 9590 3750
rect 9770 3570 9830 3750
rect 9350 3560 9830 3570
rect 9900 3120 10100 8600
rect 12550 7780 12850 7810
rect 12550 7540 12580 7780
rect 12800 7540 12850 7780
rect 12550 6710 12850 7540
rect 10190 4680 10410 4700
rect 10190 4500 10200 4680
rect 10380 4500 10410 4680
rect 10190 4490 10390 4500
rect 12600 4060 12800 6000
rect 10190 3750 10410 3760
rect 10190 3570 10210 3750
rect 10390 3570 10410 3750
rect 10190 3560 10410 3570
rect 13180 3120 13380 8600
rect 15850 7670 16150 7710
rect 15850 7550 15880 7670
rect 16090 7550 16150 7670
rect 15850 6610 16150 7550
rect 13490 4690 13710 4700
rect 13490 4510 13510 4690
rect 13690 4510 13710 4690
rect 13490 4500 13710 4510
rect 15900 4060 16100 6000
rect 13490 3750 13710 3760
rect 13490 3570 13500 3750
rect 13680 3570 13710 3750
rect 13490 3560 13710 3570
rect 16410 3120 16610 8600
rect 19150 7790 19450 7830
rect 19150 7530 19190 7790
rect 19390 7530 19450 7790
rect 19150 6730 19450 7530
rect 16790 4690 17010 4700
rect 16790 4510 16810 4690
rect 16990 4510 17010 4690
rect 16790 4500 17010 4510
rect 19200 4060 19400 6000
rect 16790 3750 17010 3760
rect 16790 3570 16810 3750
rect 16990 3570 17010 3750
rect 16790 3560 17010 3570
rect 19650 3120 19850 8600
rect 22460 7850 22760 7950
rect 22460 7540 22510 7850
rect 22710 7540 22760 7850
rect 22460 6850 22760 7540
rect 20090 4690 20310 4700
rect 20090 4510 20110 4690
rect 20290 4510 20310 4690
rect 20090 4500 20310 4510
rect 22500 4060 22700 6000
rect 20090 3750 20310 3760
rect 20090 3570 20110 3750
rect 20290 3570 20310 3750
rect 20090 3560 20310 3570
rect 23160 3120 23360 8600
rect 26000 7870 26350 7920
rect 26000 7560 26080 7870
rect 26300 7560 26350 7870
rect 26000 7520 26350 7560
rect 23690 4690 23910 4700
rect 23690 4510 23710 4690
rect 23890 4510 23910 4690
rect 23690 4500 23910 4510
rect 26100 4060 26300 6000
rect 23690 3750 23910 3760
rect 23690 3570 23700 3750
rect 23880 3570 23910 3750
rect 23690 3560 23910 3570
rect 26700 3120 26900 8600
rect 28600 7840 29020 7900
rect 28600 7550 28640 7840
rect 28970 7550 29020 7840
rect 28600 6300 29020 7550
rect 29400 7410 29730 7770
rect 28600 5880 29410 6300
rect 27190 4690 27410 4700
rect 27190 4510 27210 4690
rect 27390 4510 27410 4690
rect 27190 4500 27410 4510
rect 29600 4060 29800 6000
rect 27190 3740 27410 3760
rect 27190 3560 27210 3740
rect 27390 3560 27410 3740
rect 27200 3550 27400 3560
rect 30330 3120 30530 8600
rect 31665 7840 32075 7905
rect 31665 7560 31710 7840
rect 32010 7560 32075 7840
rect 31665 6280 32075 7560
rect 32500 7390 32830 7750
rect 33140 7410 33470 7770
rect 31665 5870 32510 6280
rect 32810 5870 33140 6230
rect 30890 4690 31110 4700
rect 30890 4510 30910 4690
rect 31090 4510 31110 4690
rect 30890 4500 31110 4510
rect 33300 4060 33500 6000
rect 30890 3750 31110 3760
rect 30890 3570 30910 3750
rect 31090 3570 31110 3750
rect 30890 3560 31110 3570
rect 33860 3120 34060 8600
rect 37480 7910 37850 7930
rect 34275 7770 34705 7835
rect 34275 7550 34320 7770
rect 34650 7550 34705 7770
rect 34275 6300 34705 7550
rect 35000 7420 35330 7780
rect 35630 7400 35960 7760
rect 36280 7400 36580 7800
rect 36900 7400 37230 7800
rect 37480 7580 37530 7910
rect 37740 7810 37850 7910
rect 37740 7610 38050 7810
rect 37740 7580 37850 7610
rect 37480 7540 37850 7580
rect 34275 5870 35020 6300
rect 35320 5890 35650 6250
rect 35950 5890 36280 6250
rect 36600 5880 36900 6280
rect 34690 4690 34910 4700
rect 34690 4510 34710 4690
rect 34890 4510 34910 4690
rect 34690 4500 34910 4510
rect 37100 4060 37300 6000
rect 34690 3750 34910 3760
rect 34690 3570 34710 3750
rect 34890 3570 34910 3750
rect 34690 3560 34910 3570
rect 9900 2920 10400 3120
rect 12600 2310 12800 2980
rect 13180 2920 13700 3120
rect 15900 2310 16100 2980
rect 16410 2920 17000 3120
rect 19200 2310 19400 2980
rect 19650 2920 20300 3120
rect 22500 2310 22700 2980
rect 23160 2920 23900 3120
rect 26100 2310 26300 2980
rect 26700 2920 27400 3120
rect 29600 2310 29800 2980
rect 30330 2920 31100 3120
rect 33300 2310 33500 2980
rect 33860 2920 34900 3120
rect 37100 2310 37300 2980
rect 12600 2110 37300 2310
rect 23200 1550 23400 2110
<< via1 >>
rect 9580 4510 9760 4690
rect 9590 3570 9770 3750
rect 12580 7540 12800 7780
rect 10200 4500 10380 4680
rect 10210 3570 10390 3750
rect 15880 7550 16090 7670
rect 13510 4510 13690 4690
rect 13500 3570 13680 3750
rect 19190 7530 19390 7790
rect 16810 4510 16990 4690
rect 16810 3570 16990 3750
rect 22510 7540 22710 7850
rect 20110 4510 20290 4690
rect 20110 3570 20290 3750
rect 26080 7560 26300 7870
rect 23710 4510 23890 4690
rect 23700 3570 23880 3750
rect 28640 7550 28970 7840
rect 27210 4510 27390 4690
rect 27210 3560 27390 3740
rect 31710 7560 32010 7840
rect 30910 4510 31090 4690
rect 30910 3570 31090 3750
rect 34320 7550 34650 7770
rect 37530 7580 37740 7910
rect 34710 4510 34890 4690
rect 34710 3570 34890 3750
<< metal2 >>
rect 12550 7910 37760 7940
rect 12550 7870 37530 7910
rect 12550 7850 26080 7870
rect 12550 7790 22510 7850
rect 12550 7780 19190 7790
rect 12550 7540 12580 7780
rect 12800 7670 19190 7780
rect 12800 7550 15880 7670
rect 16090 7550 19190 7670
rect 12800 7540 19190 7550
rect 12550 7530 19190 7540
rect 19390 7540 22510 7790
rect 22710 7560 26080 7850
rect 26300 7840 37530 7870
rect 26300 7560 28640 7840
rect 22710 7550 28640 7560
rect 28970 7560 31710 7840
rect 32010 7770 37530 7840
rect 32010 7560 34320 7770
rect 28970 7550 34320 7560
rect 34650 7580 37530 7770
rect 37740 7580 37760 7910
rect 34650 7550 37760 7580
rect 22710 7540 37760 7550
rect 19390 7530 37760 7540
rect 12550 7520 37760 7530
rect 9570 4690 9770 4700
rect 13500 4690 13700 4700
rect 9570 4510 9580 4690
rect 9760 4510 9770 4690
rect 9570 4500 9770 4510
rect 10190 4680 10390 4690
rect 10190 4500 10200 4680
rect 10380 4500 10390 4680
rect 13500 4510 13510 4690
rect 13690 4510 13700 4690
rect 13500 4500 13700 4510
rect 16800 4690 17000 4700
rect 16800 4510 16810 4690
rect 16990 4510 17000 4690
rect 16800 4500 17000 4510
rect 20100 4690 20300 4700
rect 20100 4510 20110 4690
rect 20290 4510 20300 4690
rect 20100 4500 20300 4510
rect 23700 4690 23900 4700
rect 23700 4510 23710 4690
rect 23890 4510 23900 4690
rect 23700 4500 23900 4510
rect 27200 4690 27400 4700
rect 27200 4510 27210 4690
rect 27390 4510 27400 4690
rect 27200 4500 27400 4510
rect 30900 4690 31100 4700
rect 30900 4510 30910 4690
rect 31090 4510 31100 4690
rect 30900 4500 31100 4510
rect 34700 4690 34900 4700
rect 34700 4510 34710 4690
rect 34890 4510 34900 4690
rect 34700 4500 34900 4510
rect 10190 4490 10390 4500
rect 9580 3750 9800 3760
rect 9580 3570 9590 3750
rect 9770 3570 9800 3750
rect 9580 3560 9800 3570
rect 10200 3750 10400 3760
rect 10200 3570 10210 3750
rect 10390 3570 10400 3750
rect 10200 3560 10400 3570
rect 13490 3750 13690 3760
rect 13490 3570 13500 3750
rect 13680 3570 13690 3750
rect 13490 3560 13690 3570
rect 16800 3750 17000 3760
rect 16800 3570 16810 3750
rect 16990 3570 17000 3750
rect 16800 3560 17000 3570
rect 20100 3750 20300 3760
rect 20100 3570 20110 3750
rect 20290 3570 20300 3750
rect 20100 3560 20300 3570
rect 23690 3750 23890 3760
rect 30900 3750 31100 3760
rect 23690 3570 23700 3750
rect 23880 3570 23890 3750
rect 23690 3560 23890 3570
rect 27200 3740 27400 3750
rect 27200 3560 27210 3740
rect 27390 3560 27400 3740
rect 30900 3570 30910 3750
rect 31090 3570 31100 3750
rect 30900 3560 31100 3570
rect 34700 3750 34900 3760
rect 34700 3570 34710 3750
rect 34890 3570 34900 3750
rect 34700 3560 34900 3570
rect 27200 3550 27400 3560
<< via2 >>
rect 9580 4510 9760 4690
rect 10200 4500 10380 4680
rect 13510 4510 13690 4690
rect 16810 4510 16990 4690
rect 20110 4510 20290 4690
rect 23710 4510 23890 4690
rect 27210 4510 27390 4690
rect 30910 4510 31090 4690
rect 34710 4510 34890 4690
rect 9590 3570 9770 3750
rect 10210 3570 10390 3750
rect 13500 3570 13680 3750
rect 16810 3570 16990 3750
rect 20110 3570 20290 3750
rect 23700 3570 23880 3750
rect 27210 3560 27390 3740
rect 30910 3570 31090 3750
rect 34710 3570 34890 3750
<< metal3 >>
rect 9570 4690 34900 4710
rect 9570 4510 9580 4690
rect 9760 4680 13510 4690
rect 9760 4510 10200 4680
rect 9570 4500 10200 4510
rect 10380 4510 13510 4680
rect 13690 4510 16810 4690
rect 16990 4510 20110 4690
rect 20290 4510 23710 4690
rect 23890 4510 27210 4690
rect 27390 4510 30910 4690
rect 31090 4510 34710 4690
rect 34890 4510 34900 4690
rect 10380 4500 34900 4510
rect 9570 4490 34900 4500
rect 9580 3750 34900 3770
rect 9580 3570 9590 3750
rect 9770 3570 10210 3750
rect 10390 3570 13500 3750
rect 13680 3570 16810 3750
rect 16990 3570 20110 3750
rect 20290 3570 23700 3750
rect 23880 3740 30910 3750
rect 23880 3570 27210 3740
rect 9580 3560 27210 3570
rect 27390 3570 30910 3740
rect 31090 3570 34710 3750
rect 34890 3570 34900 3750
rect 27390 3560 34900 3570
rect 9580 3550 34900 3560
use sky130_fd_pr__res_high_po_0p35_52KWSA  XR1
timestamp 1698520721
transform 1 0 12701 0 1 6398
box -201 -698 201 698
use sky130_fd_pr__res_xhigh_po_0p35_9P2C6Q  XR2
timestamp 1698520721
transform 1 0 16001 0 1 6350
box -201 -650 201 650
use sky130_fd_pr__res_xhigh_po_0p35_URGAGF  XR3
timestamp 1698520721
transform 1 0 19301 0 1 6420
box -201 -720 201 720
use sky130_fd_pr__res_xhigh_po_0p35_U5HPMT  XR4
timestamp 1698520721
transform 1 0 22601 0 1 6560
box -201 -860 201 860
use sky130_fd_pr__res_xhigh_po_0p35_WZM67X  XR5
timestamp 1698520721
transform 1 0 26201 0 1 6840
box -201 -1140 201 1140
use sky130_fd_pr__res_xhigh_po_0p35_WR52AX  XR6
timestamp 1698522189
transform 1 0 29560 0 1 6840
box -360 -1140 360 1140
use sky130_fd_pr__res_xhigh_po_0p35_QD939Z  XR7
timestamp 1698522189
transform 1 0 32978 0 1 6840
box -678 -1140 678 1140
use sky130_fd_pr__res_xhigh_po_0p35_2TH3B8  XR8
timestamp 1698522189
transform 1 0 36114 0 1 6840
box -1314 -1140 1314 1140
use tg  tg_0 /foss/designs/projects/dpga2/magic/ota_digpot/digpot/tg
timestamp 1698520465
transform 1 0 14200 0 1 1920
box -700 580 1900 3660
use tg  tg_1
timestamp 1698520465
transform 1 0 10900 0 1 1920
box -700 580 1900 3660
use tg  tg_2
timestamp 1698520465
transform 1 0 17500 0 1 1920
box -700 580 1900 3660
use tg  tg_3
timestamp 1698520465
transform 1 0 20800 0 1 1920
box -700 580 1900 3660
use tg  tg_4
timestamp 1698520465
transform 1 0 35400 0 1 1920
box -700 580 1900 3660
use tg  tg_5
timestamp 1698520465
transform 1 0 24400 0 1 1920
box -700 580 1900 3660
use tg  tg_6
timestamp 1698520465
transform 1 0 27900 0 1 1920
box -700 580 1900 3660
use tg  tg_7
timestamp 1698520465
transform 1 0 31600 0 1 1920
box -700 580 1900 3660
<< labels >>
flabel metal1 33860 8400 34060 8600 0 FreeSans 256 0 0 0 c0
port 2 nsew
flabel metal1 30330 8400 30530 8600 0 FreeSans 256 0 0 0 c1
port 3 nsew
flabel metal1 26700 8400 26900 8600 0 FreeSans 256 0 0 0 c2
port 6 nsew
flabel metal1 23160 8400 23360 8600 0 FreeSans 256 0 0 0 c3
port 7 nsew
flabel metal1 19650 8400 19850 8600 0 FreeSans 256 0 0 0 c4
port 8 nsew
flabel metal1 16410 8400 16610 8600 0 FreeSans 256 0 0 0 c5
port 9 nsew
flabel metal1 13180 8400 13380 8600 0 FreeSans 256 0 0 0 c6
port 10 nsew
flabel metal1 9900 8400 10100 8600 0 FreeSans 256 0 0 0 c7
port 11 nsew
flabel metal1 23200 1550 23400 1750 0 FreeSans 256 0 0 0 n0
port 4 nsew
flabel metal1 37850 7610 38050 7810 0 FreeSans 256 0 0 0 n8
port 5 nsew
flabel metal1 9350 3560 9550 3760 0 FreeSans 256 0 0 0 gnd
port 0 nsew
flabel metal1 9350 4500 9550 4700 0 FreeSans 256 0 0 0 vd
port 1 nsew
<< end >>
