* NGSPICE file created from digpotp.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_ECDJHW a_n129_n500# a_n513_n500# a_399_n588# a_63_n500#
+ a_n225_n500# a_495_522# a_n321_n500# a_111_522# a_207_n588# a_n33_n500# a_n369_n588#
+ a_303_522# a_447_n500# a_n605_n500# a_15_n588# a_n81_522# a_n561_n588# a_543_n500#
+ a_159_n500# a_n177_n588# a_n273_522# a_255_n500# a_351_n500# a_n417_n500# a_n465_522#
+ VSUBS
X0 a_n417_n500# a_n465_522# a_n513_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X1 a_n33_n500# a_n81_522# a_n129_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X2 a_351_n500# a_303_522# a_255_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X3 a_255_n500# a_207_n588# a_159_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X4 a_n321_n500# a_n369_n588# a_n417_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.65e+12p pd=1.066e+07u as=0p ps=0u w=5e+06u l=150000u
X5 a_543_n500# a_495_522# a_447_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.55e+12p pd=1.062e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X6 a_159_n500# a_111_522# a_63_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X7 a_n225_n500# a_n273_522# a_n321_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.65e+12p pd=1.066e+07u as=0p ps=0u w=5e+06u l=150000u
X8 a_447_n500# a_399_n588# a_351_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9 a_n513_n500# a_n561_n588# a_n605_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.55e+12p ps=1.062e+07u w=5e+06u l=150000u
X10 a_63_n500# a_15_n588# a_n33_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X11 a_n129_n500# a_n177_n588# a_n225_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_8QR85J a_15_n500# w_n109_n600# a_n33_n597# a_n73_n500#
X0 a_15_n500# a_n33_n597# a_n73_n500# w_n109_n600# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_VU5CXM a_15_n500# a_n73_n500# a_n33_n588# VSUBS
X0 a_15_n500# a_n33_n588# a_n73_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_4W7PEP a_n73_n100# a_n33_n188# a_15_n100# VSUBS
X0 a_15_n100# a_n33_n188# a_n73_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_XGAKDL a_n33_n397# a_n73_n300# a_15_n300# w_n109_n400#
X0 a_15_n300# a_n33_n397# a_n73_n300# w_n109_n400# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_VQ5UWM a_15_n500# a_n73_n500# a_n33_n588# VSUBS
X0 a_15_n500# a_n33_n588# a_n73_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_UGA66J a_15_n500# w_n109_n600# a_n33_n597# a_n73_n500#
X0 a_15_n500# a_n33_n597# a_n73_n500# w_n109_n600# sky130_fd_pr__pfet_01v8 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_PM4G2P a_n129_n500# a_n513_n500# a_63_n500# a_15_n597#
+ a_n81_531# a_n225_n500# a_n177_n597# a_n561_n597# a_n273_531# a_n321_n500# w_n641_n600#
+ a_n33_n500# a_n465_531# a_447_n500# a_n605_n500# a_399_n597# a_543_n500# a_159_n500#
+ a_495_531# a_111_531# a_255_n500# a_207_n597# a_351_n500# a_n417_n500# a_n369_n597#
+ a_303_531#
X0 a_n33_n500# a_n81_531# a_n129_n500# w_n641_n600# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X1 a_351_n500# a_303_531# a_255_n500# w_n641_n600# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X2 a_255_n500# a_207_n597# a_159_n500# w_n641_n600# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X3 a_n321_n500# a_n369_n597# a_n417_n500# w_n641_n600# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X4 a_543_n500# a_495_531# a_447_n500# w_n641_n600# sky130_fd_pr__pfet_01v8 ad=1.55e+12p pd=1.062e+07u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X5 a_159_n500# a_111_531# a_63_n500# w_n641_n600# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.65e+12p ps=1.066e+07u w=5e+06u l=150000u
X6 a_n225_n500# a_n273_531# a_n321_n500# w_n641_n600# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=0p ps=0u w=5e+06u l=150000u
X7 a_447_n500# a_399_n597# a_351_n500# w_n641_n600# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8 a_n513_n500# a_n561_n597# a_n605_n500# w_n641_n600# sky130_fd_pr__pfet_01v8 ad=1.65e+12p pd=1.066e+07u as=1.55e+12p ps=1.062e+07u w=5e+06u l=150000u
X9 a_63_n500# a_15_n597# a_n33_n500# w_n641_n600# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X10 a_n129_n500# a_n177_n597# a_n225_n500# w_n641_n600# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X11 a_n417_n500# a_n465_531# a_n513_n500# w_n641_n600# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
.ends

.subckt tg vd vgnd b a ctrl
Xsky130_fd_pr__nfet_01v8_ECDJHW_0 a a ctrl a b ctrl a ctrl ctrl b ctrl ctrl a b ctrl
+ ctrl ctrl b b ctrl ctrl a b b ctrl vgnd sky130_fd_pr__nfet_01v8_ECDJHW
XXM2 vd vd vd vd sky130_fd_pr__pfet_01v8_8QR85J
Xsky130_fd_pr__nfet_01v8_VU5CXM_0 a a a vgnd sky130_fd_pr__nfet_01v8_VU5CXM
XXM3 vgnd ctrl nctrl vgnd sky130_fd_pr__nfet_01v8_4W7PEP
XXM4 ctrl vd nctrl vd sky130_fd_pr__pfet_01v8_XGAKDL
Xsky130_fd_pr__nfet_01v8_VQ5UWM_1 vgnd vgnd vgnd vgnd sky130_fd_pr__nfet_01v8_VQ5UWM
Xsky130_fd_pr__pfet_01v8_UGA66J_0 b vd b b sky130_fd_pr__pfet_01v8_UGA66J
Xsky130_fd_pr__pfet_01v8_PM4G2P_0 b b b nctrl nctrl a nctrl nctrl nctrl b vd a nctrl
+ b a nctrl a a nctrl nctrl b nctrl a a nctrl nctrl sky130_fd_pr__pfet_01v8_PM4G2P
.ends

.subckt sky130_fd_pr__res_high_po_0p35_52KWSA a_n165_n662# a_n35_n532# a_n35_100#
X0 a_n35_n532# a_n35_100# a_n165_n662# sky130_fd_pr__res_high_po_0p35 l=1e+06u
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_9P2C6Q a_n35_n484# a_n165_n614# a_n35_52#
X0 a_n35_n484# a_n35_52# a_n165_n614# sky130_fd_pr__res_xhigh_po_0p35 l=520000u
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_URGAGF a_n35_122# a_n35_n554# a_n165_n684#
X0 a_n35_n554# a_n35_122# a_n165_n684# sky130_fd_pr__res_xhigh_po_0p35 l=1.22e+06u
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_WZM67X a_n35_n974# a_n35_542# a_n165_n1104#
X0 a_n35_n974# a_n35_542# a_n165_n1104# sky130_fd_pr__res_xhigh_po_0p35 l=5.42e+06u
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_U5HPMT a_n35_n694# a_n165_n824# a_n35_262#
X0 a_n35_n694# a_n35_262# a_n165_n824# sky130_fd_pr__res_xhigh_po_0p35 l=2.62e+06u
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_WR52AX a_n194_n974# a_124_542# a_n194_542#
+ a_124_n974# a_n324_n1104#
X0 a_124_n974# a_124_542# a_n324_n1104# sky130_fd_pr__res_xhigh_po_0p35 l=5.42e+06u
X1 a_n194_n974# a_n194_542# a_n324_n1104# sky130_fd_pr__res_xhigh_po_0p35 l=5.42e+06u
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_QD939Z a_n194_n974# a_442_542# a_124_542#
+ a_n194_542# a_n642_n1104# a_n512_n974# a_124_n974# a_n512_542# a_442_n974#
X0 a_n512_n974# a_n512_542# a_n642_n1104# sky130_fd_pr__res_xhigh_po_0p35 l=5.42e+06u
X1 a_124_n974# a_124_542# a_n642_n1104# sky130_fd_pr__res_xhigh_po_0p35 l=5.42e+06u
X2 a_n194_n974# a_n194_542# a_n642_n1104# sky130_fd_pr__res_xhigh_po_0p35 l=5.42e+06u
X3 a_442_n974# a_442_542# a_n642_n1104# sky130_fd_pr__res_xhigh_po_0p35 l=5.42e+06u
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_2TH3B8 a_1078_542# a_760_542# a_1078_n974#
+ a_n194_n974# a_442_542# a_760_n974# a_124_542# a_n194_542# a_n512_n974# a_124_n974#
+ a_n1148_n974# a_n1148_542# a_n830_542# a_n1278_n1104# a_n512_542# a_n830_n974# a_442_n974#
X0 a_n830_n974# a_n830_542# a_n1278_n1104# sky130_fd_pr__res_xhigh_po_0p35 l=5.42e+06u
X1 a_n512_n974# a_n512_542# a_n1278_n1104# sky130_fd_pr__res_xhigh_po_0p35 l=5.42e+06u
X2 a_124_n974# a_124_542# a_n1278_n1104# sky130_fd_pr__res_xhigh_po_0p35 l=5.42e+06u
X3 a_n194_n974# a_n194_542# a_n1278_n1104# sky130_fd_pr__res_xhigh_po_0p35 l=5.42e+06u
X4 a_n1148_n974# a_n1148_542# a_n1278_n1104# sky130_fd_pr__res_xhigh_po_0p35 l=5.42e+06u
X5 a_442_n974# a_442_542# a_n1278_n1104# sky130_fd_pr__res_xhigh_po_0p35 l=5.42e+06u
X6 a_1078_n974# a_1078_542# a_n1278_n1104# sky130_fd_pr__res_xhigh_po_0p35 l=5.42e+06u
X7 a_760_n974# a_760_542# a_n1278_n1104# sky130_fd_pr__res_xhigh_po_0p35 l=5.42e+06u
.ends

.subckt digpotp gnd vd c0 c1 n0 n8 c2 c3 c4 c5 c6 c7
Xtg_0 vd gnd tg_0/b n0 c6 tg
Xtg_2 vd gnd tg_2/b n0 c5 tg
Xtg_1 vd gnd tg_1/b n0 c7 tg
Xtg_3 vd gnd tg_3/b n0 c4 tg
Xtg_4 vd gnd tg_4/b n0 c0 tg
Xtg_5 vd gnd tg_5/b n0 c3 tg
Xtg_6 vd gnd tg_6/b n0 c2 tg
XXR1 gnd tg_1/b n8 sky130_fd_pr__res_high_po_0p35_52KWSA
Xtg_7 vd gnd tg_7/b n0 c1 tg
XXR2 tg_0/b gnd n8 sky130_fd_pr__res_xhigh_po_0p35_9P2C6Q
XXR3 n8 tg_2/b gnd sky130_fd_pr__res_xhigh_po_0p35_URGAGF
XXR5 tg_5/b n8 gnd sky130_fd_pr__res_xhigh_po_0p35_WZM67X
XXR4 tg_3/b gnd n8 sky130_fd_pr__res_xhigh_po_0p35_U5HPMT
XXR6 n8 m1_29400_7410# m1_29400_7410# tg_6/b gnd sky130_fd_pr__res_xhigh_po_0p35_WR52AX
XXR7 m1_32810_5870# m1_33140_7410# m1_33140_7410# m1_32500_7390# gnd n8 m1_32810_5870#
+ m1_32500_7390# tg_7/b sky130_fd_pr__res_xhigh_po_0p35_QD939Z
XXR8 m1_36900_7400# m1_36900_7400# tg_4/b m1_35950_5890# m1_36280_7400# m1_36600_5880#
+ m1_36280_7400# m1_35630_7400# m1_35320_5890# m1_35950_5890# n8 m1_35000_7420# m1_35000_7420#
+ gnd m1_35630_7400# m1_35320_5890# m1_36600_5880# sky130_fd_pr__res_xhigh_po_0p35_2TH3B8
.ends

