magic
tech sky130A
magscale 1 2
timestamp 1698520721
<< pwell >>
rect -201 -5060 201 5060
<< psubdiff >>
rect -165 4990 -69 5024
rect 69 4990 165 5024
rect -165 4928 -131 4990
rect 131 4928 165 4990
rect -165 -4990 -131 -4928
rect 131 -4990 165 -4928
rect -165 -5024 -69 -4990
rect 69 -5024 165 -4990
<< psubdiffcont >>
rect -69 4990 69 5024
rect -165 -4928 -131 4928
rect 131 -4928 165 4928
rect -69 -5024 69 -4990
<< xpolycontact >>
rect -35 4462 35 4894
rect -35 -4894 35 -4462
<< xpolyres >>
rect -35 -4462 35 4462
<< locali >>
rect -165 4990 -69 5024
rect 69 4990 165 5024
rect -165 4928 -131 4990
rect 131 4928 165 4990
rect -165 -4990 -131 -4928
rect 131 -4990 165 -4928
rect -165 -5024 -69 -4990
rect 69 -5024 165 -4990
<< viali >>
rect -19 4479 19 4876
rect -19 -4876 19 -4479
<< metal1 >>
rect -25 4876 25 4888
rect -25 4479 -19 4876
rect 19 4479 25 4876
rect -25 4467 25 4479
rect -25 -4479 25 -4467
rect -25 -4876 -19 -4479
rect 19 -4876 25 -4479
rect -25 -4888 25 -4876
<< res0p35 >>
rect -37 -4464 37 4464
<< properties >>
string FIXED_BBOX -148 -5007 148 5007
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 44.62 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 256.046k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
