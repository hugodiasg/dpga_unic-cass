** sch_path: /foss/designs/projects/dpga2/xschem/digpotp.sch
.subckt digpotp gnd vd c0 c1 n0 n8 c2 c3 c4 c5 c6 c7
*.PININFO gnd:B vd:B c0:I c1:I n0:I n8:O c2:I c3:I c4:I c5:I c6:I c7:I
x9 c0 vd net2 gnd n0 tg
x10 c1 vd net1 gnd n0 tg
x7 c2 vd net3 gnd n0 tg
x8 c3 vd net4 gnd n0 tg
x11 c4 vd net5 gnd n0 tg
x12 c5 vd net6 gnd n0 tg
x1 c6 vd net7 gnd n0 tg
x2 c7 vd net8 gnd n0 tg
XR2 n8 net7 gnd sky130_fd_pr__res_xhigh_po_0p35 L=0.52 mult=1 m=1
XR3 n8 net6 gnd sky130_fd_pr__res_xhigh_po_0p35 L=1.22 mult=1 m=1
XR4 n8 net5 gnd sky130_fd_pr__res_xhigh_po_0p35 L=2.62 mult=1 m=1
XR5 n8 net4 gnd sky130_fd_pr__res_xhigh_po_0p35 L=5.42 mult=1 m=1
XR6 n8 net3 gnd sky130_fd_pr__res_xhigh_po_0p35 L=11.02 mult=1 m=1
XR7 n8 net1 gnd sky130_fd_pr__res_xhigh_po_0p35 L=22.22 mult=1 m=1
XR8 n8 net2 gnd sky130_fd_pr__res_xhigh_po_0p35 L=44.62 mult=1 m=1
XR1 n8 net8 gnd sky130_fd_pr__res_high_po_0p35 L=1 mult=1 m=1
.ends

* expanding   symbol:  projects/dpga-ieee-sscs-contest/xschem/tg.sym # of pins=5
** sym_path: /foss/designs/projects/dpga-ieee-sscs-contest/xschem/tg.sym
** sch_path: /foss/designs/projects/dpga-ieee-sscs-contest/xschem/tg.sch
.subckt tg ctrl vd b vgnd a
*.PININFO vd:B vgnd:B b:B a:B ctrl:I
XM2 b nctrl a vd sky130_fd_pr__pfet_01v8 L=0.15 W=60 nf=12 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 a ctrl b vgnd sky130_fd_pr__nfet_01v8 L=0.15 W=60 nf=12 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 nctrl ctrl vgnd vgnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 nctrl ctrl vd vd sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 vd vd vd vd sky130_fd_pr__pfet_01v8 L=0.15 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 b b b vd sky130_fd_pr__pfet_01v8 L=0.15 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 vgnd vgnd vgnd vgnd sky130_fd_pr__nfet_01v8 L=0.15 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 a a a vgnd sky130_fd_pr__nfet_01v8 L=0.15 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
