magic
tech sky130A
magscale 1 2
timestamp 1698511094
<< metal3 >>
rect -2550 1572 2549 1600
rect -2550 -1572 2465 1572
rect 2529 -1572 2549 1572
rect -2550 -1600 2549 -1572
<< via3 >>
rect 2465 -1572 2529 1572
<< mimcap >>
rect -2450 1460 2350 1500
rect -2450 -1460 -2410 1460
rect 2310 -1460 2350 1460
rect -2450 -1500 2350 -1460
<< mimcapcontact >>
rect -2410 -1460 2310 1460
<< metal4 >>
rect 2449 1572 2545 1588
rect -2411 1460 2311 1461
rect -2411 -1460 -2410 1460
rect 2310 -1460 2311 1460
rect -2411 -1461 2311 -1460
rect 2449 -1572 2465 1572
rect 2529 -1572 2545 1572
rect 2449 -1588 2545 -1572
<< properties >>
string FIXED_BBOX -2550 -1600 2450 1600
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 24 l 15 val 734.82 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
