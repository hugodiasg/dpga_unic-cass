magic
tech sky130A
magscale 1 2
timestamp 1698522189
<< pwell >>
rect -1314 -1140 1314 1140
<< psubdiff >>
rect -1278 1070 -1182 1104
rect 1182 1070 1278 1104
rect -1278 1008 -1244 1070
rect 1244 1008 1278 1070
rect -1278 -1070 -1244 -1008
rect 1244 -1070 1278 -1008
rect -1278 -1104 -1182 -1070
rect 1182 -1104 1278 -1070
<< psubdiffcont >>
rect -1182 1070 1182 1104
rect -1278 -1008 -1244 1008
rect 1244 -1008 1278 1008
rect -1182 -1104 1182 -1070
<< xpolycontact >>
rect -1148 542 -1078 974
rect -1148 -974 -1078 -542
rect -830 542 -760 974
rect -830 -974 -760 -542
rect -512 542 -442 974
rect -512 -974 -442 -542
rect -194 542 -124 974
rect -194 -974 -124 -542
rect 124 542 194 974
rect 124 -974 194 -542
rect 442 542 512 974
rect 442 -974 512 -542
rect 760 542 830 974
rect 760 -974 830 -542
rect 1078 542 1148 974
rect 1078 -974 1148 -542
<< xpolyres >>
rect -1148 -542 -1078 542
rect -830 -542 -760 542
rect -512 -542 -442 542
rect -194 -542 -124 542
rect 124 -542 194 542
rect 442 -542 512 542
rect 760 -542 830 542
rect 1078 -542 1148 542
<< locali >>
rect -1278 1070 -1182 1104
rect 1182 1070 1278 1104
rect -1278 1008 -1244 1070
rect 1244 1008 1278 1070
rect -1278 -1070 -1244 -1008
rect 1244 -1070 1278 -1008
rect -1278 -1104 -1182 -1070
rect 1182 -1104 1278 -1070
<< viali >>
rect -1132 559 -1094 956
rect -814 559 -776 956
rect -496 559 -458 956
rect -178 559 -140 956
rect 140 559 178 956
rect 458 559 496 956
rect 776 559 814 956
rect 1094 559 1132 956
rect -1132 -956 -1094 -559
rect -814 -956 -776 -559
rect -496 -956 -458 -559
rect -178 -956 -140 -559
rect 140 -956 178 -559
rect 458 -956 496 -559
rect 776 -956 814 -559
rect 1094 -956 1132 -559
<< metal1 >>
rect -1138 956 -1088 968
rect -1138 559 -1132 956
rect -1094 559 -1088 956
rect -1138 547 -1088 559
rect -820 956 -770 968
rect -820 559 -814 956
rect -776 559 -770 956
rect -820 547 -770 559
rect -502 956 -452 968
rect -502 559 -496 956
rect -458 559 -452 956
rect -502 547 -452 559
rect -184 956 -134 968
rect -184 559 -178 956
rect -140 559 -134 956
rect -184 547 -134 559
rect 134 956 184 968
rect 134 559 140 956
rect 178 559 184 956
rect 134 547 184 559
rect 452 956 502 968
rect 452 559 458 956
rect 496 559 502 956
rect 452 547 502 559
rect 770 956 820 968
rect 770 559 776 956
rect 814 559 820 956
rect 770 547 820 559
rect 1088 956 1138 968
rect 1088 559 1094 956
rect 1132 559 1138 956
rect 1088 547 1138 559
rect -1138 -559 -1088 -547
rect -1138 -956 -1132 -559
rect -1094 -956 -1088 -559
rect -1138 -968 -1088 -956
rect -820 -559 -770 -547
rect -820 -956 -814 -559
rect -776 -956 -770 -559
rect -820 -968 -770 -956
rect -502 -559 -452 -547
rect -502 -956 -496 -559
rect -458 -956 -452 -559
rect -502 -968 -452 -956
rect -184 -559 -134 -547
rect -184 -956 -178 -559
rect -140 -956 -134 -559
rect -184 -968 -134 -956
rect 134 -559 184 -547
rect 134 -956 140 -559
rect 178 -956 184 -559
rect 134 -968 184 -956
rect 452 -559 502 -547
rect 452 -956 458 -559
rect 496 -956 502 -559
rect 452 -968 502 -956
rect 770 -559 820 -547
rect 770 -956 776 -559
rect 814 -956 820 -559
rect 770 -968 820 -956
rect 1088 -559 1138 -547
rect 1088 -956 1094 -559
rect 1132 -956 1138 -559
rect 1088 -968 1138 -956
<< res0p35 >>
rect -1150 -544 -1076 544
rect -832 -544 -758 544
rect -514 -544 -440 544
rect -196 -544 -122 544
rect 122 -544 196 544
rect 440 -544 514 544
rect 758 -544 832 544
rect 1076 -544 1150 544
<< properties >>
string FIXED_BBOX -1261 -1087 1261 1087
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 5.42 m 1 nx 8 wmin 0.350 lmin 0.50 rho 2000 val 32.046k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
