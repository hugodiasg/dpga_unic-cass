magic
tech sky130A
timestamp 1698530758
<< metal1 >>
rect -100 9920 0 9940
rect -100 9875 145 9920
rect 160 9875 2480 9920
rect -100 9845 0 9875
rect -100 9650 0 9680
rect -100 9600 2480 9650
rect -100 9585 0 9600
rect 375 5080 2650 5100
rect 375 5010 2580 5080
rect 2630 5010 2650 5080
rect 375 5000 2650 5010
rect 3600 5075 3700 5100
rect 375 4600 475 5000
rect 3600 4990 3620 5075
rect 3685 4990 3700 5075
rect 3600 4850 3700 4990
rect 2015 4750 3700 4850
rect 4650 5095 4750 5150
rect 4650 5010 4670 5095
rect 4735 5010 4750 5095
rect 2015 4600 2115 4750
rect 4650 4700 4750 5010
rect 5700 5095 5800 5150
rect 5700 5010 5715 5095
rect 5780 5010 5800 5095
rect 5700 4725 5800 5010
rect 6750 5095 7105 5100
rect 6750 5010 6800 5095
rect 6865 5010 7105 5095
rect 6750 5000 7105 5010
rect 3630 4600 4750 4700
rect 5250 4625 5800 4725
rect 7005 4625 7105 5000
rect 7850 5095 7950 5150
rect 7850 5010 7860 5095
rect 7925 5010 7950 5095
rect 7850 4725 7950 5010
rect 8850 5090 9350 5100
rect 8850 5005 8905 5090
rect 8970 5005 9350 5090
rect 8850 5000 9350 5005
rect 9950 5095 12455 5100
rect 9950 5010 9970 5095
rect 10035 5010 12455 5095
rect 9950 5000 12455 5010
rect 9250 4725 9350 5000
rect 7850 4625 8875 4725
rect 9250 4625 10690 4725
rect 12355 4600 12455 5000
rect 14600 4720 14700 4820
rect 17715 2895 17815 2995
rect -100 1720 0 1820
rect -100 1250 0 1350
rect 7025 -80 7125 20
rect 14350 -100 14450 0
<< rmetal1 >>
rect 145 9875 160 9920
<< via1 >>
rect 2580 5010 2630 5080
rect 3620 4990 3685 5075
rect 4670 5010 4735 5095
rect 5715 5010 5780 5095
rect 6800 5010 6865 5095
rect 7860 5010 7925 5095
rect 8905 5005 8970 5090
rect 9970 5010 10035 5095
<< metal2 >>
rect 3000 14755 3100 14850
rect 5160 14735 5260 14830
rect 7325 14735 7425 14830
rect 9490 14735 9590 14830
rect 4670 5095 4735 5100
rect 2570 5080 2630 5090
rect 2570 5010 2580 5080
rect 2570 5005 2630 5010
rect 3620 5075 3685 5080
rect 4670 5005 4735 5010
rect 5715 5095 5780 5100
rect 5715 5005 5780 5010
rect 6800 5095 6865 5100
rect 6800 5005 6865 5010
rect 7860 5095 7925 5100
rect 9970 5095 10035 5100
rect 7860 5005 7925 5010
rect 8905 5090 8970 5095
rect 9970 5005 10035 5010
rect 8905 5000 8970 5005
rect 3620 4985 3685 4990
use ota_digpot  ota_digpot_0 /foss/designs/projects/dpga2/magic/ota_digpot
timestamp 1698525607
transform 1 0 100 0 1 245
box -100 -245 17615 4480
use sr  sr_0 /foss/designs/projects/dpga2/magic/spi
timestamp 1698499480
transform -1 0 10662 0 1 5000
box 528 0 8212 9828
<< labels >>
flabel space 14350 0 14450 95 0 FreeSans 800 0 0 0 inp
port 3 nsew
flabel metal2 3000 14755 3100 14850 0 FreeSans 800 0 0 0 reset
port 6 nsew
flabel metal2 5160 14735 5260 14830 0 FreeSans 800 0 0 0 sdi
port 7 nsew
flabel metal1 -100 1720 0 1820 0 FreeSans 800 0 0 0 vd
port 14 nsew
flabel metal1 -100 1250 0 1350 0 FreeSans 800 0 0 0 gnd
port 5 nsew
flabel metal1 7025 -80 7125 20 0 FreeSans 800 0 0 0 inn
port 15 nsew
flabel metal1 14350 -100 14450 0 0 FreeSans 800 0 0 0 inp
port 16 nsew
flabel metal1 17715 2895 17815 2995 0 FreeSans 800 0 0 0 out
port 17 nsew
flabel metal1 14600 4720 14700 4820 0 FreeSans 800 0 0 0 ib
port 18 nsew
flabel metal1 -100 9845 0 9940 0 FreeSans 800 0 0 0 gndd
port 9 nsew
flabel metal2 7325 14735 7425 14830 0 FreeSans 800 0 0 0 sclk
port 19 nsew
flabel metal2 9490 14735 9590 14830 0 FreeSans 800 0 0 0 ss
port 21 nsew
flabel metal1 -100 9585 0 9680 0 FreeSans 800 0 0 0 vpwr
port 11 nsew
flabel metal1 709 9885 754 9894 0 FreeSans 800 0 0 0 vgnd
<< end >>
