magic
tech sky130A
magscale 1 2
timestamp 1698520465
<< nwell >>
rect -500 2100 1700 3660
<< pwell >>
rect -500 580 1680 2100
<< psubdiff >>
rect -470 2040 1660 2070
rect -470 660 -440 2040
rect -400 2000 -360 2040
rect 1560 2030 1660 2040
rect 1560 2000 1600 2030
rect -400 1980 1600 2000
rect -400 710 -380 1980
rect 1580 710 1600 1980
rect -400 680 1600 710
rect -400 660 -360 680
rect -470 640 -360 660
rect 1560 650 1600 680
rect 1640 650 1660 2030
rect 1560 640 1660 650
rect -470 620 1660 640
<< nsubdiff >>
rect -460 3600 1660 3620
rect -460 3580 -360 3600
rect -460 2180 -440 3580
rect -400 3560 -360 3580
rect 1560 3580 1660 3600
rect 1560 3560 1600 3580
rect -400 3540 1600 3560
rect -400 2240 -380 3540
rect -400 2220 -360 2240
rect 1580 2220 1600 3540
rect -400 2200 1600 2220
rect -400 2180 -360 2200
rect -460 2160 -360 2180
rect 1560 2180 1600 2200
rect 1640 2180 1660 3580
rect 1560 2160 1660 2180
rect -460 2140 1660 2160
<< psubdiffcont >>
rect -440 660 -400 2040
rect -360 2000 1560 2040
rect -360 640 1560 680
rect 1600 650 1640 2030
<< nsubdiffcont >>
rect -440 2180 -400 3580
rect -360 3560 1560 3600
rect -360 2160 1560 2200
rect 1600 2180 1640 3580
<< poly >>
rect 150 3400 1240 3450
rect 150 3380 184 3400
rect 343 3363 373 3400
rect 535 3363 565 3400
rect 727 3363 757 3400
rect 919 3385 949 3400
rect 919 3363 945 3385
rect 1111 3380 1141 3400
rect 150 819 1146 820
rect 150 810 1158 819
rect 1211 810 1241 817
rect 150 760 1241 810
rect 150 750 1240 760
<< locali >>
rect -460 3600 1660 3620
rect -460 3580 -360 3600
rect -460 2180 -440 3580
rect -400 3560 -360 3580
rect 1560 3580 1660 3600
rect 1560 3560 1600 3580
rect -400 3540 1600 3560
rect -400 2720 -380 3540
rect -390 2630 -380 2720
rect -400 2240 -380 2630
rect -400 2220 -360 2240
rect 1580 2220 1600 3540
rect -400 2200 1600 2220
rect -400 2180 -360 2200
rect -460 2160 -360 2180
rect 1560 2180 1600 2200
rect 1640 2180 1660 3580
rect 1560 2160 1660 2180
rect -460 2140 1660 2160
rect -470 2040 1660 2070
rect -470 1810 -440 2040
rect -400 2000 -360 2040
rect 1560 2030 1660 2040
rect 1560 2000 1600 2030
rect -400 1980 1600 2000
rect -400 1810 -380 1980
rect -470 1680 -450 1810
rect -390 1680 -380 1810
rect -470 660 -440 1680
rect -400 710 -380 1680
rect 1580 710 1600 1980
rect -400 680 1600 710
rect -400 660 -360 680
rect -470 640 -360 660
rect 1560 650 1600 680
rect 1640 650 1660 2030
rect 1560 640 1660 650
rect -470 620 1660 640
<< viali >>
rect -440 2630 -400 2720
rect -400 2630 -390 2720
rect -450 1680 -440 1810
rect -440 1680 -400 1810
rect -400 1680 -390 1810
<< metal1 >>
rect -280 3450 -220 3470
rect -300 3320 -180 3450
rect 10 3410 1260 3470
rect 1420 3410 1480 3470
rect -80 3010 -20 3070
rect -700 2730 -500 2780
rect -230 2730 -90 2960
rect 10 2860 50 3410
rect 110 3190 1270 3340
rect 110 3090 140 3190
rect 280 3090 1270 3190
rect 110 3030 1270 3090
rect 100 2960 1270 3030
rect 100 2950 140 2960
rect 130 2930 140 2950
rect -700 2720 -90 2730
rect -700 2630 -440 2720
rect -390 2630 -90 2720
rect -700 2620 -90 2630
rect -700 2580 -500 2620
rect -230 2390 -90 2620
rect -300 2270 -220 2330
rect -700 1820 -500 1840
rect -310 1820 -190 1940
rect -80 1880 -20 2330
rect -700 1810 -90 1820
rect -700 1680 -450 1810
rect -390 1680 -90 1810
rect 10 1740 40 2520
rect 180 2480 1330 2690
rect 180 2410 1540 2480
rect 1230 2400 1540 2410
rect 150 2270 1160 2330
rect 1300 2240 1540 2400
rect 1700 2240 1900 2340
rect 1300 2140 1900 2240
rect 240 1880 1260 1940
rect 1300 1830 1330 2140
rect 1400 1870 1470 1940
rect 1260 1820 1330 1830
rect -700 1670 -90 1680
rect -700 1640 -500 1670
rect -330 1660 -190 1670
rect -80 1560 -20 1620
rect 120 1610 1330 1820
rect -700 1115 -500 1200
rect -70 1115 -20 1560
rect -700 1065 -20 1115
rect 170 1240 1200 1260
rect 170 1140 180 1240
rect 290 1140 1200 1240
rect 170 1120 1200 1140
rect -700 1000 -500 1065
rect -280 770 -220 830
rect -75 815 -25 1065
rect 170 1020 180 1120
rect 290 1020 1200 1120
rect 170 1010 1200 1020
rect 1700 1010 1900 1060
rect 170 1000 1900 1010
rect 170 900 180 1000
rect 290 930 1900 1000
rect 290 900 1200 930
rect 170 870 1200 900
rect -75 800 155 815
rect -75 765 1160 800
rect 1360 770 1500 930
rect 1700 860 1900 930
rect 140 740 1160 765
rect 1400 760 1460 770
<< via1 >>
rect 140 3090 280 3190
rect 180 1140 290 1240
rect 180 1020 290 1120
rect 180 900 290 1000
<< metal2 >>
rect 120 3190 300 3200
rect 120 3090 140 3190
rect 280 3090 300 3190
rect 120 3080 300 3090
rect 170 1260 250 3080
rect 170 1240 300 1260
rect 170 1140 180 1240
rect 290 1140 300 1240
rect 170 1120 300 1140
rect 170 1020 180 1120
rect 290 1020 300 1120
rect 170 1000 300 1020
rect 170 900 180 1000
rect 290 900 300 1000
rect 170 870 300 900
use sky130_fd_pr__pfet_01v8_8QR85J  XM2
timestamp 1698518340
transform 1 0 -251 0 1 2870
box -109 -600 109 600
use sky130_fd_pr__nfet_01v8_4W7PEP  XM3
timestamp 1698517357
transform 1 0 -47 0 1 1748
box -73 -188 73 188
use sky130_fd_pr__pfet_01v8_XGAKDL  XM4
timestamp 1698517357
transform 1 0 -51 0 1 2670
box -109 -400 109 400
use sky130_fd_pr__nfet_01v8_ECDJHW  sky130_fd_pr__nfet_01v8_ECDJHW_0
timestamp 1698517357
transform 1 0 698 0 1 1341
box -605 -588 605 588
use sky130_fd_pr__nfet_01v8_VQ5UWM  sky130_fd_pr__nfet_01v8_VQ5UWM_1
timestamp 1698518340
transform 1 0 -247 0 1 1348
box -73 -588 73 588
use sky130_fd_pr__nfet_01v8_VU5CXM  sky130_fd_pr__nfet_01v8_VU5CXM_0
timestamp 1698518638
transform 1 0 1433 0 1 1348
box -73 -588 73 588
use sky130_fd_pr__pfet_01v8_PM4G2P  sky130_fd_pr__pfet_01v8_PM4G2P_0
timestamp 1698517357
transform 1 0 694 0 1 2863
box -641 -600 641 600
use sky130_fd_pr__pfet_01v8_UGA66J  sky130_fd_pr__pfet_01v8_UGA66J_0
timestamp 1698517357
transform 1 0 1449 0 1 2870
box -109 -600 109 600
<< labels >>
flabel metal1 -700 2580 -500 2780 0 FreeSans 256 0 0 0 vd
port 0 nsew
flabel metal1 1700 2140 1900 2340 0 FreeSans 256 0 0 0 b
port 2 nsew
flabel metal1 -700 1640 -500 1840 0 FreeSans 256 0 0 0 vgnd
port 1 nsew
flabel metal1 -700 1000 -500 1200 0 FreeSans 256 0 0 0 ctrl
port 4 nsew
flabel metal1 1700 860 1900 1060 0 FreeSans 256 0 0 0 a
port 3 nsew
flabel metal1 20 3400 40 3410 0 FreeSans 1600 0 0 0 nctrl
<< end >>
