magic
tech sky130A
magscale 1 2
timestamp 1698525106
<< nwell >>
rect 5120 3820 10480 6060
<< pwell >>
rect 5120 2880 10480 3810
<< psubdiff >>
rect 5160 3760 10400 3780
rect 5160 3720 5260 3760
rect 10300 3740 10400 3760
rect 10300 3720 10340 3740
rect 5160 3700 10340 3720
rect 5160 3060 5180 3700
rect 5220 3060 5240 3700
rect 10320 3080 10340 3700
rect 10380 3080 10400 3740
rect 10320 3060 10400 3080
rect 5160 3040 10400 3060
rect 5160 3000 5260 3040
rect 10320 3000 10400 3040
rect 5160 2980 10400 3000
<< nsubdiff >>
rect 5180 6000 10440 6020
rect 5180 5960 5280 6000
rect 10360 5960 10440 6000
rect 5180 5940 10440 5960
rect 5180 3920 5200 5940
rect 5240 3940 5260 5940
rect 10360 5920 10440 5940
rect 10360 3980 10380 5920
rect 10420 3980 10440 5920
rect 10360 3940 10440 3980
rect 5240 3920 10440 3940
rect 5180 3880 5280 3920
rect 10380 3880 10440 3920
rect 5180 3860 10440 3880
<< psubdiffcont >>
rect 5260 3720 10300 3760
rect 5180 3060 5220 3700
rect 10340 3080 10380 3740
rect 5260 3000 10320 3040
<< nsubdiffcont >>
rect 5280 5960 10360 6000
rect 5200 3920 5240 5940
rect 10380 3980 10420 5920
rect 5280 3880 10380 3920
<< poly >>
rect 5890 3990 6120 4060
rect 6280 4000 6540 4060
<< locali >>
rect 5180 6000 10440 6020
rect 5180 5960 5280 6000
rect 10360 5960 10440 6000
rect 5180 5940 10440 5960
rect 5180 3920 5200 5940
rect 5240 3940 5260 5940
rect 10360 5920 10440 5940
rect 10360 3980 10380 5920
rect 10420 3980 10440 5920
rect 10360 3940 10440 3980
rect 5240 3920 10440 3940
rect 5180 3880 5280 3920
rect 10380 3880 10440 3920
rect 5180 3860 10440 3880
rect 5160 3760 10400 3780
rect 5160 3720 5260 3760
rect 10300 3740 10400 3760
rect 10300 3720 10340 3740
rect 5160 3700 10340 3720
rect 5160 3060 5180 3700
rect 5220 3060 5240 3700
rect 10320 3080 10340 3700
rect 10380 3080 10400 3740
rect 10320 3060 10400 3080
rect 5160 3040 10400 3060
rect 5160 3000 5260 3040
rect 10320 3000 10400 3040
rect 5160 2980 10400 3000
<< viali >>
rect 5380 5960 5980 6000
rect 5500 3000 5760 3040
<< metal1 >>
rect 7650 6120 7850 6320
rect 7700 6020 7820 6120
rect 5320 6000 10280 6020
rect 5320 5960 5380 6000
rect 5980 5960 10280 6000
rect 5320 5940 10280 5960
rect 5320 5900 10290 5940
rect 5360 5620 5650 5900
rect 5720 5640 5760 5900
rect 6360 5660 6400 5900
rect 7260 5660 7300 5900
rect 5720 5520 6300 5640
rect 6360 5540 6960 5660
rect 7260 5560 9900 5660
rect 9980 5580 10290 5900
rect 9430 5310 9560 5330
rect 6640 5240 7200 5280
rect 9430 5250 9450 5310
rect 4800 5060 5000 5140
rect 6000 5060 6040 5220
rect 6640 5160 6860 5240
rect 6940 5160 7200 5240
rect 6640 5120 7200 5160
rect 7520 5150 9450 5250
rect 9550 5250 9560 5310
rect 9550 5150 9640 5250
rect 7520 5140 9640 5150
rect 4800 5000 5370 5060
rect 4800 4940 5000 5000
rect 5310 4980 5370 5000
rect 5670 5000 9880 5060
rect 5670 4980 5730 5000
rect 5310 4920 5730 4980
rect 5070 4820 6040 4890
rect 4810 4640 5010 4710
rect 5070 4640 5120 4820
rect 5660 4770 5720 4780
rect 4810 4570 5120 4640
rect 5620 4620 5750 4770
rect 5970 4730 6040 4820
rect 5980 4720 6040 4730
rect 6160 4880 6260 4900
rect 10630 4880 10830 4950
rect 6160 4800 6180 4880
rect 6240 4800 6260 4880
rect 6160 4640 6260 4800
rect 10505 4860 10830 4880
rect 10505 4780 10520 4860
rect 10610 4780 10830 4860
rect 6380 4720 6440 4780
rect 6680 4760 6740 4780
rect 10505 4770 10830 4780
rect 5860 4630 6560 4640
rect 6670 4630 6750 4760
rect 10630 4750 10830 4770
rect 5860 4620 6780 4630
rect 5620 4610 6780 4620
rect 4810 4510 5010 4570
rect 5720 4500 6780 4610
rect 5860 4480 6780 4500
rect 5960 4100 6160 4240
rect 5660 3980 5720 4040
rect 5880 3980 5940 4040
rect 4810 3820 5010 3870
rect 5080 3820 5160 3830
rect 4810 3770 5090 3820
rect 4810 3670 5010 3770
rect 5080 3760 5090 3770
rect 5150 3760 5160 3820
rect 5980 3780 6020 4100
rect 6260 4080 6480 4240
rect 6080 3980 6140 4040
rect 6270 4030 6350 4040
rect 6270 3970 6280 4030
rect 6340 3970 6350 4030
rect 6270 3960 6350 3970
rect 5080 3750 5160 3760
rect 5820 3740 6020 3780
rect 6380 3780 6420 4080
rect 6480 3980 6540 4040
rect 6680 3980 6740 4040
rect 6380 3740 6580 3780
rect 5820 3580 5860 3740
rect 6540 3590 6580 3740
rect 5820 3540 6500 3580
rect 6540 3550 8940 3590
rect 5820 3480 5860 3540
rect 6540 3510 6580 3550
rect 5470 3040 5770 3400
rect 5840 3340 5880 3480
rect 6120 3400 6280 3500
rect 6100 3360 6280 3400
rect 6120 3300 6280 3360
rect 4800 2990 5000 3030
rect 5470 3000 5500 3040
rect 5760 3000 5770 3040
rect 5470 2990 5770 3000
rect 6180 2990 6220 3300
rect 6530 3170 6590 3510
rect 6640 3490 8740 3510
rect 6640 3470 8550 3490
rect 8540 3410 8550 3470
rect 8630 3470 8740 3490
rect 8630 3410 8640 3470
rect 8540 3400 8640 3410
rect 6880 3310 9000 3350
rect 6500 3160 6650 3170
rect 6500 3040 6520 3160
rect 6640 3040 6650 3160
rect 6500 3030 6650 3040
rect 8970 2990 9000 3310
rect 9070 3200 9360 3350
rect 9050 3120 9360 3200
rect 9050 2990 9350 3120
rect 4800 2870 9350 2990
rect 4800 2830 5000 2870
<< via1 >>
rect 6860 5160 6940 5240
rect 9450 5150 9550 5310
rect 6180 4800 6240 4880
rect 10520 4780 10610 4860
rect 5090 3760 5150 3820
rect 6280 3970 6340 4030
rect 8550 3410 8630 3490
rect 6520 3040 6640 3160
<< metal2 >>
rect 9430 5310 9560 5330
rect 6840 5240 6960 5260
rect 6840 5160 6860 5240
rect 6940 5160 6960 5240
rect 6840 5140 6960 5160
rect 9430 5150 9450 5310
rect 9550 5150 9560 5310
rect 9430 5140 9560 5150
rect 6860 4900 6940 5140
rect 6160 4880 6940 4900
rect 9440 4880 9550 5140
rect 6160 4800 6180 4880
rect 6240 4820 6940 4880
rect 8535 4860 10615 4880
rect 6240 4800 6260 4820
rect 6160 4780 6260 4800
rect 8535 4780 10520 4860
rect 10610 4780 10615 4860
rect 8535 4770 10615 4780
rect 6270 4030 6350 4040
rect 6270 3970 6280 4030
rect 6340 3970 6350 4030
rect 6270 3960 6350 3970
rect 5080 3820 5160 3830
rect 6290 3820 6340 3960
rect 5080 3760 5090 3820
rect 5150 3770 6340 3820
rect 5150 3760 5160 3770
rect 5080 3750 5160 3760
rect 8535 3490 8645 4770
rect 8535 3410 8550 3490
rect 8630 3410 8645 3490
rect 8535 3365 8645 3410
rect 6500 3160 6650 3170
rect 6500 3040 6520 3160
rect 6640 3040 6650 3160
rect 8540 3150 8640 3365
rect 8540 3050 8550 3150
rect 8630 3050 8640 3150
rect 8540 3040 8640 3050
rect 6500 3030 6650 3040
<< via2 >>
rect 6520 3040 6640 3160
rect 8550 3050 8630 3150
<< metal3 >>
rect 6500 3160 6650 3170
rect 6500 3040 6520 3160
rect 6640 3040 6650 3160
rect 8540 3150 8640 3160
rect 8540 3050 8550 3150
rect 8630 3050 8640 3150
rect 8540 3040 8640 3050
rect 6500 3030 6650 3040
<< via3 >>
rect 6520 3040 6640 3160
rect 8550 3050 8630 3150
<< metal4 >>
rect 6500 3160 6650 3170
rect 6500 3040 6520 3160
rect 6640 3040 6650 3160
rect 6500 2990 6650 3040
rect 5265 2900 6650 2990
rect 8540 3150 8640 3160
rect 8540 3050 8550 3150
rect 8630 3050 8640 3150
rect 5265 2625 5400 2900
rect 8540 2530 8640 3050
use sky130_fd_pr__cap_mim_m3_1_VTBF8H  XCC
timestamp 1698511094
transform -1 0 7869 0 1 1340
box -2550 -1500 2549 1500
use sky130_fd_pr__nfet_01v8_UFMA4B  XM3
timestamp 1698511094
transform 1 0 5618 0 1 3408
box -158 -188 158 188
use sky130_fd_pr__pfet_01v8_FRJNPM  XM6
timestamp 1698511094
transform 1 0 6792 0 1 5400
box -452 -400 452 400
use sky130_fd_pr__nfet_01v8_Q7RUWS  XM7
timestamp 1698513452
transform 1 0 7810 0 1 3408
box -1190 -188 1190 188
use sky130_fd_pr__pfet_01v8_WM6J89  XM8
timestamp 1698511094
transform 1 0 8595 0 1 5400
box -1355 -400 1355 400
use sky130_fd_pr__pfet_01v8_3HT9FS  XPD1
timestamp 1698511094
transform 1 0 5514 0 1 5400
box -194 -400 194 400
use sky130_fd_pr__nfet_01v8_UFMA4B  sky130_fd_pr__nfet_01v8_UFMA4B_0
timestamp 1698511094
transform 1 0 6398 0 1 3408
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_UFMA4B  sky130_fd_pr__nfet_01v8_UFMA4B_1
timestamp 1698511094
transform 1 0 5998 0 1 3408
box -158 -188 158 188
use sky130_fd_pr__nfet_01v8_UFMA4B  sky130_fd_pr__nfet_01v8_UFMA4B_2
timestamp 1698511094
transform 1 0 9218 0 1 3408
box -158 -188 158 188
use sky130_fd_pr__pfet_01v8_3HT9FS  sky130_fd_pr__pfet_01v8_3HT9FS_0
timestamp 1698511094
transform 1 0 10134 0 1 5400
box -194 -400 194 400
use sky130_fd_pr__pfet_01v8_FRN4QM  sky130_fd_pr__pfet_01v8_FRN4QM_0
timestamp 1698511094
transform 1 0 6023 0 1 5400
box -323 -400 323 400
use sky130_fd_pr__pfet_01v8_KRRM6L  sky130_fd_pr__pfet_01v8_KRRM6L_0
timestamp 1698525106
transform 1 0 6709 0 1 4380
box -109 -400 109 400
use sky130_fd_pr__pfet_01v8_KRRM6L  sky130_fd_pr__pfet_01v8_KRRM6L_1
timestamp 1698525106
transform 1 0 5689 0 1 4380
box -109 -400 109 400
use sky130_fd_pr__pfet_01v8_KRZE7L  sky130_fd_pr__pfet_01v8_KRZE7L_1
timestamp 1698511094
transform 1 0 6009 0 1 4380
box -209 -400 209 400
use sky130_fd_pr__pfet_01v8_KVZW6L  sky130_fd_pr__pfet_01v8_KVZW6L_0
timestamp 1698513452
transform 1 0 6409 0 1 4380
box -209 -400 209 400
<< labels >>
flabel metal1 4800 2830 5000 3030 0 FreeSans 256 0 0 0 vs
port 1 nsew
flabel metal1 4810 4510 5010 4710 0 FreeSans 256 0 0 0 inn
port 3 nsew
flabel metal1 4810 3670 5010 3870 0 FreeSans 256 0 0 0 inp
port 4 nsew
flabel metal1 4800 4940 5000 5140 0 FreeSans 256 0 0 0 ib
port 2 nsew
flabel metal1 7650 6120 7850 6320 0 FreeSans 256 0 0 0 vd
port 0 nsew
flabel metal1 10630 4750 10830 4950 0 FreeSans 256 0 0 0 out
port 5 nsew
flabel metal1 6540 3640 6580 3660 0 FreeSans 1600 0 0 0 d
flabel metal1 5840 3640 5840 3660 0 FreeSans 1600 0 0 0 c
flabel metal2 6360 4860 6380 4880 0 FreeSans 1600 0 0 0 b
<< end >>
