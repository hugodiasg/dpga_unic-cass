magic
tech sky130A
magscale 1 2
timestamp 1698520721
<< pwell >>
rect -201 -720 201 720
<< psubdiff >>
rect -165 650 -69 684
rect 69 650 165 684
rect -165 588 -131 650
rect 131 588 165 650
rect -165 -650 -131 -588
rect 131 -650 165 -588
rect -165 -684 -69 -650
rect 69 -684 165 -650
<< psubdiffcont >>
rect -69 650 69 684
rect -165 -588 -131 588
rect 131 -588 165 588
rect -69 -684 69 -650
<< xpolycontact >>
rect -35 122 35 554
rect -35 -554 35 -122
<< xpolyres >>
rect -35 -122 35 122
<< locali >>
rect -165 650 -69 684
rect 69 650 165 684
rect -165 588 -131 650
rect 131 588 165 650
rect -165 -650 -131 -588
rect 131 -650 165 -588
rect -165 -684 -69 -650
rect 69 -684 165 -650
<< viali >>
rect -19 139 19 536
rect -19 -536 19 -139
<< metal1 >>
rect -25 536 25 548
rect -25 139 -19 536
rect 19 139 25 536
rect -25 127 25 139
rect -25 -139 25 -127
rect -25 -536 -19 -139
rect 19 -536 25 -139
rect -25 -548 25 -536
<< res0p35 >>
rect -37 -124 37 124
<< properties >>
string FIXED_BBOX -148 -667 148 667
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 1.22 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 8.046k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
