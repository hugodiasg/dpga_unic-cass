magic
tech sky130A
magscale 1 2
timestamp 1698511094
<< nwell >>
rect -452 -400 452 400
<< pmos >>
rect -358 -300 -158 300
rect -100 -300 100 300
rect 158 -300 358 300
<< pdiff >>
rect -416 288 -358 300
rect -416 -288 -404 288
rect -370 -288 -358 288
rect -416 -300 -358 -288
rect -158 288 -100 300
rect -158 -288 -146 288
rect -112 -288 -100 288
rect -158 -300 -100 -288
rect 100 288 158 300
rect 100 -288 112 288
rect 146 -288 158 288
rect 100 -300 158 -288
rect 358 288 416 300
rect 358 -288 370 288
rect 404 -288 416 288
rect 358 -300 416 -288
<< pdiffc >>
rect -404 -288 -370 288
rect -146 -288 -112 288
rect 112 -288 146 288
rect 370 -288 404 288
<< poly >>
rect -358 381 -158 397
rect -358 347 -342 381
rect -174 347 -158 381
rect -358 300 -158 347
rect -100 381 100 397
rect -100 347 -84 381
rect 84 347 100 381
rect -100 300 100 347
rect 158 381 358 397
rect 158 347 174 381
rect 342 347 358 381
rect 158 300 358 347
rect -358 -347 -158 -300
rect -358 -381 -342 -347
rect -174 -381 -158 -347
rect -358 -397 -158 -381
rect -100 -347 100 -300
rect -100 -381 -84 -347
rect 84 -381 100 -347
rect -100 -397 100 -381
rect 158 -347 358 -300
rect 158 -381 174 -347
rect 342 -381 358 -347
rect 158 -397 358 -381
<< polycont >>
rect -342 347 -174 381
rect -84 347 84 381
rect 174 347 342 381
rect -342 -381 -174 -347
rect -84 -381 84 -347
rect 174 -381 342 -347
<< locali >>
rect -358 347 -342 381
rect -174 347 -158 381
rect -100 347 -84 381
rect 84 347 100 381
rect 158 347 174 381
rect 342 347 358 381
rect -404 288 -370 304
rect -404 -304 -370 -288
rect -146 288 -112 304
rect -146 -304 -112 -288
rect 112 288 146 304
rect 112 -304 146 -288
rect 370 288 404 304
rect 370 -304 404 -288
rect -358 -381 -342 -347
rect -174 -381 -158 -347
rect -100 -381 -84 -347
rect 84 -381 100 -347
rect 158 -381 174 -347
rect 342 -381 358 -347
<< viali >>
rect -342 347 -174 381
rect -84 347 84 381
rect 174 347 342 381
rect -404 -17 -370 271
rect -146 -271 -112 17
rect 112 -17 146 271
rect 370 -271 404 17
rect -342 -381 -174 -347
rect -84 -381 84 -347
rect 174 -381 342 -347
<< metal1 >>
rect -354 381 -162 387
rect -354 347 -342 381
rect -174 347 -162 381
rect -354 341 -162 347
rect -96 381 96 387
rect -96 347 -84 381
rect 84 347 96 381
rect -96 341 96 347
rect 162 381 354 387
rect 162 347 174 381
rect 342 347 354 381
rect 162 341 354 347
rect -410 271 -364 283
rect -410 -17 -404 271
rect -370 -17 -364 271
rect 106 271 152 283
rect -410 -29 -364 -17
rect -152 17 -106 29
rect -152 -271 -146 17
rect -112 -271 -106 17
rect 106 -17 112 271
rect 146 -17 152 271
rect 106 -29 152 -17
rect 364 17 410 29
rect -152 -283 -106 -271
rect 364 -271 370 17
rect 404 -271 410 17
rect 364 -283 410 -271
rect -354 -347 -162 -341
rect -354 -381 -342 -347
rect -174 -381 -162 -347
rect -354 -387 -162 -381
rect -96 -347 96 -341
rect -96 -381 -84 -347
rect 84 -381 96 -347
rect -96 -387 96 -381
rect 162 -347 354 -341
rect 162 -381 174 -347
rect 342 -381 354 -347
rect 162 -387 354 -381
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.0 l 1.0 m 1 nf 3 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc +50 viadrn -50 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
