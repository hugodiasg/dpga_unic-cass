magic
tech sky130A
magscale 1 2
timestamp 1698517357
<< error_p >>
rect -461 572 -403 578
rect -269 572 -211 578
rect -77 572 -19 578
rect 115 572 173 578
rect 307 572 365 578
rect 499 572 557 578
rect -461 538 -449 572
rect -269 538 -257 572
rect -77 538 -65 572
rect 115 538 127 572
rect 307 538 319 572
rect 499 538 511 572
rect -461 532 -403 538
rect -269 532 -211 538
rect -77 532 -19 538
rect 115 532 173 538
rect 307 532 365 538
rect 499 532 557 538
rect -557 -538 -499 -532
rect -365 -538 -307 -532
rect -173 -538 -115 -532
rect 19 -538 77 -532
rect 211 -538 269 -532
rect 403 -538 461 -532
rect -557 -572 -545 -538
rect -365 -572 -353 -538
rect -173 -572 -161 -538
rect 19 -572 31 -538
rect 211 -572 223 -538
rect 403 -572 415 -538
rect -557 -578 -499 -572
rect -365 -578 -307 -572
rect -173 -578 -115 -572
rect 19 -578 77 -572
rect 211 -578 269 -572
rect 403 -578 461 -572
<< nmos >>
rect -543 -500 -513 500
rect -447 -500 -417 500
rect -351 -500 -321 500
rect -255 -500 -225 500
rect -159 -500 -129 500
rect -63 -500 -33 500
rect 33 -500 63 500
rect 129 -500 159 500
rect 225 -500 255 500
rect 321 -500 351 500
rect 417 -500 447 500
rect 513 -500 543 500
<< ndiff >>
rect -605 488 -543 500
rect -605 -488 -593 488
rect -559 -488 -543 488
rect -605 -500 -543 -488
rect -513 488 -447 500
rect -513 -488 -497 488
rect -463 -488 -447 488
rect -513 -500 -447 -488
rect -417 488 -351 500
rect -417 -488 -401 488
rect -367 -488 -351 488
rect -417 -500 -351 -488
rect -321 488 -255 500
rect -321 -488 -305 488
rect -271 -488 -255 488
rect -321 -500 -255 -488
rect -225 488 -159 500
rect -225 -488 -209 488
rect -175 -488 -159 488
rect -225 -500 -159 -488
rect -129 488 -63 500
rect -129 -488 -113 488
rect -79 -488 -63 488
rect -129 -500 -63 -488
rect -33 488 33 500
rect -33 -488 -17 488
rect 17 -488 33 488
rect -33 -500 33 -488
rect 63 488 129 500
rect 63 -488 79 488
rect 113 -488 129 488
rect 63 -500 129 -488
rect 159 488 225 500
rect 159 -488 175 488
rect 209 -488 225 488
rect 159 -500 225 -488
rect 255 488 321 500
rect 255 -488 271 488
rect 305 -488 321 488
rect 255 -500 321 -488
rect 351 488 417 500
rect 351 -488 367 488
rect 401 -488 417 488
rect 351 -500 417 -488
rect 447 488 513 500
rect 447 -488 463 488
rect 497 -488 513 488
rect 447 -500 513 -488
rect 543 488 605 500
rect 543 -488 559 488
rect 593 -488 605 488
rect 543 -500 605 -488
<< ndiffc >>
rect -593 -488 -559 488
rect -497 -488 -463 488
rect -401 -488 -367 488
rect -305 -488 -271 488
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
rect 271 -488 305 488
rect 367 -488 401 488
rect 463 -488 497 488
rect 559 -488 593 488
<< poly >>
rect -465 572 -399 588
rect -465 538 -449 572
rect -415 538 -399 572
rect -543 500 -513 526
rect -465 522 -399 538
rect -273 572 -207 588
rect -273 538 -257 572
rect -223 538 -207 572
rect -447 500 -417 522
rect -351 500 -321 526
rect -273 522 -207 538
rect -81 572 -15 588
rect -81 538 -65 572
rect -31 538 -15 572
rect -255 500 -225 522
rect -159 500 -129 526
rect -81 522 -15 538
rect 111 572 177 588
rect 111 538 127 572
rect 161 538 177 572
rect -63 500 -33 522
rect 33 500 63 526
rect 111 522 177 538
rect 303 572 369 588
rect 303 538 319 572
rect 353 538 369 572
rect 129 500 159 522
rect 225 500 255 526
rect 303 522 369 538
rect 495 572 561 588
rect 495 538 511 572
rect 545 538 561 572
rect 321 500 351 522
rect 417 500 447 526
rect 495 522 561 538
rect 513 500 543 522
rect -543 -522 -513 -500
rect -561 -538 -495 -522
rect -447 -526 -417 -500
rect -351 -522 -321 -500
rect -561 -572 -545 -538
rect -511 -572 -495 -538
rect -561 -588 -495 -572
rect -369 -538 -303 -522
rect -255 -526 -225 -500
rect -159 -522 -129 -500
rect -369 -572 -353 -538
rect -319 -572 -303 -538
rect -369 -588 -303 -572
rect -177 -538 -111 -522
rect -63 -526 -33 -500
rect 33 -522 63 -500
rect -177 -572 -161 -538
rect -127 -572 -111 -538
rect -177 -588 -111 -572
rect 15 -538 81 -522
rect 129 -526 159 -500
rect 225 -522 255 -500
rect 15 -572 31 -538
rect 65 -572 81 -538
rect 15 -588 81 -572
rect 207 -538 273 -522
rect 321 -526 351 -500
rect 417 -522 447 -500
rect 207 -572 223 -538
rect 257 -572 273 -538
rect 207 -588 273 -572
rect 399 -538 465 -522
rect 513 -526 543 -500
rect 399 -572 415 -538
rect 449 -572 465 -538
rect 399 -588 465 -572
<< polycont >>
rect -449 538 -415 572
rect -257 538 -223 572
rect -65 538 -31 572
rect 127 538 161 572
rect 319 538 353 572
rect 511 538 545 572
rect -545 -572 -511 -538
rect -353 -572 -319 -538
rect -161 -572 -127 -538
rect 31 -572 65 -538
rect 223 -572 257 -538
rect 415 -572 449 -538
<< locali >>
rect -465 538 -449 572
rect -415 538 -399 572
rect -273 538 -257 572
rect -223 538 -207 572
rect -81 538 -65 572
rect -31 538 -15 572
rect 111 538 127 572
rect 161 538 177 572
rect 303 538 319 572
rect 353 538 369 572
rect 495 538 511 572
rect 545 538 561 572
rect -593 488 -559 504
rect -593 -504 -559 -488
rect -497 488 -463 504
rect -497 -504 -463 -488
rect -401 488 -367 504
rect -401 -504 -367 -488
rect -305 488 -271 504
rect -305 -504 -271 -488
rect -209 488 -175 504
rect -209 -504 -175 -488
rect -113 488 -79 504
rect -113 -504 -79 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 79 488 113 504
rect 79 -504 113 -488
rect 175 488 209 504
rect 175 -504 209 -488
rect 271 488 305 504
rect 271 -504 305 -488
rect 367 488 401 504
rect 367 -504 401 -488
rect 463 488 497 504
rect 463 -504 497 -488
rect 559 488 593 504
rect 559 -504 593 -488
rect -561 -572 -545 -538
rect -511 -572 -495 -538
rect -369 -572 -353 -538
rect -319 -572 -303 -538
rect -177 -572 -161 -538
rect -127 -572 -111 -538
rect 15 -572 31 -538
rect 65 -572 81 -538
rect 207 -572 223 -538
rect 257 -572 273 -538
rect 399 -572 415 -538
rect 449 -572 465 -538
<< viali >>
rect -449 538 -415 572
rect -257 538 -223 572
rect -65 538 -31 572
rect 127 538 161 572
rect 319 538 353 572
rect 511 538 545 572
rect -593 -17 -559 471
rect -497 -471 -463 17
rect -401 -17 -367 471
rect -305 -471 -271 17
rect -209 -17 -175 471
rect -113 -471 -79 17
rect -17 -17 17 471
rect 79 -471 113 17
rect 175 -17 209 471
rect 271 -471 305 17
rect 367 -17 401 471
rect 463 -471 497 17
rect 559 -17 593 471
rect -545 -572 -511 -538
rect -353 -572 -319 -538
rect -161 -572 -127 -538
rect 31 -572 65 -538
rect 223 -572 257 -538
rect 415 -572 449 -538
<< metal1 >>
rect -461 572 -403 578
rect -461 538 -449 572
rect -415 538 -403 572
rect -461 532 -403 538
rect -269 572 -211 578
rect -269 538 -257 572
rect -223 538 -211 572
rect -269 532 -211 538
rect -77 572 -19 578
rect -77 538 -65 572
rect -31 538 -19 572
rect -77 532 -19 538
rect 115 572 173 578
rect 115 538 127 572
rect 161 538 173 572
rect 115 532 173 538
rect 307 572 365 578
rect 307 538 319 572
rect 353 538 365 572
rect 307 532 365 538
rect 499 572 557 578
rect 499 538 511 572
rect 545 538 557 572
rect 499 532 557 538
rect -599 471 -553 483
rect -599 -17 -593 471
rect -559 -17 -553 471
rect -407 471 -361 483
rect -599 -29 -553 -17
rect -503 17 -457 29
rect -503 -471 -497 17
rect -463 -471 -457 17
rect -407 -17 -401 471
rect -367 -17 -361 471
rect -215 471 -169 483
rect -407 -29 -361 -17
rect -311 17 -265 29
rect -503 -483 -457 -471
rect -311 -471 -305 17
rect -271 -471 -265 17
rect -215 -17 -209 471
rect -175 -17 -169 471
rect -23 471 23 483
rect -215 -29 -169 -17
rect -119 17 -73 29
rect -311 -483 -265 -471
rect -119 -471 -113 17
rect -79 -471 -73 17
rect -23 -17 -17 471
rect 17 -17 23 471
rect 169 471 215 483
rect -23 -29 23 -17
rect 73 17 119 29
rect -119 -483 -73 -471
rect 73 -471 79 17
rect 113 -471 119 17
rect 169 -17 175 471
rect 209 -17 215 471
rect 361 471 407 483
rect 169 -29 215 -17
rect 265 17 311 29
rect 73 -483 119 -471
rect 265 -471 271 17
rect 305 -471 311 17
rect 361 -17 367 471
rect 401 -17 407 471
rect 553 471 599 483
rect 361 -29 407 -17
rect 457 17 503 29
rect 265 -483 311 -471
rect 457 -471 463 17
rect 497 -471 503 17
rect 553 -17 559 471
rect 593 -17 599 471
rect 553 -29 599 -17
rect 457 -483 503 -471
rect -557 -538 -499 -532
rect -557 -572 -545 -538
rect -511 -572 -499 -538
rect -557 -578 -499 -572
rect -365 -538 -307 -532
rect -365 -572 -353 -538
rect -319 -572 -307 -538
rect -365 -578 -307 -572
rect -173 -538 -115 -532
rect -173 -572 -161 -538
rect -127 -572 -115 -538
rect -173 -578 -115 -572
rect 19 -538 77 -532
rect 19 -572 31 -538
rect 65 -572 77 -538
rect 19 -578 77 -572
rect 211 -538 269 -532
rect 211 -572 223 -538
rect 257 -572 269 -538
rect 211 -578 269 -572
rect 403 -538 461 -532
rect 403 -572 415 -538
rect 449 -572 461 -538
rect 403 -578 461 -572
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.0 l 0.15 m 1 nf 12 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc +50 viadrn -50 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
