magic
tech sky130A
magscale 1 2
timestamp 1698511094
<< nwell >>
rect -1355 -400 1355 400
<< pmos >>
rect -1261 -300 -1061 300
rect -1003 -300 -803 300
rect -745 -300 -545 300
rect -487 -300 -287 300
rect -229 -300 -29 300
rect 29 -300 229 300
rect 287 -300 487 300
rect 545 -300 745 300
rect 803 -300 1003 300
rect 1061 -300 1261 300
<< pdiff >>
rect -1319 288 -1261 300
rect -1319 -288 -1307 288
rect -1273 -288 -1261 288
rect -1319 -300 -1261 -288
rect -1061 288 -1003 300
rect -1061 -288 -1049 288
rect -1015 -288 -1003 288
rect -1061 -300 -1003 -288
rect -803 288 -745 300
rect -803 -288 -791 288
rect -757 -288 -745 288
rect -803 -300 -745 -288
rect -545 288 -487 300
rect -545 -288 -533 288
rect -499 -288 -487 288
rect -545 -300 -487 -288
rect -287 288 -229 300
rect -287 -288 -275 288
rect -241 -288 -229 288
rect -287 -300 -229 -288
rect -29 288 29 300
rect -29 -288 -17 288
rect 17 -288 29 288
rect -29 -300 29 -288
rect 229 288 287 300
rect 229 -288 241 288
rect 275 -288 287 288
rect 229 -300 287 -288
rect 487 288 545 300
rect 487 -288 499 288
rect 533 -288 545 288
rect 487 -300 545 -288
rect 745 288 803 300
rect 745 -288 757 288
rect 791 -288 803 288
rect 745 -300 803 -288
rect 1003 288 1061 300
rect 1003 -288 1015 288
rect 1049 -288 1061 288
rect 1003 -300 1061 -288
rect 1261 288 1319 300
rect 1261 -288 1273 288
rect 1307 -288 1319 288
rect 1261 -300 1319 -288
<< pdiffc >>
rect -1307 -288 -1273 288
rect -1049 -288 -1015 288
rect -791 -288 -757 288
rect -533 -288 -499 288
rect -275 -288 -241 288
rect -17 -288 17 288
rect 241 -288 275 288
rect 499 -288 533 288
rect 757 -288 791 288
rect 1015 -288 1049 288
rect 1273 -288 1307 288
<< poly >>
rect -1261 381 -1061 397
rect -1261 347 -1245 381
rect -1077 347 -1061 381
rect -1261 300 -1061 347
rect -1003 381 -803 397
rect -1003 347 -987 381
rect -819 347 -803 381
rect -1003 300 -803 347
rect -745 381 -545 397
rect -745 347 -729 381
rect -561 347 -545 381
rect -745 300 -545 347
rect -487 381 -287 397
rect -487 347 -471 381
rect -303 347 -287 381
rect -487 300 -287 347
rect -229 381 -29 397
rect -229 347 -213 381
rect -45 347 -29 381
rect -229 300 -29 347
rect 29 381 229 397
rect 29 347 45 381
rect 213 347 229 381
rect 29 300 229 347
rect 287 381 487 397
rect 287 347 303 381
rect 471 347 487 381
rect 287 300 487 347
rect 545 381 745 397
rect 545 347 561 381
rect 729 347 745 381
rect 545 300 745 347
rect 803 381 1003 397
rect 803 347 819 381
rect 987 347 1003 381
rect 803 300 1003 347
rect 1061 381 1261 397
rect 1061 347 1077 381
rect 1245 347 1261 381
rect 1061 300 1261 347
rect -1261 -347 -1061 -300
rect -1261 -381 -1245 -347
rect -1077 -381 -1061 -347
rect -1261 -397 -1061 -381
rect -1003 -347 -803 -300
rect -1003 -381 -987 -347
rect -819 -381 -803 -347
rect -1003 -397 -803 -381
rect -745 -347 -545 -300
rect -745 -381 -729 -347
rect -561 -381 -545 -347
rect -745 -397 -545 -381
rect -487 -347 -287 -300
rect -487 -381 -471 -347
rect -303 -381 -287 -347
rect -487 -397 -287 -381
rect -229 -347 -29 -300
rect -229 -381 -213 -347
rect -45 -381 -29 -347
rect -229 -397 -29 -381
rect 29 -347 229 -300
rect 29 -381 45 -347
rect 213 -381 229 -347
rect 29 -397 229 -381
rect 287 -347 487 -300
rect 287 -381 303 -347
rect 471 -381 487 -347
rect 287 -397 487 -381
rect 545 -347 745 -300
rect 545 -381 561 -347
rect 729 -381 745 -347
rect 545 -397 745 -381
rect 803 -347 1003 -300
rect 803 -381 819 -347
rect 987 -381 1003 -347
rect 803 -397 1003 -381
rect 1061 -347 1261 -300
rect 1061 -381 1077 -347
rect 1245 -381 1261 -347
rect 1061 -397 1261 -381
<< polycont >>
rect -1245 347 -1077 381
rect -987 347 -819 381
rect -729 347 -561 381
rect -471 347 -303 381
rect -213 347 -45 381
rect 45 347 213 381
rect 303 347 471 381
rect 561 347 729 381
rect 819 347 987 381
rect 1077 347 1245 381
rect -1245 -381 -1077 -347
rect -987 -381 -819 -347
rect -729 -381 -561 -347
rect -471 -381 -303 -347
rect -213 -381 -45 -347
rect 45 -381 213 -347
rect 303 -381 471 -347
rect 561 -381 729 -347
rect 819 -381 987 -347
rect 1077 -381 1245 -347
<< locali >>
rect -1261 347 -1245 381
rect -1077 347 -1061 381
rect -1003 347 -987 381
rect -819 347 -803 381
rect -745 347 -729 381
rect -561 347 -545 381
rect -487 347 -471 381
rect -303 347 -287 381
rect -229 347 -213 381
rect -45 347 -29 381
rect 29 347 45 381
rect 213 347 229 381
rect 287 347 303 381
rect 471 347 487 381
rect 545 347 561 381
rect 729 347 745 381
rect 803 347 819 381
rect 987 347 1003 381
rect 1061 347 1077 381
rect 1245 347 1261 381
rect -1307 288 -1273 304
rect -1307 -304 -1273 -288
rect -1049 288 -1015 304
rect -1049 -304 -1015 -288
rect -791 288 -757 304
rect -791 -304 -757 -288
rect -533 288 -499 304
rect -533 -304 -499 -288
rect -275 288 -241 304
rect -275 -304 -241 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 241 288 275 304
rect 241 -304 275 -288
rect 499 288 533 304
rect 499 -304 533 -288
rect 757 288 791 304
rect 757 -304 791 -288
rect 1015 288 1049 304
rect 1015 -304 1049 -288
rect 1273 288 1307 304
rect 1273 -304 1307 -288
rect -1261 -381 -1245 -347
rect -1077 -381 -1061 -347
rect -1003 -381 -987 -347
rect -819 -381 -803 -347
rect -745 -381 -729 -347
rect -561 -381 -545 -347
rect -487 -381 -471 -347
rect -303 -381 -287 -347
rect -229 -381 -213 -347
rect -45 -381 -29 -347
rect 29 -381 45 -347
rect 213 -381 229 -347
rect 287 -381 303 -347
rect 471 -381 487 -347
rect 545 -381 561 -347
rect 729 -381 745 -347
rect 803 -381 819 -347
rect 987 -381 1003 -347
rect 1061 -381 1077 -347
rect 1245 -381 1261 -347
<< viali >>
rect -1245 347 -1077 381
rect -987 347 -819 381
rect -729 347 -561 381
rect -471 347 -303 381
rect -213 347 -45 381
rect 45 347 213 381
rect 303 347 471 381
rect 561 347 729 381
rect 819 347 987 381
rect 1077 347 1245 381
rect -1307 -17 -1273 271
rect -1049 -271 -1015 17
rect -791 -17 -757 271
rect -533 -271 -499 17
rect -275 -17 -241 271
rect -17 -271 17 17
rect 241 -17 275 271
rect 499 -271 533 17
rect 757 -17 791 271
rect 1015 -271 1049 17
rect 1273 -17 1307 271
rect -1245 -381 -1077 -347
rect -987 -381 -819 -347
rect -729 -381 -561 -347
rect -471 -381 -303 -347
rect -213 -381 -45 -347
rect 45 -381 213 -347
rect 303 -381 471 -347
rect 561 -381 729 -347
rect 819 -381 987 -347
rect 1077 -381 1245 -347
<< metal1 >>
rect -1257 381 -1065 387
rect -1257 347 -1245 381
rect -1077 347 -1065 381
rect -1257 341 -1065 347
rect -999 381 -807 387
rect -999 347 -987 381
rect -819 347 -807 381
rect -999 341 -807 347
rect -741 381 -549 387
rect -741 347 -729 381
rect -561 347 -549 381
rect -741 341 -549 347
rect -483 381 -291 387
rect -483 347 -471 381
rect -303 347 -291 381
rect -483 341 -291 347
rect -225 381 -33 387
rect -225 347 -213 381
rect -45 347 -33 381
rect -225 341 -33 347
rect 33 381 225 387
rect 33 347 45 381
rect 213 347 225 381
rect 33 341 225 347
rect 291 381 483 387
rect 291 347 303 381
rect 471 347 483 381
rect 291 341 483 347
rect 549 381 741 387
rect 549 347 561 381
rect 729 347 741 381
rect 549 341 741 347
rect 807 381 999 387
rect 807 347 819 381
rect 987 347 999 381
rect 807 341 999 347
rect 1065 381 1257 387
rect 1065 347 1077 381
rect 1245 347 1257 381
rect 1065 341 1257 347
rect -1313 271 -1267 283
rect -1313 -17 -1307 271
rect -1273 -17 -1267 271
rect -797 271 -751 283
rect -1313 -29 -1267 -17
rect -1055 17 -1009 29
rect -1055 -271 -1049 17
rect -1015 -271 -1009 17
rect -797 -17 -791 271
rect -757 -17 -751 271
rect -281 271 -235 283
rect -797 -29 -751 -17
rect -539 17 -493 29
rect -1055 -283 -1009 -271
rect -539 -271 -533 17
rect -499 -271 -493 17
rect -281 -17 -275 271
rect -241 -17 -235 271
rect 235 271 281 283
rect -281 -29 -235 -17
rect -23 17 23 29
rect -539 -283 -493 -271
rect -23 -271 -17 17
rect 17 -271 23 17
rect 235 -17 241 271
rect 275 -17 281 271
rect 751 271 797 283
rect 235 -29 281 -17
rect 493 17 539 29
rect -23 -283 23 -271
rect 493 -271 499 17
rect 533 -271 539 17
rect 751 -17 757 271
rect 791 -17 797 271
rect 1267 271 1313 283
rect 751 -29 797 -17
rect 1009 17 1055 29
rect 493 -283 539 -271
rect 1009 -271 1015 17
rect 1049 -271 1055 17
rect 1267 -17 1273 271
rect 1307 -17 1313 271
rect 1267 -29 1313 -17
rect 1009 -283 1055 -271
rect -1257 -347 -1065 -341
rect -1257 -381 -1245 -347
rect -1077 -381 -1065 -347
rect -1257 -387 -1065 -381
rect -999 -347 -807 -341
rect -999 -381 -987 -347
rect -819 -381 -807 -347
rect -999 -387 -807 -381
rect -741 -347 -549 -341
rect -741 -381 -729 -347
rect -561 -381 -549 -347
rect -741 -387 -549 -381
rect -483 -347 -291 -341
rect -483 -381 -471 -347
rect -303 -381 -291 -347
rect -483 -387 -291 -381
rect -225 -347 -33 -341
rect -225 -381 -213 -347
rect -45 -381 -33 -347
rect -225 -387 -33 -381
rect 33 -347 225 -341
rect 33 -381 45 -347
rect 213 -381 225 -347
rect 33 -387 225 -381
rect 291 -347 483 -341
rect 291 -381 303 -347
rect 471 -381 483 -347
rect 291 -387 483 -381
rect 549 -347 741 -341
rect 549 -381 561 -347
rect 729 -381 741 -347
rect 549 -387 741 -381
rect 807 -347 999 -341
rect 807 -381 819 -347
rect 987 -381 999 -347
rect 807 -387 999 -381
rect 1065 -347 1257 -341
rect 1065 -381 1077 -347
rect 1245 -381 1257 -347
rect 1065 -387 1257 -381
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.0 l 1.0 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc +50 viadrn -50 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
