magic
tech sky130A
timestamp 1698511094
<< pwell >>
rect -664 -155 664 155
<< nmos >>
rect -566 -50 -466 50
rect -437 -50 -337 50
rect -308 -50 -208 50
rect -179 -50 -79 50
rect -50 -50 50 50
rect 79 -50 179 50
rect 208 -50 308 50
rect 337 -50 437 50
rect 466 -50 566 50
<< ndiff >>
rect -595 44 -566 50
rect -595 -44 -589 44
rect -572 -44 -566 44
rect -595 -50 -566 -44
rect -466 44 -437 50
rect -466 -44 -460 44
rect -443 -44 -437 44
rect -466 -50 -437 -44
rect -337 44 -308 50
rect -337 -44 -331 44
rect -314 -44 -308 44
rect -337 -50 -308 -44
rect -208 44 -179 50
rect -208 -44 -202 44
rect -185 -44 -179 44
rect -208 -50 -179 -44
rect -79 44 -50 50
rect -79 -44 -73 44
rect -56 -44 -50 44
rect -79 -50 -50 -44
rect 50 44 79 50
rect 50 -44 56 44
rect 73 -44 79 44
rect 50 -50 79 -44
rect 179 44 208 50
rect 179 -44 185 44
rect 202 -44 208 44
rect 179 -50 208 -44
rect 308 44 337 50
rect 308 -44 314 44
rect 331 -44 337 44
rect 308 -50 337 -44
rect 437 44 466 50
rect 437 -44 443 44
rect 460 -44 466 44
rect 437 -50 466 -44
rect 566 44 595 50
rect 566 -44 572 44
rect 589 -44 595 44
rect 566 -50 595 -44
<< ndiffc >>
rect -589 -44 -572 44
rect -460 -44 -443 44
rect -331 -44 -314 44
rect -202 -44 -185 44
rect -73 -44 -56 44
rect 56 -44 73 44
rect 185 -44 202 44
rect 314 -44 331 44
rect 443 -44 460 44
rect 572 -44 589 44
<< psubdiff >>
rect -646 120 -598 137
rect 598 120 646 137
rect -646 89 -629 120
rect 629 89 646 120
rect -646 -120 -629 -89
rect 629 -120 646 -89
rect -646 -137 -598 -120
rect 598 -137 646 -120
<< psubdiffcont >>
rect -598 120 598 137
rect -646 -89 -629 89
rect 629 -89 646 89
rect -598 -137 598 -120
<< poly >>
rect -566 86 -466 94
rect -566 69 -558 86
rect -474 69 -466 86
rect -566 50 -466 69
rect -437 86 -337 94
rect -437 69 -429 86
rect -345 69 -337 86
rect -437 50 -337 69
rect -308 86 -208 94
rect -308 69 -300 86
rect -216 69 -208 86
rect -308 50 -208 69
rect -179 86 -79 94
rect -179 69 -171 86
rect -87 69 -79 86
rect -179 50 -79 69
rect -50 86 50 94
rect -50 69 -42 86
rect 42 69 50 86
rect -50 50 50 69
rect 79 86 179 94
rect 79 69 87 86
rect 171 69 179 86
rect 79 50 179 69
rect 208 86 308 94
rect 208 69 216 86
rect 300 69 308 86
rect 208 50 308 69
rect 337 86 437 94
rect 337 69 345 86
rect 429 69 437 86
rect 337 50 437 69
rect 466 86 566 94
rect 466 69 474 86
rect 558 69 566 86
rect 466 50 566 69
rect -566 -69 -466 -50
rect -566 -86 -558 -69
rect -474 -86 -466 -69
rect -566 -94 -466 -86
rect -437 -69 -337 -50
rect -437 -86 -429 -69
rect -345 -86 -337 -69
rect -437 -94 -337 -86
rect -308 -69 -208 -50
rect -308 -86 -300 -69
rect -216 -86 -208 -69
rect -308 -94 -208 -86
rect -179 -69 -79 -50
rect -179 -86 -171 -69
rect -87 -86 -79 -69
rect -179 -94 -79 -86
rect -50 -69 50 -50
rect -50 -86 -42 -69
rect 42 -86 50 -69
rect -50 -94 50 -86
rect 79 -69 179 -50
rect 79 -86 87 -69
rect 171 -86 179 -69
rect 79 -94 179 -86
rect 208 -69 308 -50
rect 208 -86 216 -69
rect 300 -86 308 -69
rect 208 -94 308 -86
rect 337 -69 437 -50
rect 337 -86 345 -69
rect 429 -86 437 -69
rect 337 -94 437 -86
rect 466 -69 566 -50
rect 466 -86 474 -69
rect 558 -86 566 -69
rect 466 -94 566 -86
<< polycont >>
rect -558 69 -474 86
rect -429 69 -345 86
rect -300 69 -216 86
rect -171 69 -87 86
rect -42 69 42 86
rect 87 69 171 86
rect 216 69 300 86
rect 345 69 429 86
rect 474 69 558 86
rect -558 -86 -474 -69
rect -429 -86 -345 -69
rect -300 -86 -216 -69
rect -171 -86 -87 -69
rect -42 -86 42 -69
rect 87 -86 171 -69
rect 216 -86 300 -69
rect 345 -86 429 -69
rect 474 -86 558 -69
<< locali >>
rect -646 120 -598 137
rect 598 120 646 137
rect -646 89 -629 120
rect 629 89 646 120
rect -566 69 -558 86
rect -474 69 -466 86
rect -437 69 -429 86
rect -345 69 -337 86
rect -308 69 -300 86
rect -216 69 -208 86
rect -179 69 -171 86
rect -87 69 -79 86
rect -50 69 -42 86
rect 42 69 50 86
rect 79 69 87 86
rect 171 69 179 86
rect 208 69 216 86
rect 300 69 308 86
rect 337 69 345 86
rect 429 69 437 86
rect 466 69 474 86
rect 558 69 566 86
rect -589 44 -572 52
rect -589 -52 -572 -44
rect -460 44 -443 52
rect -460 -52 -443 -44
rect -331 44 -314 52
rect -331 -52 -314 -44
rect -202 44 -185 52
rect -202 -52 -185 -44
rect -73 44 -56 52
rect -73 -52 -56 -44
rect 56 44 73 52
rect 56 -52 73 -44
rect 185 44 202 52
rect 185 -52 202 -44
rect 314 44 331 52
rect 314 -52 331 -44
rect 443 44 460 52
rect 443 -52 460 -44
rect 572 44 589 52
rect 572 -52 589 -44
rect -566 -86 -558 -69
rect -474 -86 -466 -69
rect -437 -86 -429 -69
rect -345 -86 -337 -69
rect -308 -86 -300 -69
rect -216 -86 -208 -69
rect -179 -86 -171 -69
rect -87 -86 -79 -69
rect -50 -86 -42 -69
rect 42 -86 50 -69
rect 79 -86 87 -69
rect 171 -86 179 -69
rect 208 -86 216 -69
rect 300 -86 308 -69
rect 337 -86 345 -69
rect 429 -86 437 -69
rect 466 -86 474 -69
rect 558 -86 566 -69
rect -646 -120 -629 -89
rect 629 -120 646 -89
rect -646 -137 -598 -120
rect 598 -137 646 -120
<< viali >>
rect -558 69 -474 86
rect -429 69 -345 86
rect -300 69 -216 86
rect -171 69 -87 86
rect -42 69 42 86
rect 87 69 171 86
rect 216 69 300 86
rect 345 69 429 86
rect 474 69 558 86
rect -589 -44 -572 44
rect -460 -44 -443 44
rect -331 -44 -314 44
rect -202 -44 -185 44
rect -73 -44 -56 44
rect 56 -44 73 44
rect 185 -44 202 44
rect 314 -44 331 44
rect 443 -44 460 44
rect 572 -44 589 44
rect -558 -86 -474 -69
rect -429 -86 -345 -69
rect -300 -86 -216 -69
rect -171 -86 -87 -69
rect -42 -86 42 -69
rect 87 -86 171 -69
rect 216 -86 300 -69
rect 345 -86 429 -69
rect 474 -86 558 -69
<< metal1 >>
rect -564 86 -468 89
rect -564 69 -558 86
rect -474 69 -468 86
rect -564 66 -468 69
rect -435 86 -339 89
rect -435 69 -429 86
rect -345 69 -339 86
rect -435 66 -339 69
rect -306 86 -210 89
rect -306 69 -300 86
rect -216 69 -210 86
rect -306 66 -210 69
rect -177 86 -81 89
rect -177 69 -171 86
rect -87 69 -81 86
rect -177 66 -81 69
rect -48 86 48 89
rect -48 69 -42 86
rect 42 69 48 86
rect -48 66 48 69
rect 81 86 177 89
rect 81 69 87 86
rect 171 69 177 86
rect 81 66 177 69
rect 210 86 306 89
rect 210 69 216 86
rect 300 69 306 86
rect 210 66 306 69
rect 339 86 435 89
rect 339 69 345 86
rect 429 69 435 86
rect 339 66 435 69
rect 468 86 564 89
rect 468 69 474 86
rect 558 69 564 86
rect 468 66 564 69
rect -592 44 -569 50
rect -592 -44 -589 44
rect -572 -44 -569 44
rect -592 -50 -569 -44
rect -463 44 -440 50
rect -463 -44 -460 44
rect -443 -44 -440 44
rect -463 -50 -440 -44
rect -334 44 -311 50
rect -334 -44 -331 44
rect -314 -44 -311 44
rect -334 -50 -311 -44
rect -205 44 -182 50
rect -205 -44 -202 44
rect -185 -44 -182 44
rect -205 -50 -182 -44
rect -76 44 -53 50
rect -76 -44 -73 44
rect -56 -44 -53 44
rect -76 -50 -53 -44
rect 53 44 76 50
rect 53 -44 56 44
rect 73 -44 76 44
rect 53 -50 76 -44
rect 182 44 205 50
rect 182 -44 185 44
rect 202 -44 205 44
rect 182 -50 205 -44
rect 311 44 334 50
rect 311 -44 314 44
rect 331 -44 334 44
rect 311 -50 334 -44
rect 440 44 463 50
rect 440 -44 443 44
rect 460 -44 463 44
rect 440 -50 463 -44
rect 569 44 592 50
rect 569 -44 572 44
rect 589 -44 592 44
rect 569 -50 592 -44
rect -564 -69 -468 -66
rect -564 -86 -558 -69
rect -474 -86 -468 -69
rect -564 -89 -468 -86
rect -435 -69 -339 -66
rect -435 -86 -429 -69
rect -345 -86 -339 -69
rect -435 -89 -339 -86
rect -306 -69 -210 -66
rect -306 -86 -300 -69
rect -216 -86 -210 -69
rect -306 -89 -210 -86
rect -177 -69 -81 -66
rect -177 -86 -171 -69
rect -87 -86 -81 -69
rect -177 -89 -81 -86
rect -48 -69 48 -66
rect -48 -86 -42 -69
rect 42 -86 48 -69
rect -48 -89 48 -86
rect 81 -69 177 -66
rect 81 -86 87 -69
rect 171 -86 177 -69
rect 81 -89 177 -86
rect 210 -69 306 -66
rect 210 -86 216 -69
rect 300 -86 306 -69
rect 210 -89 306 -86
rect 339 -69 435 -66
rect 339 -86 345 -69
rect 429 -86 435 -69
rect 339 -89 435 -86
rect 468 -69 564 -66
rect 468 -86 474 -69
rect 558 -86 564 -69
rect 468 -89 564 -86
<< properties >>
string FIXED_BBOX -637 -128 637 128
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 1.0 m 1 nf 9 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
