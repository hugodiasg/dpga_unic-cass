magic
tech sky130A
magscale 1 2
timestamp 1698525607
<< metal1 >>
rect 550 6840 750 8960
rect 3830 6840 4030 8960
rect 7060 6820 7260 8960
rect 10300 6850 10500 8960
rect 13810 6850 14010 8960
rect 17350 6850 17550 8960
rect 20980 6850 21180 8960
rect 24510 6850 24710 8960
rect 25660 8210 26020 8580
rect 26300 8200 26660 8570
rect 26930 8200 27290 8570
rect 27560 8200 27920 8570
rect 24965 7050 25730 7060
rect 24965 6920 25010 7050
rect 25140 7040 25730 7050
rect 25140 6920 25210 7040
rect 24965 6910 25210 6920
rect 25340 7030 25730 7040
rect 25340 6910 25400 7030
rect 24965 6900 25400 6910
rect 25530 6900 25730 7030
rect 24965 6870 25730 6900
rect 24965 6740 25020 6870
rect 25150 6850 25730 6870
rect 25150 6740 25200 6850
rect 24965 6720 25200 6740
rect 25330 6840 25730 6850
rect 25330 6720 25380 6840
rect 24965 6710 25380 6720
rect 25510 6710 25730 6840
rect 24965 6650 25730 6710
rect 25980 6690 26340 7060
rect 26610 6670 26970 7040
rect 27250 6670 27610 7040
rect 28430 7030 28700 7040
rect 27850 6630 28700 7030
rect 28430 5990 28700 6630
rect 28500 5270 28700 5990
rect 29000 5500 29200 8950
rect 31850 6830 32050 7050
rect 31850 6690 31880 6830
rect 32030 6690 32050 6830
rect 31850 6680 32050 6690
rect 35030 5310 35230 5500
rect 28500 5070 29210 5270
rect 28500 4230 29210 4430
rect -200 2950 0 3150
rect -200 2010 0 2200
rect 13850 -450 14050 40
rect 28500 -490 28700 4230
rect 28890 3400 28900 3600
rect 29200 3400 29210 3600
<< via1 >>
rect 25010 6920 25140 7050
rect 25210 6910 25340 7040
rect 25400 6900 25530 7030
rect 25020 6740 25150 6870
rect 25200 6720 25330 6850
rect 25380 6710 25510 6840
rect 31880 6690 32030 6830
rect 28900 3400 29200 3600
<< metal2 >>
rect 28330 7290 34810 7710
rect 28330 7080 28750 7290
rect 24990 7050 28750 7080
rect 24990 6920 25010 7050
rect 25140 7040 28750 7050
rect 25140 6920 25210 7040
rect 24990 6910 25210 6920
rect 25340 7030 28750 7040
rect 25340 6910 25400 7030
rect 24990 6900 25400 6910
rect 25530 6900 28750 7030
rect 24990 6870 28750 6900
rect 24990 6740 25020 6870
rect 25150 6850 28750 6870
rect 25150 6740 25200 6850
rect 24990 6720 25200 6740
rect 25330 6840 28750 6850
rect 25330 6720 25380 6840
rect 24990 6710 25380 6720
rect 25510 6710 28750 6840
rect 24990 6690 28750 6710
rect 31860 6840 32060 6850
rect 31860 6700 31870 6840
rect 32020 6830 32060 6840
rect 31860 6690 31880 6700
rect 32030 6690 32060 6830
rect 24990 6660 28700 6690
rect 31860 6660 32060 6690
rect 34730 5340 34810 7290
rect 28900 3600 29200 3610
rect 28900 3390 29200 3400
<< via2 >>
rect 31870 6830 32020 6840
rect 31870 6700 31880 6830
rect 31880 6700 32020 6830
rect 28900 3400 29200 3600
<< metal3 >>
rect 28110 6840 32030 6860
rect 28110 6700 31870 6840
rect 32020 6700 32030 6840
rect 28110 6640 32030 6700
rect 28110 3160 28330 6640
rect 25080 2940 28330 3160
rect 28890 3605 29110 3710
rect 28890 3600 29210 3605
rect 28890 3400 28900 3600
rect 29200 3400 29210 3600
rect 28890 3395 29210 3400
rect 28890 2220 29110 3395
rect 24890 2000 29110 2220
use sky130_fd_pr__res_xhigh_po_0p35_2TH3B8  XR8 /foss/designs/projects/dpga2/magic/ota_digpot/digpot
timestamp 1698522189
transform 1 0 26794 0 1 7630
box -1314 -1140 1314 1140
use digpotp  digpotp_0 /foss/designs/projects/dpga2/magic/ota_digpot/digpot
timestamp 1698522569
transform 1 0 -9350 0 1 -1550
box 9350 1550 38050 8600
use ota  ota_0 /foss/designs/projects/dpga2/magic/ota_digpot/ota
timestamp 1698525106
transform 1 0 24200 0 1 560
box 4800 -160 10830 6320
<< labels >>
flabel metal1 35030 5310 35230 5500 0 FreeSans 1600 0 0 0 out
port 4 nsew
flabel metal1 -200 2010 0 2200 0 FreeSans 1600 0 0 0 gnd
port 5 nsew
flabel metal1 -200 2950 0 3150 0 FreeSans 1600 0 0 0 vd
port 14 nsew
flabel metal1 28500 -490 28700 -300 0 FreeSans 1600 0 0 0 inp
port 2 nsew
flabel metal1 13850 -450 14050 -260 0 FreeSans 1600 0 0 0 inn
port 1 nsew
flabel metal1 29000 8760 29200 8950 0 FreeSans 1600 0 0 0 ib
port 3 nsew
flabel metal1 24510 8760 24710 8960 0 FreeSans 1600 0 0 0 c0
port 6 nsew
flabel metal1 20980 8760 21180 8960 0 FreeSans 1600 0 0 0 c1
port 7 nsew
flabel metal1 17350 8760 17550 8960 0 FreeSans 1600 0 0 0 c2
port 8 nsew
flabel metal1 13810 8760 14010 8960 0 FreeSans 1600 0 0 0 c3
port 9 nsew
flabel metal1 10300 8760 10500 8960 0 FreeSans 1600 0 0 0 c4
port 10 nsew
flabel metal1 7060 8760 7260 8960 0 FreeSans 1600 0 0 0 c5
port 11 nsew
flabel metal1 3830 8760 4030 8960 0 FreeSans 1600 0 0 0 c6
port 12 nsew
flabel metal1 550 8760 750 8960 0 FreeSans 1600 0 0 0 c7
port 13 nsew
<< end >>
