magic
tech sky130A
magscale 1 2
timestamp 1698520721
<< pwell >>
rect -201 -1140 201 1140
<< psubdiff >>
rect -165 1070 -69 1104
rect 69 1070 165 1104
rect -165 1008 -131 1070
rect 131 1008 165 1070
rect -165 -1070 -131 -1008
rect 131 -1070 165 -1008
rect -165 -1104 -69 -1070
rect 69 -1104 165 -1070
<< psubdiffcont >>
rect -69 1070 69 1104
rect -165 -1008 -131 1008
rect 131 -1008 165 1008
rect -69 -1104 69 -1070
<< xpolycontact >>
rect -35 542 35 974
rect -35 -974 35 -542
<< xpolyres >>
rect -35 -542 35 542
<< locali >>
rect -165 1070 -69 1104
rect 69 1070 165 1104
rect -165 1008 -131 1070
rect 131 1008 165 1070
rect -165 -1070 -131 -1008
rect 131 -1070 165 -1008
rect -165 -1104 -69 -1070
rect 69 -1104 165 -1070
<< viali >>
rect -19 559 19 956
rect -19 -956 19 -559
<< metal1 >>
rect -25 956 25 968
rect -25 559 -19 956
rect 19 559 25 956
rect -25 547 25 559
rect -25 -559 25 -547
rect -25 -956 -19 -559
rect 19 -956 25 -559
rect -25 -968 25 -956
<< res0p35 >>
rect -37 -544 37 544
<< properties >>
string FIXED_BBOX -148 -1087 148 1087
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 5.42 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 32.046k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
