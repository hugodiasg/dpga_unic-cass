magic
tech sky130A
magscale 1 2
timestamp 1698430756
<< obsli1 >>
rect 1104 2159 16376 17425
<< obsm1 >>
rect 1104 2128 16376 17456
<< metal2 >>
rect 2226 18856 2282 19656
rect 6550 18856 6606 19656
rect 10874 18856 10930 19656
rect 15198 18856 15254 19656
rect 1306 0 1362 800
rect 3422 0 3478 800
rect 5538 0 5594 800
rect 7654 0 7710 800
rect 9770 0 9826 800
rect 11886 0 11942 800
rect 14002 0 14058 800
rect 16118 0 16174 800
<< obsm2 >>
rect 1308 18800 2170 18986
rect 2338 18800 6494 18986
rect 6662 18800 10818 18986
rect 10986 18800 15142 18986
rect 15310 18800 16160 18986
rect 1308 856 16160 18800
rect 1418 800 3366 856
rect 3534 800 5482 856
rect 5650 800 7598 856
rect 7766 800 9714 856
rect 9882 800 11830 856
rect 11998 800 13946 856
rect 14114 800 16062 856
<< obsm3 >>
rect 2855 2143 15285 17441
<< metal4 >>
rect 2853 2128 3173 17456
rect 3513 2128 3833 17456
rect 6671 2128 6991 17456
rect 7331 2128 7651 17456
rect 10489 2128 10809 17456
rect 11149 2128 11469 17456
rect 14307 2128 14627 17456
rect 14967 2128 15287 17456
<< metal5 >>
rect 1056 16004 16424 16324
rect 1056 15344 16424 15664
rect 1056 12196 16424 12516
rect 1056 11536 16424 11856
rect 1056 8388 16424 8708
rect 1056 7728 16424 8048
rect 1056 4580 16424 4900
rect 1056 3920 16424 4240
<< labels >>
rlabel metal4 s 3513 2128 3833 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7331 2128 7651 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 11149 2128 11469 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 14967 2128 15287 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 4580 16424 4900 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 8388 16424 8708 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 12196 16424 12516 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 16004 16424 16324 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 2853 2128 3173 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 6671 2128 6991 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 10489 2128 10809 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 14307 2128 14627 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3920 16424 4240 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 7728 16424 8048 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 11536 16424 11856 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 15344 16424 15664 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 1306 0 1362 800 6 data[0]
port 3 nsew signal output
rlabel metal2 s 3422 0 3478 800 6 data[1]
port 4 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 data[2]
port 5 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 data[3]
port 6 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 data[4]
port 7 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 data[5]
port 8 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 data[6]
port 9 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 data[7]
port 10 nsew signal output
rlabel metal2 s 15198 18856 15254 19656 6 reset
port 11 nsew signal input
rlabel metal2 s 6550 18856 6606 19656 6 sclk
port 12 nsew signal input
rlabel metal2 s 10874 18856 10930 19656 6 sdi
port 13 nsew signal input
rlabel metal2 s 2226 18856 2282 19656 6 ss
port 14 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 17512 19656
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 311804
string GDS_FILE /shift/openlane/sr/runs/RUN_2023.10.27_18.18.11/results/signoff/sr.magic.gds
string GDS_START 77600
<< end >>

