magic
tech sky130A
magscale 1 2
timestamp 1698520721
<< pwell >>
rect -201 -2820 201 2820
<< psubdiff >>
rect -165 2750 -69 2784
rect 69 2750 165 2784
rect -165 2688 -131 2750
rect 131 2688 165 2750
rect -165 -2750 -131 -2688
rect 131 -2750 165 -2688
rect -165 -2784 -69 -2750
rect 69 -2784 165 -2750
<< psubdiffcont >>
rect -69 2750 69 2784
rect -165 -2688 -131 2688
rect 131 -2688 165 2688
rect -69 -2784 69 -2750
<< xpolycontact >>
rect -35 2222 35 2654
rect -35 -2654 35 -2222
<< xpolyres >>
rect -35 -2222 35 2222
<< locali >>
rect -165 2750 -69 2784
rect 69 2750 165 2784
rect -165 2688 -131 2750
rect 131 2688 165 2750
rect -165 -2750 -131 -2688
rect 131 -2750 165 -2688
rect -165 -2784 -69 -2750
rect 69 -2784 165 -2750
<< viali >>
rect -19 2239 19 2636
rect -19 -2636 19 -2239
<< metal1 >>
rect -25 2636 25 2648
rect -25 2239 -19 2636
rect 19 2239 25 2636
rect -25 2227 25 2239
rect -25 -2239 25 -2227
rect -25 -2636 -19 -2239
rect 19 -2636 25 -2239
rect -25 -2648 25 -2636
<< res0p35 >>
rect -37 -2224 37 2224
<< properties >>
string FIXED_BBOX -148 -2767 148 2767
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 22.22 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 128.046k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
